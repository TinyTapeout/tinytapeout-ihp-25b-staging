module tt_um_rejunity_atari2600 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire \atari2600.address_bus_r[0] ;
 wire \atari2600.address_bus_r[10] ;
 wire \atari2600.address_bus_r[11] ;
 wire \atari2600.address_bus_r[12] ;
 wire \atari2600.address_bus_r[1] ;
 wire \atari2600.address_bus_r[2] ;
 wire \atari2600.address_bus_r[3] ;
 wire \atari2600.address_bus_r[4] ;
 wire \atari2600.address_bus_r[5] ;
 wire \atari2600.address_bus_r[6] ;
 wire \atari2600.address_bus_r[7] ;
 wire \atari2600.address_bus_r[8] ;
 wire \atari2600.address_bus_r[9] ;
 wire \atari2600.clk_counter[0] ;
 wire \atari2600.clk_counter[1] ;
 wire \atari2600.clk_counter[2] ;
 wire \atari2600.clk_counter[3] ;
 wire \atari2600.clk_counter[4] ;
 wire \atari2600.clk_counter[5] ;
 wire \atari2600.clk_counter[6] ;
 wire \atari2600.clk_counter[7] ;
 wire \atari2600.clk_counter[8] ;
 wire \atari2600.cpu.ABH[0] ;
 wire \atari2600.cpu.ABH[1] ;
 wire \atari2600.cpu.ABH[2] ;
 wire \atari2600.cpu.ABH[3] ;
 wire \atari2600.cpu.ABH[4] ;
 wire \atari2600.cpu.ABH[5] ;
 wire \atari2600.cpu.ABH[6] ;
 wire \atari2600.cpu.ABH[7] ;
 wire \atari2600.cpu.ABL[0] ;
 wire \atari2600.cpu.ABL[1] ;
 wire \atari2600.cpu.ABL[2] ;
 wire \atari2600.cpu.ABL[3] ;
 wire \atari2600.cpu.ABL[4] ;
 wire \atari2600.cpu.ABL[5] ;
 wire \atari2600.cpu.ABL[6] ;
 wire \atari2600.cpu.ABL[7] ;
 wire \atari2600.cpu.ADD[0] ;
 wire \atari2600.cpu.ADD[1] ;
 wire \atari2600.cpu.ADD[2] ;
 wire \atari2600.cpu.ADD[3] ;
 wire \atari2600.cpu.ADD[4] ;
 wire \atari2600.cpu.ADD[5] ;
 wire \atari2600.cpu.ADD[6] ;
 wire \atari2600.cpu.ADD[7] ;
 wire \atari2600.cpu.ALU.AI7 ;
 wire \atari2600.cpu.ALU.BI7 ;
 wire \atari2600.cpu.ALU.CO ;
 wire \atari2600.cpu.ALU.HC ;
 wire \atari2600.cpu.AXYS[0][0] ;
 wire \atari2600.cpu.AXYS[0][1] ;
 wire \atari2600.cpu.AXYS[0][2] ;
 wire \atari2600.cpu.AXYS[0][3] ;
 wire \atari2600.cpu.AXYS[0][4] ;
 wire \atari2600.cpu.AXYS[0][5] ;
 wire \atari2600.cpu.AXYS[0][6] ;
 wire \atari2600.cpu.AXYS[0][7] ;
 wire \atari2600.cpu.AXYS[1][0] ;
 wire \atari2600.cpu.AXYS[1][1] ;
 wire \atari2600.cpu.AXYS[1][2] ;
 wire \atari2600.cpu.AXYS[1][3] ;
 wire \atari2600.cpu.AXYS[1][4] ;
 wire \atari2600.cpu.AXYS[1][5] ;
 wire \atari2600.cpu.AXYS[1][6] ;
 wire \atari2600.cpu.AXYS[1][7] ;
 wire \atari2600.cpu.AXYS[2][0] ;
 wire \atari2600.cpu.AXYS[2][1] ;
 wire \atari2600.cpu.AXYS[2][2] ;
 wire \atari2600.cpu.AXYS[2][3] ;
 wire \atari2600.cpu.AXYS[2][4] ;
 wire \atari2600.cpu.AXYS[2][5] ;
 wire \atari2600.cpu.AXYS[2][6] ;
 wire \atari2600.cpu.AXYS[2][7] ;
 wire \atari2600.cpu.AXYS[3][0] ;
 wire \atari2600.cpu.AXYS[3][1] ;
 wire \atari2600.cpu.AXYS[3][2] ;
 wire \atari2600.cpu.AXYS[3][3] ;
 wire \atari2600.cpu.AXYS[3][4] ;
 wire \atari2600.cpu.AXYS[3][5] ;
 wire \atari2600.cpu.AXYS[3][6] ;
 wire \atari2600.cpu.AXYS[3][7] ;
 wire \atari2600.cpu.C ;
 wire \atari2600.cpu.D ;
 wire \atari2600.cpu.DIHOLD[0] ;
 wire \atari2600.cpu.DIHOLD[1] ;
 wire \atari2600.cpu.DIHOLD[2] ;
 wire \atari2600.cpu.DIHOLD[3] ;
 wire \atari2600.cpu.DIHOLD[4] ;
 wire \atari2600.cpu.DIHOLD[5] ;
 wire \atari2600.cpu.DIHOLD[6] ;
 wire \atari2600.cpu.DIHOLD[7] ;
 wire \atari2600.cpu.DIMUX[0] ;
 wire \atari2600.cpu.DIMUX[1] ;
 wire \atari2600.cpu.DIMUX[2] ;
 wire \atari2600.cpu.DIMUX[3] ;
 wire \atari2600.cpu.DIMUX[4] ;
 wire \atari2600.cpu.DIMUX[5] ;
 wire \atari2600.cpu.DIMUX[6] ;
 wire \atari2600.cpu.DIMUX[7] ;
 wire \atari2600.cpu.DI[0] ;
 wire \atari2600.cpu.DI[1] ;
 wire \atari2600.cpu.DI[2] ;
 wire \atari2600.cpu.DI[3] ;
 wire \atari2600.cpu.DI[4] ;
 wire \atari2600.cpu.DI[5] ;
 wire \atari2600.cpu.DI[6] ;
 wire \atari2600.cpu.DI[7] ;
 wire \atari2600.cpu.I ;
 wire \atari2600.cpu.IRHOLD[0] ;
 wire \atari2600.cpu.IRHOLD[1] ;
 wire \atari2600.cpu.IRHOLD[2] ;
 wire \atari2600.cpu.IRHOLD[3] ;
 wire \atari2600.cpu.IRHOLD[4] ;
 wire \atari2600.cpu.IRHOLD[5] ;
 wire \atari2600.cpu.IRHOLD[6] ;
 wire \atari2600.cpu.IRHOLD[7] ;
 wire \atari2600.cpu.IRHOLD_valid ;
 wire \atari2600.cpu.N ;
 wire \atari2600.cpu.PC[0] ;
 wire \atari2600.cpu.PC[10] ;
 wire \atari2600.cpu.PC[11] ;
 wire \atari2600.cpu.PC[12] ;
 wire \atari2600.cpu.PC[13] ;
 wire \atari2600.cpu.PC[14] ;
 wire \atari2600.cpu.PC[15] ;
 wire \atari2600.cpu.PC[1] ;
 wire \atari2600.cpu.PC[2] ;
 wire \atari2600.cpu.PC[3] ;
 wire \atari2600.cpu.PC[4] ;
 wire \atari2600.cpu.PC[5] ;
 wire \atari2600.cpu.PC[6] ;
 wire \atari2600.cpu.PC[7] ;
 wire \atari2600.cpu.PC[8] ;
 wire \atari2600.cpu.PC[9] ;
 wire \atari2600.cpu.V ;
 wire \atari2600.cpu.Z ;
 wire \atari2600.cpu.adc_bcd ;
 wire \atari2600.cpu.adc_sbc ;
 wire \atari2600.cpu.adj_bcd ;
 wire \atari2600.cpu.backwards ;
 wire \atari2600.cpu.bit_ins ;
 wire \atari2600.cpu.clc ;
 wire \atari2600.cpu.cld ;
 wire \atari2600.cpu.cli ;
 wire \atari2600.cpu.clv ;
 wire \atari2600.cpu.compare ;
 wire \atari2600.cpu.cond_code[0] ;
 wire \atari2600.cpu.cond_code[1] ;
 wire \atari2600.cpu.cond_code[2] ;
 wire \atari2600.cpu.dst_reg[0] ;
 wire \atari2600.cpu.dst_reg[1] ;
 wire \atari2600.cpu.inc ;
 wire \atari2600.cpu.index_y ;
 wire \atari2600.cpu.load_only ;
 wire \atari2600.cpu.load_reg ;
 wire \atari2600.cpu.op[0] ;
 wire \atari2600.cpu.op[1] ;
 wire \atari2600.cpu.op[2] ;
 wire \atari2600.cpu.op[3] ;
 wire \atari2600.cpu.php ;
 wire \atari2600.cpu.plp ;
 wire \atari2600.cpu.res ;
 wire \atari2600.cpu.rotate ;
 wire \atari2600.cpu.sec ;
 wire \atari2600.cpu.sed ;
 wire \atari2600.cpu.sei ;
 wire \atari2600.cpu.shift ;
 wire \atari2600.cpu.shift_right ;
 wire \atari2600.cpu.src_reg[0] ;
 wire \atari2600.cpu.src_reg[1] ;
 wire \atari2600.cpu.state[0] ;
 wire \atari2600.cpu.state[1] ;
 wire \atari2600.cpu.state[2] ;
 wire \atari2600.cpu.state[3] ;
 wire \atari2600.cpu.state[4] ;
 wire \atari2600.cpu.state[5] ;
 wire \atari2600.cpu.store ;
 wire \atari2600.cpu.write_back ;
 wire \atari2600.input_switches[0] ;
 wire \atari2600.input_switches[1] ;
 wire \atari2600.input_switches[2] ;
 wire \atari2600.input_switches[3] ;
 wire \atari2600.pia.dat_o[0] ;
 wire \atari2600.pia.dat_o[1] ;
 wire \atari2600.pia.dat_o[2] ;
 wire \atari2600.pia.dat_o[3] ;
 wire \atari2600.pia.dat_o[4] ;
 wire \atari2600.pia.dat_o[5] ;
 wire \atari2600.pia.dat_o[6] ;
 wire \atari2600.pia.dat_o[7] ;
 wire \atari2600.pia.diag[0] ;
 wire \atari2600.pia.diag[1] ;
 wire \atari2600.pia.diag[2] ;
 wire \atari2600.pia.diag[3] ;
 wire \atari2600.pia.diag[4] ;
 wire \atari2600.pia.diag[5] ;
 wire \atari2600.pia.diag[6] ;
 wire \atari2600.pia.diag[7] ;
 wire \atari2600.pia.instat[0] ;
 wire \atari2600.pia.instat[1] ;
 wire \atari2600.pia.interval[0] ;
 wire \atari2600.pia.interval[10] ;
 wire \atari2600.pia.interval[3] ;
 wire \atari2600.pia.interval[6] ;
 wire \atari2600.pia.reset_timer[0] ;
 wire \atari2600.pia.reset_timer[1] ;
 wire \atari2600.pia.reset_timer[2] ;
 wire \atari2600.pia.reset_timer[3] ;
 wire \atari2600.pia.reset_timer[4] ;
 wire \atari2600.pia.reset_timer[5] ;
 wire \atari2600.pia.reset_timer[6] ;
 wire \atari2600.pia.reset_timer[7] ;
 wire \atari2600.pia.swa_dir[0] ;
 wire \atari2600.pia.swa_dir[1] ;
 wire \atari2600.pia.swa_dir[2] ;
 wire \atari2600.pia.swa_dir[3] ;
 wire \atari2600.pia.swa_dir[4] ;
 wire \atari2600.pia.swa_dir[5] ;
 wire \atari2600.pia.swa_dir[6] ;
 wire \atari2600.pia.swa_dir[7] ;
 wire \atari2600.pia.swb_dir[2] ;
 wire \atari2600.pia.swb_dir[4] ;
 wire \atari2600.pia.swb_dir[5] ;
 wire \atari2600.pia.time_counter[0] ;
 wire \atari2600.pia.time_counter[10] ;
 wire \atari2600.pia.time_counter[11] ;
 wire \atari2600.pia.time_counter[12] ;
 wire \atari2600.pia.time_counter[13] ;
 wire \atari2600.pia.time_counter[14] ;
 wire \atari2600.pia.time_counter[15] ;
 wire \atari2600.pia.time_counter[16] ;
 wire \atari2600.pia.time_counter[17] ;
 wire \atari2600.pia.time_counter[18] ;
 wire \atari2600.pia.time_counter[19] ;
 wire \atari2600.pia.time_counter[1] ;
 wire \atari2600.pia.time_counter[20] ;
 wire \atari2600.pia.time_counter[21] ;
 wire \atari2600.pia.time_counter[22] ;
 wire \atari2600.pia.time_counter[23] ;
 wire \atari2600.pia.time_counter[2] ;
 wire \atari2600.pia.time_counter[3] ;
 wire \atari2600.pia.time_counter[4] ;
 wire \atari2600.pia.time_counter[5] ;
 wire \atari2600.pia.time_counter[6] ;
 wire \atari2600.pia.time_counter[7] ;
 wire \atari2600.pia.time_counter[8] ;
 wire \atari2600.pia.time_counter[9] ;
 wire \atari2600.pia.underflow ;
 wire \atari2600.ram[0][0] ;
 wire \atari2600.ram[0][1] ;
 wire \atari2600.ram[0][2] ;
 wire \atari2600.ram[0][3] ;
 wire \atari2600.ram[0][4] ;
 wire \atari2600.ram[0][5] ;
 wire \atari2600.ram[0][6] ;
 wire \atari2600.ram[0][7] ;
 wire \atari2600.ram[100][0] ;
 wire \atari2600.ram[100][1] ;
 wire \atari2600.ram[100][2] ;
 wire \atari2600.ram[100][3] ;
 wire \atari2600.ram[100][4] ;
 wire \atari2600.ram[100][5] ;
 wire \atari2600.ram[100][6] ;
 wire \atari2600.ram[100][7] ;
 wire \atari2600.ram[101][0] ;
 wire \atari2600.ram[101][1] ;
 wire \atari2600.ram[101][2] ;
 wire \atari2600.ram[101][3] ;
 wire \atari2600.ram[101][4] ;
 wire \atari2600.ram[101][5] ;
 wire \atari2600.ram[101][6] ;
 wire \atari2600.ram[101][7] ;
 wire \atari2600.ram[102][0] ;
 wire \atari2600.ram[102][1] ;
 wire \atari2600.ram[102][2] ;
 wire \atari2600.ram[102][3] ;
 wire \atari2600.ram[102][4] ;
 wire \atari2600.ram[102][5] ;
 wire \atari2600.ram[102][6] ;
 wire \atari2600.ram[102][7] ;
 wire \atari2600.ram[103][0] ;
 wire \atari2600.ram[103][1] ;
 wire \atari2600.ram[103][2] ;
 wire \atari2600.ram[103][3] ;
 wire \atari2600.ram[103][4] ;
 wire \atari2600.ram[103][5] ;
 wire \atari2600.ram[103][6] ;
 wire \atari2600.ram[103][7] ;
 wire \atari2600.ram[104][0] ;
 wire \atari2600.ram[104][1] ;
 wire \atari2600.ram[104][2] ;
 wire \atari2600.ram[104][3] ;
 wire \atari2600.ram[104][4] ;
 wire \atari2600.ram[104][5] ;
 wire \atari2600.ram[104][6] ;
 wire \atari2600.ram[104][7] ;
 wire \atari2600.ram[105][0] ;
 wire \atari2600.ram[105][1] ;
 wire \atari2600.ram[105][2] ;
 wire \atari2600.ram[105][3] ;
 wire \atari2600.ram[105][4] ;
 wire \atari2600.ram[105][5] ;
 wire \atari2600.ram[105][6] ;
 wire \atari2600.ram[105][7] ;
 wire \atari2600.ram[106][0] ;
 wire \atari2600.ram[106][1] ;
 wire \atari2600.ram[106][2] ;
 wire \atari2600.ram[106][3] ;
 wire \atari2600.ram[106][4] ;
 wire \atari2600.ram[106][5] ;
 wire \atari2600.ram[106][6] ;
 wire \atari2600.ram[106][7] ;
 wire \atari2600.ram[107][0] ;
 wire \atari2600.ram[107][1] ;
 wire \atari2600.ram[107][2] ;
 wire \atari2600.ram[107][3] ;
 wire \atari2600.ram[107][4] ;
 wire \atari2600.ram[107][5] ;
 wire \atari2600.ram[107][6] ;
 wire \atari2600.ram[107][7] ;
 wire \atari2600.ram[108][0] ;
 wire \atari2600.ram[108][1] ;
 wire \atari2600.ram[108][2] ;
 wire \atari2600.ram[108][3] ;
 wire \atari2600.ram[108][4] ;
 wire \atari2600.ram[108][5] ;
 wire \atari2600.ram[108][6] ;
 wire \atari2600.ram[108][7] ;
 wire \atari2600.ram[109][0] ;
 wire \atari2600.ram[109][1] ;
 wire \atari2600.ram[109][2] ;
 wire \atari2600.ram[109][3] ;
 wire \atari2600.ram[109][4] ;
 wire \atari2600.ram[109][5] ;
 wire \atari2600.ram[109][6] ;
 wire \atari2600.ram[109][7] ;
 wire \atari2600.ram[10][0] ;
 wire \atari2600.ram[10][1] ;
 wire \atari2600.ram[10][2] ;
 wire \atari2600.ram[10][3] ;
 wire \atari2600.ram[10][4] ;
 wire \atari2600.ram[10][5] ;
 wire \atari2600.ram[10][6] ;
 wire \atari2600.ram[10][7] ;
 wire \atari2600.ram[110][0] ;
 wire \atari2600.ram[110][1] ;
 wire \atari2600.ram[110][2] ;
 wire \atari2600.ram[110][3] ;
 wire \atari2600.ram[110][4] ;
 wire \atari2600.ram[110][5] ;
 wire \atari2600.ram[110][6] ;
 wire \atari2600.ram[110][7] ;
 wire \atari2600.ram[111][0] ;
 wire \atari2600.ram[111][1] ;
 wire \atari2600.ram[111][2] ;
 wire \atari2600.ram[111][3] ;
 wire \atari2600.ram[111][4] ;
 wire \atari2600.ram[111][5] ;
 wire \atari2600.ram[111][6] ;
 wire \atari2600.ram[111][7] ;
 wire \atari2600.ram[112][0] ;
 wire \atari2600.ram[112][1] ;
 wire \atari2600.ram[112][2] ;
 wire \atari2600.ram[112][3] ;
 wire \atari2600.ram[112][4] ;
 wire \atari2600.ram[112][5] ;
 wire \atari2600.ram[112][6] ;
 wire \atari2600.ram[112][7] ;
 wire \atari2600.ram[113][0] ;
 wire \atari2600.ram[113][1] ;
 wire \atari2600.ram[113][2] ;
 wire \atari2600.ram[113][3] ;
 wire \atari2600.ram[113][4] ;
 wire \atari2600.ram[113][5] ;
 wire \atari2600.ram[113][6] ;
 wire \atari2600.ram[113][7] ;
 wire \atari2600.ram[114][0] ;
 wire \atari2600.ram[114][1] ;
 wire \atari2600.ram[114][2] ;
 wire \atari2600.ram[114][3] ;
 wire \atari2600.ram[114][4] ;
 wire \atari2600.ram[114][5] ;
 wire \atari2600.ram[114][6] ;
 wire \atari2600.ram[114][7] ;
 wire \atari2600.ram[115][0] ;
 wire \atari2600.ram[115][1] ;
 wire \atari2600.ram[115][2] ;
 wire \atari2600.ram[115][3] ;
 wire \atari2600.ram[115][4] ;
 wire \atari2600.ram[115][5] ;
 wire \atari2600.ram[115][6] ;
 wire \atari2600.ram[115][7] ;
 wire \atari2600.ram[116][0] ;
 wire \atari2600.ram[116][1] ;
 wire \atari2600.ram[116][2] ;
 wire \atari2600.ram[116][3] ;
 wire \atari2600.ram[116][4] ;
 wire \atari2600.ram[116][5] ;
 wire \atari2600.ram[116][6] ;
 wire \atari2600.ram[116][7] ;
 wire \atari2600.ram[117][0] ;
 wire \atari2600.ram[117][1] ;
 wire \atari2600.ram[117][2] ;
 wire \atari2600.ram[117][3] ;
 wire \atari2600.ram[117][4] ;
 wire \atari2600.ram[117][5] ;
 wire \atari2600.ram[117][6] ;
 wire \atari2600.ram[117][7] ;
 wire \atari2600.ram[118][0] ;
 wire \atari2600.ram[118][1] ;
 wire \atari2600.ram[118][2] ;
 wire \atari2600.ram[118][3] ;
 wire \atari2600.ram[118][4] ;
 wire \atari2600.ram[118][5] ;
 wire \atari2600.ram[118][6] ;
 wire \atari2600.ram[118][7] ;
 wire \atari2600.ram[119][0] ;
 wire \atari2600.ram[119][1] ;
 wire \atari2600.ram[119][2] ;
 wire \atari2600.ram[119][3] ;
 wire \atari2600.ram[119][4] ;
 wire \atari2600.ram[119][5] ;
 wire \atari2600.ram[119][6] ;
 wire \atari2600.ram[119][7] ;
 wire \atari2600.ram[11][0] ;
 wire \atari2600.ram[11][1] ;
 wire \atari2600.ram[11][2] ;
 wire \atari2600.ram[11][3] ;
 wire \atari2600.ram[11][4] ;
 wire \atari2600.ram[11][5] ;
 wire \atari2600.ram[11][6] ;
 wire \atari2600.ram[11][7] ;
 wire \atari2600.ram[120][0] ;
 wire \atari2600.ram[120][1] ;
 wire \atari2600.ram[120][2] ;
 wire \atari2600.ram[120][3] ;
 wire \atari2600.ram[120][4] ;
 wire \atari2600.ram[120][5] ;
 wire \atari2600.ram[120][6] ;
 wire \atari2600.ram[120][7] ;
 wire \atari2600.ram[121][0] ;
 wire \atari2600.ram[121][1] ;
 wire \atari2600.ram[121][2] ;
 wire \atari2600.ram[121][3] ;
 wire \atari2600.ram[121][4] ;
 wire \atari2600.ram[121][5] ;
 wire \atari2600.ram[121][6] ;
 wire \atari2600.ram[121][7] ;
 wire \atari2600.ram[122][0] ;
 wire \atari2600.ram[122][1] ;
 wire \atari2600.ram[122][2] ;
 wire \atari2600.ram[122][3] ;
 wire \atari2600.ram[122][4] ;
 wire \atari2600.ram[122][5] ;
 wire \atari2600.ram[122][6] ;
 wire \atari2600.ram[122][7] ;
 wire \atari2600.ram[123][0] ;
 wire \atari2600.ram[123][1] ;
 wire \atari2600.ram[123][2] ;
 wire \atari2600.ram[123][3] ;
 wire \atari2600.ram[123][4] ;
 wire \atari2600.ram[123][5] ;
 wire \atari2600.ram[123][6] ;
 wire \atari2600.ram[123][7] ;
 wire \atari2600.ram[124][0] ;
 wire \atari2600.ram[124][1] ;
 wire \atari2600.ram[124][2] ;
 wire \atari2600.ram[124][3] ;
 wire \atari2600.ram[124][4] ;
 wire \atari2600.ram[124][5] ;
 wire \atari2600.ram[124][6] ;
 wire \atari2600.ram[124][7] ;
 wire \atari2600.ram[125][0] ;
 wire \atari2600.ram[125][1] ;
 wire \atari2600.ram[125][2] ;
 wire \atari2600.ram[125][3] ;
 wire \atari2600.ram[125][4] ;
 wire \atari2600.ram[125][5] ;
 wire \atari2600.ram[125][6] ;
 wire \atari2600.ram[125][7] ;
 wire \atari2600.ram[126][0] ;
 wire \atari2600.ram[126][1] ;
 wire \atari2600.ram[126][2] ;
 wire \atari2600.ram[126][3] ;
 wire \atari2600.ram[126][4] ;
 wire \atari2600.ram[126][5] ;
 wire \atari2600.ram[126][6] ;
 wire \atari2600.ram[126][7] ;
 wire \atari2600.ram[127][0] ;
 wire \atari2600.ram[127][1] ;
 wire \atari2600.ram[127][2] ;
 wire \atari2600.ram[127][3] ;
 wire \atari2600.ram[127][4] ;
 wire \atari2600.ram[127][5] ;
 wire \atari2600.ram[127][6] ;
 wire \atari2600.ram[127][7] ;
 wire \atari2600.ram[12][0] ;
 wire \atari2600.ram[12][1] ;
 wire \atari2600.ram[12][2] ;
 wire \atari2600.ram[12][3] ;
 wire \atari2600.ram[12][4] ;
 wire \atari2600.ram[12][5] ;
 wire \atari2600.ram[12][6] ;
 wire \atari2600.ram[12][7] ;
 wire \atari2600.ram[13][0] ;
 wire \atari2600.ram[13][1] ;
 wire \atari2600.ram[13][2] ;
 wire \atari2600.ram[13][3] ;
 wire \atari2600.ram[13][4] ;
 wire \atari2600.ram[13][5] ;
 wire \atari2600.ram[13][6] ;
 wire \atari2600.ram[13][7] ;
 wire \atari2600.ram[14][0] ;
 wire \atari2600.ram[14][1] ;
 wire \atari2600.ram[14][2] ;
 wire \atari2600.ram[14][3] ;
 wire \atari2600.ram[14][4] ;
 wire \atari2600.ram[14][5] ;
 wire \atari2600.ram[14][6] ;
 wire \atari2600.ram[14][7] ;
 wire \atari2600.ram[15][0] ;
 wire \atari2600.ram[15][1] ;
 wire \atari2600.ram[15][2] ;
 wire \atari2600.ram[15][3] ;
 wire \atari2600.ram[15][4] ;
 wire \atari2600.ram[15][5] ;
 wire \atari2600.ram[15][6] ;
 wire \atari2600.ram[15][7] ;
 wire \atari2600.ram[16][0] ;
 wire \atari2600.ram[16][1] ;
 wire \atari2600.ram[16][2] ;
 wire \atari2600.ram[16][3] ;
 wire \atari2600.ram[16][4] ;
 wire \atari2600.ram[16][5] ;
 wire \atari2600.ram[16][6] ;
 wire \atari2600.ram[16][7] ;
 wire \atari2600.ram[17][0] ;
 wire \atari2600.ram[17][1] ;
 wire \atari2600.ram[17][2] ;
 wire \atari2600.ram[17][3] ;
 wire \atari2600.ram[17][4] ;
 wire \atari2600.ram[17][5] ;
 wire \atari2600.ram[17][6] ;
 wire \atari2600.ram[17][7] ;
 wire \atari2600.ram[18][0] ;
 wire \atari2600.ram[18][1] ;
 wire \atari2600.ram[18][2] ;
 wire \atari2600.ram[18][3] ;
 wire \atari2600.ram[18][4] ;
 wire \atari2600.ram[18][5] ;
 wire \atari2600.ram[18][6] ;
 wire \atari2600.ram[18][7] ;
 wire \atari2600.ram[19][0] ;
 wire \atari2600.ram[19][1] ;
 wire \atari2600.ram[19][2] ;
 wire \atari2600.ram[19][3] ;
 wire \atari2600.ram[19][4] ;
 wire \atari2600.ram[19][5] ;
 wire \atari2600.ram[19][6] ;
 wire \atari2600.ram[19][7] ;
 wire \atari2600.ram[1][0] ;
 wire \atari2600.ram[1][1] ;
 wire \atari2600.ram[1][2] ;
 wire \atari2600.ram[1][3] ;
 wire \atari2600.ram[1][4] ;
 wire \atari2600.ram[1][5] ;
 wire \atari2600.ram[1][6] ;
 wire \atari2600.ram[1][7] ;
 wire \atari2600.ram[20][0] ;
 wire \atari2600.ram[20][1] ;
 wire \atari2600.ram[20][2] ;
 wire \atari2600.ram[20][3] ;
 wire \atari2600.ram[20][4] ;
 wire \atari2600.ram[20][5] ;
 wire \atari2600.ram[20][6] ;
 wire \atari2600.ram[20][7] ;
 wire \atari2600.ram[21][0] ;
 wire \atari2600.ram[21][1] ;
 wire \atari2600.ram[21][2] ;
 wire \atari2600.ram[21][3] ;
 wire \atari2600.ram[21][4] ;
 wire \atari2600.ram[21][5] ;
 wire \atari2600.ram[21][6] ;
 wire \atari2600.ram[21][7] ;
 wire \atari2600.ram[22][0] ;
 wire \atari2600.ram[22][1] ;
 wire \atari2600.ram[22][2] ;
 wire \atari2600.ram[22][3] ;
 wire \atari2600.ram[22][4] ;
 wire \atari2600.ram[22][5] ;
 wire \atari2600.ram[22][6] ;
 wire \atari2600.ram[22][7] ;
 wire \atari2600.ram[23][0] ;
 wire \atari2600.ram[23][1] ;
 wire \atari2600.ram[23][2] ;
 wire \atari2600.ram[23][3] ;
 wire \atari2600.ram[23][4] ;
 wire \atari2600.ram[23][5] ;
 wire \atari2600.ram[23][6] ;
 wire \atari2600.ram[23][7] ;
 wire \atari2600.ram[24][0] ;
 wire \atari2600.ram[24][1] ;
 wire \atari2600.ram[24][2] ;
 wire \atari2600.ram[24][3] ;
 wire \atari2600.ram[24][4] ;
 wire \atari2600.ram[24][5] ;
 wire \atari2600.ram[24][6] ;
 wire \atari2600.ram[24][7] ;
 wire \atari2600.ram[25][0] ;
 wire \atari2600.ram[25][1] ;
 wire \atari2600.ram[25][2] ;
 wire \atari2600.ram[25][3] ;
 wire \atari2600.ram[25][4] ;
 wire \atari2600.ram[25][5] ;
 wire \atari2600.ram[25][6] ;
 wire \atari2600.ram[25][7] ;
 wire \atari2600.ram[26][0] ;
 wire \atari2600.ram[26][1] ;
 wire \atari2600.ram[26][2] ;
 wire \atari2600.ram[26][3] ;
 wire \atari2600.ram[26][4] ;
 wire \atari2600.ram[26][5] ;
 wire \atari2600.ram[26][6] ;
 wire \atari2600.ram[26][7] ;
 wire \atari2600.ram[27][0] ;
 wire \atari2600.ram[27][1] ;
 wire \atari2600.ram[27][2] ;
 wire \atari2600.ram[27][3] ;
 wire \atari2600.ram[27][4] ;
 wire \atari2600.ram[27][5] ;
 wire \atari2600.ram[27][6] ;
 wire \atari2600.ram[27][7] ;
 wire \atari2600.ram[28][0] ;
 wire \atari2600.ram[28][1] ;
 wire \atari2600.ram[28][2] ;
 wire \atari2600.ram[28][3] ;
 wire \atari2600.ram[28][4] ;
 wire \atari2600.ram[28][5] ;
 wire \atari2600.ram[28][6] ;
 wire \atari2600.ram[28][7] ;
 wire \atari2600.ram[29][0] ;
 wire \atari2600.ram[29][1] ;
 wire \atari2600.ram[29][2] ;
 wire \atari2600.ram[29][3] ;
 wire \atari2600.ram[29][4] ;
 wire \atari2600.ram[29][5] ;
 wire \atari2600.ram[29][6] ;
 wire \atari2600.ram[29][7] ;
 wire \atari2600.ram[2][0] ;
 wire \atari2600.ram[2][1] ;
 wire \atari2600.ram[2][2] ;
 wire \atari2600.ram[2][3] ;
 wire \atari2600.ram[2][4] ;
 wire \atari2600.ram[2][5] ;
 wire \atari2600.ram[2][6] ;
 wire \atari2600.ram[2][7] ;
 wire \atari2600.ram[30][0] ;
 wire \atari2600.ram[30][1] ;
 wire \atari2600.ram[30][2] ;
 wire \atari2600.ram[30][3] ;
 wire \atari2600.ram[30][4] ;
 wire \atari2600.ram[30][5] ;
 wire \atari2600.ram[30][6] ;
 wire \atari2600.ram[30][7] ;
 wire \atari2600.ram[31][0] ;
 wire \atari2600.ram[31][1] ;
 wire \atari2600.ram[31][2] ;
 wire \atari2600.ram[31][3] ;
 wire \atari2600.ram[31][4] ;
 wire \atari2600.ram[31][5] ;
 wire \atari2600.ram[31][6] ;
 wire \atari2600.ram[31][7] ;
 wire \atari2600.ram[32][0] ;
 wire \atari2600.ram[32][1] ;
 wire \atari2600.ram[32][2] ;
 wire \atari2600.ram[32][3] ;
 wire \atari2600.ram[32][4] ;
 wire \atari2600.ram[32][5] ;
 wire \atari2600.ram[32][6] ;
 wire \atari2600.ram[32][7] ;
 wire \atari2600.ram[33][0] ;
 wire \atari2600.ram[33][1] ;
 wire \atari2600.ram[33][2] ;
 wire \atari2600.ram[33][3] ;
 wire \atari2600.ram[33][4] ;
 wire \atari2600.ram[33][5] ;
 wire \atari2600.ram[33][6] ;
 wire \atari2600.ram[33][7] ;
 wire \atari2600.ram[34][0] ;
 wire \atari2600.ram[34][1] ;
 wire \atari2600.ram[34][2] ;
 wire \atari2600.ram[34][3] ;
 wire \atari2600.ram[34][4] ;
 wire \atari2600.ram[34][5] ;
 wire \atari2600.ram[34][6] ;
 wire \atari2600.ram[34][7] ;
 wire \atari2600.ram[35][0] ;
 wire \atari2600.ram[35][1] ;
 wire \atari2600.ram[35][2] ;
 wire \atari2600.ram[35][3] ;
 wire \atari2600.ram[35][4] ;
 wire \atari2600.ram[35][5] ;
 wire \atari2600.ram[35][6] ;
 wire \atari2600.ram[35][7] ;
 wire \atari2600.ram[36][0] ;
 wire \atari2600.ram[36][1] ;
 wire \atari2600.ram[36][2] ;
 wire \atari2600.ram[36][3] ;
 wire \atari2600.ram[36][4] ;
 wire \atari2600.ram[36][5] ;
 wire \atari2600.ram[36][6] ;
 wire \atari2600.ram[36][7] ;
 wire \atari2600.ram[37][0] ;
 wire \atari2600.ram[37][1] ;
 wire \atari2600.ram[37][2] ;
 wire \atari2600.ram[37][3] ;
 wire \atari2600.ram[37][4] ;
 wire \atari2600.ram[37][5] ;
 wire \atari2600.ram[37][6] ;
 wire \atari2600.ram[37][7] ;
 wire \atari2600.ram[38][0] ;
 wire \atari2600.ram[38][1] ;
 wire \atari2600.ram[38][2] ;
 wire \atari2600.ram[38][3] ;
 wire \atari2600.ram[38][4] ;
 wire \atari2600.ram[38][5] ;
 wire \atari2600.ram[38][6] ;
 wire \atari2600.ram[38][7] ;
 wire \atari2600.ram[39][0] ;
 wire \atari2600.ram[39][1] ;
 wire \atari2600.ram[39][2] ;
 wire \atari2600.ram[39][3] ;
 wire \atari2600.ram[39][4] ;
 wire \atari2600.ram[39][5] ;
 wire \atari2600.ram[39][6] ;
 wire \atari2600.ram[39][7] ;
 wire \atari2600.ram[3][0] ;
 wire \atari2600.ram[3][1] ;
 wire \atari2600.ram[3][2] ;
 wire \atari2600.ram[3][3] ;
 wire \atari2600.ram[3][4] ;
 wire \atari2600.ram[3][5] ;
 wire \atari2600.ram[3][6] ;
 wire \atari2600.ram[3][7] ;
 wire \atari2600.ram[40][0] ;
 wire \atari2600.ram[40][1] ;
 wire \atari2600.ram[40][2] ;
 wire \atari2600.ram[40][3] ;
 wire \atari2600.ram[40][4] ;
 wire \atari2600.ram[40][5] ;
 wire \atari2600.ram[40][6] ;
 wire \atari2600.ram[40][7] ;
 wire \atari2600.ram[41][0] ;
 wire \atari2600.ram[41][1] ;
 wire \atari2600.ram[41][2] ;
 wire \atari2600.ram[41][3] ;
 wire \atari2600.ram[41][4] ;
 wire \atari2600.ram[41][5] ;
 wire \atari2600.ram[41][6] ;
 wire \atari2600.ram[41][7] ;
 wire \atari2600.ram[42][0] ;
 wire \atari2600.ram[42][1] ;
 wire \atari2600.ram[42][2] ;
 wire \atari2600.ram[42][3] ;
 wire \atari2600.ram[42][4] ;
 wire \atari2600.ram[42][5] ;
 wire \atari2600.ram[42][6] ;
 wire \atari2600.ram[42][7] ;
 wire \atari2600.ram[43][0] ;
 wire \atari2600.ram[43][1] ;
 wire \atari2600.ram[43][2] ;
 wire \atari2600.ram[43][3] ;
 wire \atari2600.ram[43][4] ;
 wire \atari2600.ram[43][5] ;
 wire \atari2600.ram[43][6] ;
 wire \atari2600.ram[43][7] ;
 wire \atari2600.ram[44][0] ;
 wire \atari2600.ram[44][1] ;
 wire \atari2600.ram[44][2] ;
 wire \atari2600.ram[44][3] ;
 wire \atari2600.ram[44][4] ;
 wire \atari2600.ram[44][5] ;
 wire \atari2600.ram[44][6] ;
 wire \atari2600.ram[44][7] ;
 wire \atari2600.ram[45][0] ;
 wire \atari2600.ram[45][1] ;
 wire \atari2600.ram[45][2] ;
 wire \atari2600.ram[45][3] ;
 wire \atari2600.ram[45][4] ;
 wire \atari2600.ram[45][5] ;
 wire \atari2600.ram[45][6] ;
 wire \atari2600.ram[45][7] ;
 wire \atari2600.ram[46][0] ;
 wire \atari2600.ram[46][1] ;
 wire \atari2600.ram[46][2] ;
 wire \atari2600.ram[46][3] ;
 wire \atari2600.ram[46][4] ;
 wire \atari2600.ram[46][5] ;
 wire \atari2600.ram[46][6] ;
 wire \atari2600.ram[46][7] ;
 wire \atari2600.ram[47][0] ;
 wire \atari2600.ram[47][1] ;
 wire \atari2600.ram[47][2] ;
 wire \atari2600.ram[47][3] ;
 wire \atari2600.ram[47][4] ;
 wire \atari2600.ram[47][5] ;
 wire \atari2600.ram[47][6] ;
 wire \atari2600.ram[47][7] ;
 wire \atari2600.ram[48][0] ;
 wire \atari2600.ram[48][1] ;
 wire \atari2600.ram[48][2] ;
 wire \atari2600.ram[48][3] ;
 wire \atari2600.ram[48][4] ;
 wire \atari2600.ram[48][5] ;
 wire \atari2600.ram[48][6] ;
 wire \atari2600.ram[48][7] ;
 wire \atari2600.ram[49][0] ;
 wire \atari2600.ram[49][1] ;
 wire \atari2600.ram[49][2] ;
 wire \atari2600.ram[49][3] ;
 wire \atari2600.ram[49][4] ;
 wire \atari2600.ram[49][5] ;
 wire \atari2600.ram[49][6] ;
 wire \atari2600.ram[49][7] ;
 wire \atari2600.ram[4][0] ;
 wire \atari2600.ram[4][1] ;
 wire \atari2600.ram[4][2] ;
 wire \atari2600.ram[4][3] ;
 wire \atari2600.ram[4][4] ;
 wire \atari2600.ram[4][5] ;
 wire \atari2600.ram[4][6] ;
 wire \atari2600.ram[4][7] ;
 wire \atari2600.ram[50][0] ;
 wire \atari2600.ram[50][1] ;
 wire \atari2600.ram[50][2] ;
 wire \atari2600.ram[50][3] ;
 wire \atari2600.ram[50][4] ;
 wire \atari2600.ram[50][5] ;
 wire \atari2600.ram[50][6] ;
 wire \atari2600.ram[50][7] ;
 wire \atari2600.ram[51][0] ;
 wire \atari2600.ram[51][1] ;
 wire \atari2600.ram[51][2] ;
 wire \atari2600.ram[51][3] ;
 wire \atari2600.ram[51][4] ;
 wire \atari2600.ram[51][5] ;
 wire \atari2600.ram[51][6] ;
 wire \atari2600.ram[51][7] ;
 wire \atari2600.ram[52][0] ;
 wire \atari2600.ram[52][1] ;
 wire \atari2600.ram[52][2] ;
 wire \atari2600.ram[52][3] ;
 wire \atari2600.ram[52][4] ;
 wire \atari2600.ram[52][5] ;
 wire \atari2600.ram[52][6] ;
 wire \atari2600.ram[52][7] ;
 wire \atari2600.ram[53][0] ;
 wire \atari2600.ram[53][1] ;
 wire \atari2600.ram[53][2] ;
 wire \atari2600.ram[53][3] ;
 wire \atari2600.ram[53][4] ;
 wire \atari2600.ram[53][5] ;
 wire \atari2600.ram[53][6] ;
 wire \atari2600.ram[53][7] ;
 wire \atari2600.ram[54][0] ;
 wire \atari2600.ram[54][1] ;
 wire \atari2600.ram[54][2] ;
 wire \atari2600.ram[54][3] ;
 wire \atari2600.ram[54][4] ;
 wire \atari2600.ram[54][5] ;
 wire \atari2600.ram[54][6] ;
 wire \atari2600.ram[54][7] ;
 wire \atari2600.ram[55][0] ;
 wire \atari2600.ram[55][1] ;
 wire \atari2600.ram[55][2] ;
 wire \atari2600.ram[55][3] ;
 wire \atari2600.ram[55][4] ;
 wire \atari2600.ram[55][5] ;
 wire \atari2600.ram[55][6] ;
 wire \atari2600.ram[55][7] ;
 wire \atari2600.ram[56][0] ;
 wire \atari2600.ram[56][1] ;
 wire \atari2600.ram[56][2] ;
 wire \atari2600.ram[56][3] ;
 wire \atari2600.ram[56][4] ;
 wire \atari2600.ram[56][5] ;
 wire \atari2600.ram[56][6] ;
 wire \atari2600.ram[56][7] ;
 wire \atari2600.ram[57][0] ;
 wire \atari2600.ram[57][1] ;
 wire \atari2600.ram[57][2] ;
 wire \atari2600.ram[57][3] ;
 wire \atari2600.ram[57][4] ;
 wire \atari2600.ram[57][5] ;
 wire \atari2600.ram[57][6] ;
 wire \atari2600.ram[57][7] ;
 wire \atari2600.ram[58][0] ;
 wire \atari2600.ram[58][1] ;
 wire \atari2600.ram[58][2] ;
 wire \atari2600.ram[58][3] ;
 wire \atari2600.ram[58][4] ;
 wire \atari2600.ram[58][5] ;
 wire \atari2600.ram[58][6] ;
 wire \atari2600.ram[58][7] ;
 wire \atari2600.ram[59][0] ;
 wire \atari2600.ram[59][1] ;
 wire \atari2600.ram[59][2] ;
 wire \atari2600.ram[59][3] ;
 wire \atari2600.ram[59][4] ;
 wire \atari2600.ram[59][5] ;
 wire \atari2600.ram[59][6] ;
 wire \atari2600.ram[59][7] ;
 wire \atari2600.ram[5][0] ;
 wire \atari2600.ram[5][1] ;
 wire \atari2600.ram[5][2] ;
 wire \atari2600.ram[5][3] ;
 wire \atari2600.ram[5][4] ;
 wire \atari2600.ram[5][5] ;
 wire \atari2600.ram[5][6] ;
 wire \atari2600.ram[5][7] ;
 wire \atari2600.ram[60][0] ;
 wire \atari2600.ram[60][1] ;
 wire \atari2600.ram[60][2] ;
 wire \atari2600.ram[60][3] ;
 wire \atari2600.ram[60][4] ;
 wire \atari2600.ram[60][5] ;
 wire \atari2600.ram[60][6] ;
 wire \atari2600.ram[60][7] ;
 wire \atari2600.ram[61][0] ;
 wire \atari2600.ram[61][1] ;
 wire \atari2600.ram[61][2] ;
 wire \atari2600.ram[61][3] ;
 wire \atari2600.ram[61][4] ;
 wire \atari2600.ram[61][5] ;
 wire \atari2600.ram[61][6] ;
 wire \atari2600.ram[61][7] ;
 wire \atari2600.ram[62][0] ;
 wire \atari2600.ram[62][1] ;
 wire \atari2600.ram[62][2] ;
 wire \atari2600.ram[62][3] ;
 wire \atari2600.ram[62][4] ;
 wire \atari2600.ram[62][5] ;
 wire \atari2600.ram[62][6] ;
 wire \atari2600.ram[62][7] ;
 wire \atari2600.ram[63][0] ;
 wire \atari2600.ram[63][1] ;
 wire \atari2600.ram[63][2] ;
 wire \atari2600.ram[63][3] ;
 wire \atari2600.ram[63][4] ;
 wire \atari2600.ram[63][5] ;
 wire \atari2600.ram[63][6] ;
 wire \atari2600.ram[63][7] ;
 wire \atari2600.ram[64][0] ;
 wire \atari2600.ram[64][1] ;
 wire \atari2600.ram[64][2] ;
 wire \atari2600.ram[64][3] ;
 wire \atari2600.ram[64][4] ;
 wire \atari2600.ram[64][5] ;
 wire \atari2600.ram[64][6] ;
 wire \atari2600.ram[64][7] ;
 wire \atari2600.ram[65][0] ;
 wire \atari2600.ram[65][1] ;
 wire \atari2600.ram[65][2] ;
 wire \atari2600.ram[65][3] ;
 wire \atari2600.ram[65][4] ;
 wire \atari2600.ram[65][5] ;
 wire \atari2600.ram[65][6] ;
 wire \atari2600.ram[65][7] ;
 wire \atari2600.ram[66][0] ;
 wire \atari2600.ram[66][1] ;
 wire \atari2600.ram[66][2] ;
 wire \atari2600.ram[66][3] ;
 wire \atari2600.ram[66][4] ;
 wire \atari2600.ram[66][5] ;
 wire \atari2600.ram[66][6] ;
 wire \atari2600.ram[66][7] ;
 wire \atari2600.ram[67][0] ;
 wire \atari2600.ram[67][1] ;
 wire \atari2600.ram[67][2] ;
 wire \atari2600.ram[67][3] ;
 wire \atari2600.ram[67][4] ;
 wire \atari2600.ram[67][5] ;
 wire \atari2600.ram[67][6] ;
 wire \atari2600.ram[67][7] ;
 wire \atari2600.ram[68][0] ;
 wire \atari2600.ram[68][1] ;
 wire \atari2600.ram[68][2] ;
 wire \atari2600.ram[68][3] ;
 wire \atari2600.ram[68][4] ;
 wire \atari2600.ram[68][5] ;
 wire \atari2600.ram[68][6] ;
 wire \atari2600.ram[68][7] ;
 wire \atari2600.ram[69][0] ;
 wire \atari2600.ram[69][1] ;
 wire \atari2600.ram[69][2] ;
 wire \atari2600.ram[69][3] ;
 wire \atari2600.ram[69][4] ;
 wire \atari2600.ram[69][5] ;
 wire \atari2600.ram[69][6] ;
 wire \atari2600.ram[69][7] ;
 wire \atari2600.ram[6][0] ;
 wire \atari2600.ram[6][1] ;
 wire \atari2600.ram[6][2] ;
 wire \atari2600.ram[6][3] ;
 wire \atari2600.ram[6][4] ;
 wire \atari2600.ram[6][5] ;
 wire \atari2600.ram[6][6] ;
 wire \atari2600.ram[6][7] ;
 wire \atari2600.ram[70][0] ;
 wire \atari2600.ram[70][1] ;
 wire \atari2600.ram[70][2] ;
 wire \atari2600.ram[70][3] ;
 wire \atari2600.ram[70][4] ;
 wire \atari2600.ram[70][5] ;
 wire \atari2600.ram[70][6] ;
 wire \atari2600.ram[70][7] ;
 wire \atari2600.ram[71][0] ;
 wire \atari2600.ram[71][1] ;
 wire \atari2600.ram[71][2] ;
 wire \atari2600.ram[71][3] ;
 wire \atari2600.ram[71][4] ;
 wire \atari2600.ram[71][5] ;
 wire \atari2600.ram[71][6] ;
 wire \atari2600.ram[71][7] ;
 wire \atari2600.ram[72][0] ;
 wire \atari2600.ram[72][1] ;
 wire \atari2600.ram[72][2] ;
 wire \atari2600.ram[72][3] ;
 wire \atari2600.ram[72][4] ;
 wire \atari2600.ram[72][5] ;
 wire \atari2600.ram[72][6] ;
 wire \atari2600.ram[72][7] ;
 wire \atari2600.ram[73][0] ;
 wire \atari2600.ram[73][1] ;
 wire \atari2600.ram[73][2] ;
 wire \atari2600.ram[73][3] ;
 wire \atari2600.ram[73][4] ;
 wire \atari2600.ram[73][5] ;
 wire \atari2600.ram[73][6] ;
 wire \atari2600.ram[73][7] ;
 wire \atari2600.ram[74][0] ;
 wire \atari2600.ram[74][1] ;
 wire \atari2600.ram[74][2] ;
 wire \atari2600.ram[74][3] ;
 wire \atari2600.ram[74][4] ;
 wire \atari2600.ram[74][5] ;
 wire \atari2600.ram[74][6] ;
 wire \atari2600.ram[74][7] ;
 wire \atari2600.ram[75][0] ;
 wire \atari2600.ram[75][1] ;
 wire \atari2600.ram[75][2] ;
 wire \atari2600.ram[75][3] ;
 wire \atari2600.ram[75][4] ;
 wire \atari2600.ram[75][5] ;
 wire \atari2600.ram[75][6] ;
 wire \atari2600.ram[75][7] ;
 wire \atari2600.ram[76][0] ;
 wire \atari2600.ram[76][1] ;
 wire \atari2600.ram[76][2] ;
 wire \atari2600.ram[76][3] ;
 wire \atari2600.ram[76][4] ;
 wire \atari2600.ram[76][5] ;
 wire \atari2600.ram[76][6] ;
 wire \atari2600.ram[76][7] ;
 wire \atari2600.ram[77][0] ;
 wire \atari2600.ram[77][1] ;
 wire \atari2600.ram[77][2] ;
 wire \atari2600.ram[77][3] ;
 wire \atari2600.ram[77][4] ;
 wire \atari2600.ram[77][5] ;
 wire \atari2600.ram[77][6] ;
 wire \atari2600.ram[77][7] ;
 wire \atari2600.ram[78][0] ;
 wire \atari2600.ram[78][1] ;
 wire \atari2600.ram[78][2] ;
 wire \atari2600.ram[78][3] ;
 wire \atari2600.ram[78][4] ;
 wire \atari2600.ram[78][5] ;
 wire \atari2600.ram[78][6] ;
 wire \atari2600.ram[78][7] ;
 wire \atari2600.ram[79][0] ;
 wire \atari2600.ram[79][1] ;
 wire \atari2600.ram[79][2] ;
 wire \atari2600.ram[79][3] ;
 wire \atari2600.ram[79][4] ;
 wire \atari2600.ram[79][5] ;
 wire \atari2600.ram[79][6] ;
 wire \atari2600.ram[79][7] ;
 wire \atari2600.ram[7][0] ;
 wire \atari2600.ram[7][1] ;
 wire \atari2600.ram[7][2] ;
 wire \atari2600.ram[7][3] ;
 wire \atari2600.ram[7][4] ;
 wire \atari2600.ram[7][5] ;
 wire \atari2600.ram[7][6] ;
 wire \atari2600.ram[7][7] ;
 wire \atari2600.ram[80][0] ;
 wire \atari2600.ram[80][1] ;
 wire \atari2600.ram[80][2] ;
 wire \atari2600.ram[80][3] ;
 wire \atari2600.ram[80][4] ;
 wire \atari2600.ram[80][5] ;
 wire \atari2600.ram[80][6] ;
 wire \atari2600.ram[80][7] ;
 wire \atari2600.ram[81][0] ;
 wire \atari2600.ram[81][1] ;
 wire \atari2600.ram[81][2] ;
 wire \atari2600.ram[81][3] ;
 wire \atari2600.ram[81][4] ;
 wire \atari2600.ram[81][5] ;
 wire \atari2600.ram[81][6] ;
 wire \atari2600.ram[81][7] ;
 wire \atari2600.ram[82][0] ;
 wire \atari2600.ram[82][1] ;
 wire \atari2600.ram[82][2] ;
 wire \atari2600.ram[82][3] ;
 wire \atari2600.ram[82][4] ;
 wire \atari2600.ram[82][5] ;
 wire \atari2600.ram[82][6] ;
 wire \atari2600.ram[82][7] ;
 wire \atari2600.ram[83][0] ;
 wire \atari2600.ram[83][1] ;
 wire \atari2600.ram[83][2] ;
 wire \atari2600.ram[83][3] ;
 wire \atari2600.ram[83][4] ;
 wire \atari2600.ram[83][5] ;
 wire \atari2600.ram[83][6] ;
 wire \atari2600.ram[83][7] ;
 wire \atari2600.ram[84][0] ;
 wire \atari2600.ram[84][1] ;
 wire \atari2600.ram[84][2] ;
 wire \atari2600.ram[84][3] ;
 wire \atari2600.ram[84][4] ;
 wire \atari2600.ram[84][5] ;
 wire \atari2600.ram[84][6] ;
 wire \atari2600.ram[84][7] ;
 wire \atari2600.ram[85][0] ;
 wire \atari2600.ram[85][1] ;
 wire \atari2600.ram[85][2] ;
 wire \atari2600.ram[85][3] ;
 wire \atari2600.ram[85][4] ;
 wire \atari2600.ram[85][5] ;
 wire \atari2600.ram[85][6] ;
 wire \atari2600.ram[85][7] ;
 wire \atari2600.ram[86][0] ;
 wire \atari2600.ram[86][1] ;
 wire \atari2600.ram[86][2] ;
 wire \atari2600.ram[86][3] ;
 wire \atari2600.ram[86][4] ;
 wire \atari2600.ram[86][5] ;
 wire \atari2600.ram[86][6] ;
 wire \atari2600.ram[86][7] ;
 wire \atari2600.ram[87][0] ;
 wire \atari2600.ram[87][1] ;
 wire \atari2600.ram[87][2] ;
 wire \atari2600.ram[87][3] ;
 wire \atari2600.ram[87][4] ;
 wire \atari2600.ram[87][5] ;
 wire \atari2600.ram[87][6] ;
 wire \atari2600.ram[87][7] ;
 wire \atari2600.ram[88][0] ;
 wire \atari2600.ram[88][1] ;
 wire \atari2600.ram[88][2] ;
 wire \atari2600.ram[88][3] ;
 wire \atari2600.ram[88][4] ;
 wire \atari2600.ram[88][5] ;
 wire \atari2600.ram[88][6] ;
 wire \atari2600.ram[88][7] ;
 wire \atari2600.ram[89][0] ;
 wire \atari2600.ram[89][1] ;
 wire \atari2600.ram[89][2] ;
 wire \atari2600.ram[89][3] ;
 wire \atari2600.ram[89][4] ;
 wire \atari2600.ram[89][5] ;
 wire \atari2600.ram[89][6] ;
 wire \atari2600.ram[89][7] ;
 wire \atari2600.ram[8][0] ;
 wire \atari2600.ram[8][1] ;
 wire \atari2600.ram[8][2] ;
 wire \atari2600.ram[8][3] ;
 wire \atari2600.ram[8][4] ;
 wire \atari2600.ram[8][5] ;
 wire \atari2600.ram[8][6] ;
 wire \atari2600.ram[8][7] ;
 wire \atari2600.ram[90][0] ;
 wire \atari2600.ram[90][1] ;
 wire \atari2600.ram[90][2] ;
 wire \atari2600.ram[90][3] ;
 wire \atari2600.ram[90][4] ;
 wire \atari2600.ram[90][5] ;
 wire \atari2600.ram[90][6] ;
 wire \atari2600.ram[90][7] ;
 wire \atari2600.ram[91][0] ;
 wire \atari2600.ram[91][1] ;
 wire \atari2600.ram[91][2] ;
 wire \atari2600.ram[91][3] ;
 wire \atari2600.ram[91][4] ;
 wire \atari2600.ram[91][5] ;
 wire \atari2600.ram[91][6] ;
 wire \atari2600.ram[91][7] ;
 wire \atari2600.ram[92][0] ;
 wire \atari2600.ram[92][1] ;
 wire \atari2600.ram[92][2] ;
 wire \atari2600.ram[92][3] ;
 wire \atari2600.ram[92][4] ;
 wire \atari2600.ram[92][5] ;
 wire \atari2600.ram[92][6] ;
 wire \atari2600.ram[92][7] ;
 wire \atari2600.ram[93][0] ;
 wire \atari2600.ram[93][1] ;
 wire \atari2600.ram[93][2] ;
 wire \atari2600.ram[93][3] ;
 wire \atari2600.ram[93][4] ;
 wire \atari2600.ram[93][5] ;
 wire \atari2600.ram[93][6] ;
 wire \atari2600.ram[93][7] ;
 wire \atari2600.ram[94][0] ;
 wire \atari2600.ram[94][1] ;
 wire \atari2600.ram[94][2] ;
 wire \atari2600.ram[94][3] ;
 wire \atari2600.ram[94][4] ;
 wire \atari2600.ram[94][5] ;
 wire \atari2600.ram[94][6] ;
 wire \atari2600.ram[94][7] ;
 wire \atari2600.ram[95][0] ;
 wire \atari2600.ram[95][1] ;
 wire \atari2600.ram[95][2] ;
 wire \atari2600.ram[95][3] ;
 wire \atari2600.ram[95][4] ;
 wire \atari2600.ram[95][5] ;
 wire \atari2600.ram[95][6] ;
 wire \atari2600.ram[95][7] ;
 wire \atari2600.ram[96][0] ;
 wire \atari2600.ram[96][1] ;
 wire \atari2600.ram[96][2] ;
 wire \atari2600.ram[96][3] ;
 wire \atari2600.ram[96][4] ;
 wire \atari2600.ram[96][5] ;
 wire \atari2600.ram[96][6] ;
 wire \atari2600.ram[96][7] ;
 wire \atari2600.ram[97][0] ;
 wire \atari2600.ram[97][1] ;
 wire \atari2600.ram[97][2] ;
 wire \atari2600.ram[97][3] ;
 wire \atari2600.ram[97][4] ;
 wire \atari2600.ram[97][5] ;
 wire \atari2600.ram[97][6] ;
 wire \atari2600.ram[97][7] ;
 wire \atari2600.ram[98][0] ;
 wire \atari2600.ram[98][1] ;
 wire \atari2600.ram[98][2] ;
 wire \atari2600.ram[98][3] ;
 wire \atari2600.ram[98][4] ;
 wire \atari2600.ram[98][5] ;
 wire \atari2600.ram[98][6] ;
 wire \atari2600.ram[98][7] ;
 wire \atari2600.ram[99][0] ;
 wire \atari2600.ram[99][1] ;
 wire \atari2600.ram[99][2] ;
 wire \atari2600.ram[99][3] ;
 wire \atari2600.ram[99][4] ;
 wire \atari2600.ram[99][5] ;
 wire \atari2600.ram[99][6] ;
 wire \atari2600.ram[99][7] ;
 wire \atari2600.ram[9][0] ;
 wire \atari2600.ram[9][1] ;
 wire \atari2600.ram[9][2] ;
 wire \atari2600.ram[9][3] ;
 wire \atari2600.ram[9][4] ;
 wire \atari2600.ram[9][5] ;
 wire \atari2600.ram[9][6] ;
 wire \atari2600.ram[9][7] ;
 wire \atari2600.ram_data[0] ;
 wire \atari2600.ram_data[1] ;
 wire \atari2600.ram_data[2] ;
 wire \atari2600.ram_data[3] ;
 wire \atari2600.ram_data[4] ;
 wire \atari2600.ram_data[5] ;
 wire \atari2600.ram_data[6] ;
 wire \atari2600.ram_data[7] ;
 wire \atari2600.stall_cpu ;
 wire \atari2600.tia.audc0[0] ;
 wire \atari2600.tia.audc0[1] ;
 wire \atari2600.tia.audc0[2] ;
 wire \atari2600.tia.audc0[3] ;
 wire \atari2600.tia.audc1[0] ;
 wire \atari2600.tia.audc1[1] ;
 wire \atari2600.tia.audc1[2] ;
 wire \atari2600.tia.audc1[3] ;
 wire \atari2600.tia.audf0[0] ;
 wire \atari2600.tia.audf0[1] ;
 wire \atari2600.tia.audf0[2] ;
 wire \atari2600.tia.audf0[3] ;
 wire \atari2600.tia.audf0[4] ;
 wire \atari2600.tia.audf1[0] ;
 wire \atari2600.tia.audf1[1] ;
 wire \atari2600.tia.audf1[2] ;
 wire \atari2600.tia.audf1[3] ;
 wire \atari2600.tia.audf1[4] ;
 wire \atari2600.tia.audio_l ;
 wire \atari2600.tia.audio_left_counter[0] ;
 wire \atari2600.tia.audio_left_counter[10] ;
 wire \atari2600.tia.audio_left_counter[11] ;
 wire \atari2600.tia.audio_left_counter[12] ;
 wire \atari2600.tia.audio_left_counter[13] ;
 wire \atari2600.tia.audio_left_counter[14] ;
 wire \atari2600.tia.audio_left_counter[15] ;
 wire \atari2600.tia.audio_left_counter[1] ;
 wire \atari2600.tia.audio_left_counter[2] ;
 wire \atari2600.tia.audio_left_counter[3] ;
 wire \atari2600.tia.audio_left_counter[4] ;
 wire \atari2600.tia.audio_left_counter[5] ;
 wire \atari2600.tia.audio_left_counter[6] ;
 wire \atari2600.tia.audio_left_counter[7] ;
 wire \atari2600.tia.audio_left_counter[8] ;
 wire \atari2600.tia.audio_left_counter[9] ;
 wire \atari2600.tia.audio_r ;
 wire \atari2600.tia.audio_right_counter[0] ;
 wire \atari2600.tia.audio_right_counter[10] ;
 wire \atari2600.tia.audio_right_counter[11] ;
 wire \atari2600.tia.audio_right_counter[12] ;
 wire \atari2600.tia.audio_right_counter[13] ;
 wire \atari2600.tia.audio_right_counter[14] ;
 wire \atari2600.tia.audio_right_counter[15] ;
 wire \atari2600.tia.audio_right_counter[1] ;
 wire \atari2600.tia.audio_right_counter[2] ;
 wire \atari2600.tia.audio_right_counter[3] ;
 wire \atari2600.tia.audio_right_counter[4] ;
 wire \atari2600.tia.audio_right_counter[5] ;
 wire \atari2600.tia.audio_right_counter[6] ;
 wire \atari2600.tia.audio_right_counter[7] ;
 wire \atari2600.tia.audio_right_counter[8] ;
 wire \atari2600.tia.audio_right_counter[9] ;
 wire \atari2600.tia.audv0[0] ;
 wire \atari2600.tia.audv0[1] ;
 wire \atari2600.tia.audv0[2] ;
 wire \atari2600.tia.audv0[3] ;
 wire \atari2600.tia.audv1[0] ;
 wire \atari2600.tia.audv1[1] ;
 wire \atari2600.tia.audv1[2] ;
 wire \atari2600.tia.audv1[3] ;
 wire \atari2600.tia.ball_w[0] ;
 wire \atari2600.tia.ball_w[1] ;
 wire \atari2600.tia.ball_w[2] ;
 wire \atari2600.tia.ball_w[3] ;
 wire \atari2600.tia.colubk[0] ;
 wire \atari2600.tia.colubk[1] ;
 wire \atari2600.tia.colubk[2] ;
 wire \atari2600.tia.colubk[3] ;
 wire \atari2600.tia.colubk[4] ;
 wire \atari2600.tia.colubk[5] ;
 wire \atari2600.tia.colubk[6] ;
 wire \atari2600.tia.colup0[0] ;
 wire \atari2600.tia.colup0[1] ;
 wire \atari2600.tia.colup0[2] ;
 wire \atari2600.tia.colup0[3] ;
 wire \atari2600.tia.colup0[4] ;
 wire \atari2600.tia.colup0[5] ;
 wire \atari2600.tia.colup0[6] ;
 wire \atari2600.tia.colup1[0] ;
 wire \atari2600.tia.colup1[1] ;
 wire \atari2600.tia.colup1[2] ;
 wire \atari2600.tia.colup1[3] ;
 wire \atari2600.tia.colup1[4] ;
 wire \atari2600.tia.colup1[5] ;
 wire \atari2600.tia.colup1[6] ;
 wire \atari2600.tia.colupf[0] ;
 wire \atari2600.tia.colupf[1] ;
 wire \atari2600.tia.colupf[2] ;
 wire \atari2600.tia.colupf[3] ;
 wire \atari2600.tia.colupf[4] ;
 wire \atari2600.tia.colupf[5] ;
 wire \atari2600.tia.colupf[6] ;
 wire \atari2600.tia.cx[0] ;
 wire \atari2600.tia.cx[10] ;
 wire \atari2600.tia.cx[11] ;
 wire \atari2600.tia.cx[12] ;
 wire \atari2600.tia.cx[13] ;
 wire \atari2600.tia.cx[14] ;
 wire \atari2600.tia.cx[1] ;
 wire \atari2600.tia.cx[2] ;
 wire \atari2600.tia.cx[3] ;
 wire \atari2600.tia.cx[4] ;
 wire \atari2600.tia.cx[5] ;
 wire \atari2600.tia.cx[6] ;
 wire \atari2600.tia.cx[7] ;
 wire \atari2600.tia.cx[8] ;
 wire \atari2600.tia.cx[9] ;
 wire \atari2600.tia.cx_clr ;
 wire \atari2600.tia.dat_o[6] ;
 wire \atari2600.tia.dat_o[7] ;
 wire \atari2600.tia.diag[100] ;
 wire \atari2600.tia.diag[101] ;
 wire \atari2600.tia.diag[102] ;
 wire \atari2600.tia.diag[103] ;
 wire \atari2600.tia.diag[104] ;
 wire \atari2600.tia.diag[105] ;
 wire \atari2600.tia.diag[106] ;
 wire \atari2600.tia.diag[107] ;
 wire \atari2600.tia.diag[108] ;
 wire \atari2600.tia.diag[109] ;
 wire \atari2600.tia.diag[110] ;
 wire \atari2600.tia.diag[111] ;
 wire \atari2600.tia.diag[32] ;
 wire \atari2600.tia.diag[33] ;
 wire \atari2600.tia.diag[34] ;
 wire \atari2600.tia.diag[35] ;
 wire \atari2600.tia.diag[36] ;
 wire \atari2600.tia.diag[37] ;
 wire \atari2600.tia.diag[38] ;
 wire \atari2600.tia.diag[39] ;
 wire \atari2600.tia.diag[40] ;
 wire \atari2600.tia.diag[41] ;
 wire \atari2600.tia.diag[42] ;
 wire \atari2600.tia.diag[43] ;
 wire \atari2600.tia.diag[44] ;
 wire \atari2600.tia.diag[45] ;
 wire \atari2600.tia.diag[46] ;
 wire \atari2600.tia.diag[47] ;
 wire \atari2600.tia.diag[48] ;
 wire \atari2600.tia.diag[49] ;
 wire \atari2600.tia.diag[50] ;
 wire \atari2600.tia.diag[51] ;
 wire \atari2600.tia.diag[52] ;
 wire \atari2600.tia.diag[53] ;
 wire \atari2600.tia.diag[54] ;
 wire \atari2600.tia.diag[55] ;
 wire \atari2600.tia.diag[56] ;
 wire \atari2600.tia.diag[57] ;
 wire \atari2600.tia.diag[58] ;
 wire \atari2600.tia.diag[59] ;
 wire \atari2600.tia.diag[60] ;
 wire \atari2600.tia.diag[61] ;
 wire \atari2600.tia.diag[62] ;
 wire \atari2600.tia.diag[63] ;
 wire \atari2600.tia.diag[64] ;
 wire \atari2600.tia.diag[65] ;
 wire \atari2600.tia.diag[66] ;
 wire \atari2600.tia.diag[67] ;
 wire \atari2600.tia.diag[68] ;
 wire \atari2600.tia.diag[69] ;
 wire \atari2600.tia.diag[70] ;
 wire \atari2600.tia.diag[71] ;
 wire \atari2600.tia.diag[76] ;
 wire \atari2600.tia.diag[77] ;
 wire \atari2600.tia.diag[78] ;
 wire \atari2600.tia.diag[79] ;
 wire \atari2600.tia.diag[80] ;
 wire \atari2600.tia.diag[81] ;
 wire \atari2600.tia.diag[82] ;
 wire \atari2600.tia.diag[83] ;
 wire \atari2600.tia.diag[84] ;
 wire \atari2600.tia.diag[85] ;
 wire \atari2600.tia.diag[86] ;
 wire \atari2600.tia.diag[87] ;
 wire \atari2600.tia.diag[88] ;
 wire \atari2600.tia.diag[89] ;
 wire \atari2600.tia.diag[90] ;
 wire \atari2600.tia.diag[91] ;
 wire \atari2600.tia.diag[92] ;
 wire \atari2600.tia.diag[93] ;
 wire \atari2600.tia.diag[94] ;
 wire \atari2600.tia.diag[95] ;
 wire \atari2600.tia.diag[96] ;
 wire \atari2600.tia.diag[97] ;
 wire \atari2600.tia.diag[98] ;
 wire \atari2600.tia.diag[99] ;
 wire \atari2600.tia.enabl ;
 wire \atari2600.tia.enam0 ;
 wire \atari2600.tia.enam1 ;
 wire \atari2600.tia.hmbl[0] ;
 wire \atari2600.tia.hmbl[1] ;
 wire \atari2600.tia.hmbl[2] ;
 wire \atari2600.tia.hmbl[3] ;
 wire \atari2600.tia.hmm0[0] ;
 wire \atari2600.tia.hmm0[1] ;
 wire \atari2600.tia.hmm0[2] ;
 wire \atari2600.tia.hmm0[3] ;
 wire \atari2600.tia.hmm1[0] ;
 wire \atari2600.tia.hmm1[1] ;
 wire \atari2600.tia.hmm1[2] ;
 wire \atari2600.tia.hmm1[3] ;
 wire \atari2600.tia.hmp0[0] ;
 wire \atari2600.tia.hmp0[1] ;
 wire \atari2600.tia.hmp0[2] ;
 wire \atari2600.tia.hmp0[3] ;
 wire \atari2600.tia.hmp1[0] ;
 wire \atari2600.tia.hmp1[1] ;
 wire \atari2600.tia.hmp1[2] ;
 wire \atari2600.tia.hmp1[3] ;
 wire \atari2600.tia.m0_w[0] ;
 wire \atari2600.tia.m0_w[1] ;
 wire \atari2600.tia.m0_w[2] ;
 wire \atari2600.tia.m0_w[3] ;
 wire \atari2600.tia.m1_w[0] ;
 wire \atari2600.tia.m1_w[1] ;
 wire \atari2600.tia.m1_w[2] ;
 wire \atari2600.tia.m1_w[3] ;
 wire \atari2600.tia.old_grp0[0] ;
 wire \atari2600.tia.old_grp0[1] ;
 wire \atari2600.tia.old_grp0[2] ;
 wire \atari2600.tia.old_grp0[3] ;
 wire \atari2600.tia.old_grp0[4] ;
 wire \atari2600.tia.old_grp0[5] ;
 wire \atari2600.tia.old_grp0[6] ;
 wire \atari2600.tia.old_grp0[7] ;
 wire \atari2600.tia.old_grp1[0] ;
 wire \atari2600.tia.old_grp1[1] ;
 wire \atari2600.tia.old_grp1[2] ;
 wire \atari2600.tia.old_grp1[3] ;
 wire \atari2600.tia.old_grp1[4] ;
 wire \atari2600.tia.old_grp1[5] ;
 wire \atari2600.tia.old_grp1[6] ;
 wire \atari2600.tia.old_grp1[7] ;
 wire \atari2600.tia.p0_copies[1] ;
 wire \atari2600.tia.p0_copies[2] ;
 wire \atari2600.tia.p0_scale[0] ;
 wire \atari2600.tia.p0_scale[1] ;
 wire \atari2600.tia.p0_spacing[4] ;
 wire \atari2600.tia.p0_spacing[5] ;
 wire \atari2600.tia.p0_spacing[6] ;
 wire \atari2600.tia.p0_w[3] ;
 wire \atari2600.tia.p0_w[4] ;
 wire \atari2600.tia.p0_w[5] ;
 wire \atari2600.tia.p1_copies[1] ;
 wire \atari2600.tia.p1_copies[2] ;
 wire \atari2600.tia.p1_scale[0] ;
 wire \atari2600.tia.p1_scale[1] ;
 wire \atari2600.tia.p1_spacing[4] ;
 wire \atari2600.tia.p1_spacing[5] ;
 wire \atari2600.tia.p1_spacing[6] ;
 wire \atari2600.tia.p1_w[3] ;
 wire \atari2600.tia.p1_w[4] ;
 wire \atari2600.tia.p1_w[5] ;
 wire \atari2600.tia.p4_l ;
 wire \atari2600.tia.p4_r ;
 wire \atari2600.tia.p5_l ;
 wire \atari2600.tia.p5_r ;
 wire \atari2600.tia.p9_l ;
 wire \atari2600.tia.p9_r ;
 wire \atari2600.tia.pf_priority ;
 wire \atari2600.tia.poly4_l.x[1] ;
 wire \atari2600.tia.poly4_l.x[2] ;
 wire \atari2600.tia.poly4_l.x[3] ;
 wire \atari2600.tia.poly4_r.x[1] ;
 wire \atari2600.tia.poly4_r.x[2] ;
 wire \atari2600.tia.poly4_r.x[3] ;
 wire \atari2600.tia.poly5_l.x[1] ;
 wire \atari2600.tia.poly5_l.x[2] ;
 wire \atari2600.tia.poly5_l.x[3] ;
 wire \atari2600.tia.poly5_l.x[4] ;
 wire \atari2600.tia.poly5_r.x[1] ;
 wire \atari2600.tia.poly5_r.x[2] ;
 wire \atari2600.tia.poly5_r.x[3] ;
 wire \atari2600.tia.poly5_r.x[4] ;
 wire \atari2600.tia.poly9_l.x[1] ;
 wire \atari2600.tia.poly9_l.x[2] ;
 wire \atari2600.tia.poly9_l.x[3] ;
 wire \atari2600.tia.poly9_l.x[4] ;
 wire \atari2600.tia.poly9_l.x[5] ;
 wire \atari2600.tia.poly9_l.x[6] ;
 wire \atari2600.tia.poly9_l.x[7] ;
 wire \atari2600.tia.poly9_l.x[8] ;
 wire \atari2600.tia.poly9_r.x[1] ;
 wire \atari2600.tia.poly9_r.x[2] ;
 wire \atari2600.tia.poly9_r.x[3] ;
 wire \atari2600.tia.poly9_r.x[4] ;
 wire \atari2600.tia.poly9_r.x[5] ;
 wire \atari2600.tia.poly9_r.x[6] ;
 wire \atari2600.tia.poly9_r.x[7] ;
 wire \atari2600.tia.poly9_r.x[8] ;
 wire \atari2600.tia.refp0 ;
 wire \atari2600.tia.refp1 ;
 wire \atari2600.tia.refpf ;
 wire \atari2600.tia.scorepf ;
 wire \atari2600.tia.vblank ;
 wire \atari2600.tia.vdelp0 ;
 wire \atari2600.tia.vdelp1 ;
 wire \atari2600.tia.vid_out[0] ;
 wire \atari2600.tia.vid_out[1] ;
 wire \atari2600.tia.vid_out[2] ;
 wire \atari2600.tia.vid_out[3] ;
 wire \atari2600.tia.vid_out[4] ;
 wire \atari2600.tia.vid_out[5] ;
 wire \atari2600.tia.vid_out[6] ;
 wire \atari2600.tia.vid_vsync ;
 wire \atari2600.tia.vid_xpos[0] ;
 wire \atari2600.tia.vid_xpos[1] ;
 wire \atari2600.tia.vid_xpos[2] ;
 wire \atari2600.tia.vid_xpos[3] ;
 wire \atari2600.tia.vid_xpos[4] ;
 wire \atari2600.tia.vid_xpos[5] ;
 wire \atari2600.tia.vid_xpos[6] ;
 wire \atari2600.tia.vid_xpos[7] ;
 wire \atari2600.tia.vid_ypos[0] ;
 wire \atari2600.tia.vid_ypos[1] ;
 wire \atari2600.tia.vid_ypos[2] ;
 wire \atari2600.tia.vid_ypos[3] ;
 wire \atari2600.tia.vid_ypos[4] ;
 wire \atari2600.tia.vid_ypos[5] ;
 wire \atari2600.tia.vid_ypos[6] ;
 wire \atari2600.tia.vid_ypos[7] ;
 wire \atari2600.tia.vid_ypos[8] ;
 wire audio_pwm;
 wire \audio_pwm_accumulator[0] ;
 wire \audio_pwm_accumulator[1] ;
 wire \audio_pwm_accumulator[2] ;
 wire \audio_pwm_accumulator[3] ;
 wire \audio_pwm_accumulator[4] ;
 wire \b_pwm_even[1] ;
 wire \b_pwm_even[2] ;
 wire \b_pwm_even[3] ;
 wire \b_pwm_even[4] ;
 wire \b_pwm_even[5] ;
 wire \b_pwm_even[6] ;
 wire \b_pwm_even[7] ;
 wire \b_pwm_even[8] ;
 wire \b_pwm_even[9] ;
 wire \b_pwm_odd[1] ;
 wire \b_pwm_odd[2] ;
 wire \b_pwm_odd[3] ;
 wire \b_pwm_odd[4] ;
 wire \b_pwm_odd[5] ;
 wire \b_pwm_odd[6] ;
 wire \b_pwm_odd[7] ;
 wire \b_pwm_odd[8] ;
 wire \b_pwm_odd[9] ;
 wire \external_rom_data[0] ;
 wire \external_rom_data[1] ;
 wire \external_rom_data[2] ;
 wire \external_rom_data[3] ;
 wire \external_rom_data[4] ;
 wire \external_rom_data[5] ;
 wire \external_rom_data[6] ;
 wire \external_rom_data[7] ;
 wire \flash_rom.addr[0] ;
 wire \flash_rom.addr[10] ;
 wire \flash_rom.addr[11] ;
 wire \flash_rom.addr[12] ;
 wire \flash_rom.addr[13] ;
 wire \flash_rom.addr[14] ;
 wire \flash_rom.addr[15] ;
 wire \flash_rom.addr[16] ;
 wire \flash_rom.addr[17] ;
 wire \flash_rom.addr[18] ;
 wire \flash_rom.addr[19] ;
 wire \flash_rom.addr[1] ;
 wire \flash_rom.addr[20] ;
 wire \flash_rom.addr[21] ;
 wire \flash_rom.addr[22] ;
 wire \flash_rom.addr[23] ;
 wire \flash_rom.addr[2] ;
 wire \flash_rom.addr[3] ;
 wire \flash_rom.addr[4] ;
 wire \flash_rom.addr[5] ;
 wire \flash_rom.addr[6] ;
 wire \flash_rom.addr[7] ;
 wire \flash_rom.addr[8] ;
 wire \flash_rom.addr[9] ;
 wire \flash_rom.addr_in[16] ;
 wire \flash_rom.addr_in[17] ;
 wire \flash_rom.addr_in[18] ;
 wire \flash_rom.addr_in[19] ;
 wire \flash_rom.data_ready ;
 wire \flash_rom.fsm_state[0] ;
 wire \flash_rom.fsm_state[1] ;
 wire \flash_rom.fsm_state[2] ;
 wire \flash_rom.nibbles_remaining[0] ;
 wire \flash_rom.nibbles_remaining[1] ;
 wire \flash_rom.nibbles_remaining[2] ;
 wire \flash_rom.spi_clk_out ;
 wire \flash_rom.spi_select ;
 wire \flash_rom.stall_read ;
 wire \frame_counter[0] ;
 wire \frame_counter[1] ;
 wire \frame_counter[2] ;
 wire \g_pwm_even[1] ;
 wire \g_pwm_even[2] ;
 wire \g_pwm_even[3] ;
 wire \g_pwm_even[4] ;
 wire \g_pwm_even[5] ;
 wire \g_pwm_even[6] ;
 wire \g_pwm_even[7] ;
 wire \g_pwm_even[8] ;
 wire \g_pwm_even[9] ;
 wire \g_pwm_odd[1] ;
 wire \g_pwm_odd[2] ;
 wire \g_pwm_odd[3] ;
 wire \g_pwm_odd[4] ;
 wire \g_pwm_odd[5] ;
 wire \g_pwm_odd[6] ;
 wire \g_pwm_odd[7] ;
 wire \g_pwm_odd[8] ;
 wire \g_pwm_odd[9] ;
 wire \gamepad_pmod.decoder.data_reg[0] ;
 wire \gamepad_pmod.decoder.data_reg[10] ;
 wire \gamepad_pmod.decoder.data_reg[11] ;
 wire \gamepad_pmod.decoder.data_reg[1] ;
 wire \gamepad_pmod.decoder.data_reg[2] ;
 wire \gamepad_pmod.decoder.data_reg[3] ;
 wire \gamepad_pmod.decoder.data_reg[4] ;
 wire \gamepad_pmod.decoder.data_reg[5] ;
 wire \gamepad_pmod.decoder.data_reg[6] ;
 wire \gamepad_pmod.decoder.data_reg[7] ;
 wire \gamepad_pmod.decoder.data_reg[8] ;
 wire \gamepad_pmod.decoder.data_reg[9] ;
 wire \gamepad_pmod.driver.pmod_clk_prev ;
 wire \gamepad_pmod.driver.pmod_clk_sync[0] ;
 wire \gamepad_pmod.driver.pmod_clk_sync[1] ;
 wire \gamepad_pmod.driver.pmod_data_sync[0] ;
 wire \gamepad_pmod.driver.pmod_data_sync[1] ;
 wire \gamepad_pmod.driver.pmod_latch_prev ;
 wire \gamepad_pmod.driver.pmod_latch_sync[0] ;
 wire \gamepad_pmod.driver.pmod_latch_sync[1] ;
 wire \gamepad_pmod.driver.shift_reg[0] ;
 wire \gamepad_pmod.driver.shift_reg[10] ;
 wire \gamepad_pmod.driver.shift_reg[11] ;
 wire \gamepad_pmod.driver.shift_reg[1] ;
 wire \gamepad_pmod.driver.shift_reg[2] ;
 wire \gamepad_pmod.driver.shift_reg[3] ;
 wire \gamepad_pmod.driver.shift_reg[4] ;
 wire \gamepad_pmod.driver.shift_reg[5] ;
 wire \gamepad_pmod.driver.shift_reg[6] ;
 wire \gamepad_pmod.driver.shift_reg[7] ;
 wire \gamepad_pmod.driver.shift_reg[8] ;
 wire \gamepad_pmod.driver.shift_reg[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vga.vpos[0] ;
 wire \hvsync_gen.vga.vpos[1] ;
 wire \hvsync_gen.vga.vpos[2] ;
 wire \hvsync_gen.vga.vpos[3] ;
 wire \hvsync_gen.vga.vpos[4] ;
 wire \hvsync_gen.vga.vpos[5] ;
 wire \hvsync_gen.vga.vpos[6] ;
 wire \hvsync_gen.vga.vpos[7] ;
 wire \hvsync_gen.vga.vpos[8] ;
 wire \hvsync_gen.vga.vpos[9] ;
 wire \hvsync_gen.vga.vsync ;
 wire \internal_rom_data[0] ;
 wire \internal_rom_data[1] ;
 wire \internal_rom_data[2] ;
 wire \internal_rom_data[3] ;
 wire \internal_rom_data[4] ;
 wire \internal_rom_data[5] ;
 wire \internal_rom_data[6] ;
 wire \internal_rom_data[7] ;
 wire \r_pwm_even[1] ;
 wire \r_pwm_even[2] ;
 wire \r_pwm_even[3] ;
 wire \r_pwm_even[4] ;
 wire \r_pwm_even[5] ;
 wire \r_pwm_even[6] ;
 wire \r_pwm_even[7] ;
 wire \r_pwm_even[8] ;
 wire \r_pwm_even[9] ;
 wire \r_pwm_odd[1] ;
 wire \r_pwm_odd[2] ;
 wire \r_pwm_odd[3] ;
 wire \r_pwm_odd[4] ;
 wire \r_pwm_odd[5] ;
 wire \r_pwm_odd[6] ;
 wire \r_pwm_odd[7] ;
 wire \r_pwm_odd[8] ;
 wire \r_pwm_odd[9] ;
 wire rom_data_pending;
 wire \rom_last_read_addr[0] ;
 wire \rom_last_read_addr[10] ;
 wire \rom_last_read_addr[11] ;
 wire \rom_last_read_addr[1] ;
 wire \rom_last_read_addr[2] ;
 wire \rom_last_read_addr[3] ;
 wire \rom_last_read_addr[4] ;
 wire \rom_last_read_addr[5] ;
 wire \rom_last_read_addr[6] ;
 wire \rom_last_read_addr[7] ;
 wire \rom_last_read_addr[8] ;
 wire \rom_last_read_addr[9] ;
 wire \rom_next_addr_in_queue[0] ;
 wire \rom_next_addr_in_queue[10] ;
 wire \rom_next_addr_in_queue[11] ;
 wire \rom_next_addr_in_queue[1] ;
 wire \rom_next_addr_in_queue[2] ;
 wire \rom_next_addr_in_queue[3] ;
 wire \rom_next_addr_in_queue[4] ;
 wire \rom_next_addr_in_queue[5] ;
 wire \rom_next_addr_in_queue[6] ;
 wire \rom_next_addr_in_queue[7] ;
 wire \rom_next_addr_in_queue[8] ;
 wire \rom_next_addr_in_queue[9] ;
 wire \scanline[0][0] ;
 wire \scanline[0][1] ;
 wire \scanline[0][2] ;
 wire \scanline[0][3] ;
 wire \scanline[0][4] ;
 wire \scanline[0][5] ;
 wire \scanline[0][6] ;
 wire \scanline[100][0] ;
 wire \scanline[100][1] ;
 wire \scanline[100][2] ;
 wire \scanline[100][3] ;
 wire \scanline[100][4] ;
 wire \scanline[100][5] ;
 wire \scanline[100][6] ;
 wire \scanline[101][0] ;
 wire \scanline[101][1] ;
 wire \scanline[101][2] ;
 wire \scanline[101][3] ;
 wire \scanline[101][4] ;
 wire \scanline[101][5] ;
 wire \scanline[101][6] ;
 wire \scanline[102][0] ;
 wire \scanline[102][1] ;
 wire \scanline[102][2] ;
 wire \scanline[102][3] ;
 wire \scanline[102][4] ;
 wire \scanline[102][5] ;
 wire \scanline[102][6] ;
 wire \scanline[103][0] ;
 wire \scanline[103][1] ;
 wire \scanline[103][2] ;
 wire \scanline[103][3] ;
 wire \scanline[103][4] ;
 wire \scanline[103][5] ;
 wire \scanline[103][6] ;
 wire \scanline[104][0] ;
 wire \scanline[104][1] ;
 wire \scanline[104][2] ;
 wire \scanline[104][3] ;
 wire \scanline[104][4] ;
 wire \scanline[104][5] ;
 wire \scanline[104][6] ;
 wire \scanline[105][0] ;
 wire \scanline[105][1] ;
 wire \scanline[105][2] ;
 wire \scanline[105][3] ;
 wire \scanline[105][4] ;
 wire \scanline[105][5] ;
 wire \scanline[105][6] ;
 wire \scanline[106][0] ;
 wire \scanline[106][1] ;
 wire \scanline[106][2] ;
 wire \scanline[106][3] ;
 wire \scanline[106][4] ;
 wire \scanline[106][5] ;
 wire \scanline[106][6] ;
 wire \scanline[107][0] ;
 wire \scanline[107][1] ;
 wire \scanline[107][2] ;
 wire \scanline[107][3] ;
 wire \scanline[107][4] ;
 wire \scanline[107][5] ;
 wire \scanline[107][6] ;
 wire \scanline[108][0] ;
 wire \scanline[108][1] ;
 wire \scanline[108][2] ;
 wire \scanline[108][3] ;
 wire \scanline[108][4] ;
 wire \scanline[108][5] ;
 wire \scanline[108][6] ;
 wire \scanline[109][0] ;
 wire \scanline[109][1] ;
 wire \scanline[109][2] ;
 wire \scanline[109][3] ;
 wire \scanline[109][4] ;
 wire \scanline[109][5] ;
 wire \scanline[109][6] ;
 wire \scanline[10][0] ;
 wire \scanline[10][1] ;
 wire \scanline[10][2] ;
 wire \scanline[10][3] ;
 wire \scanline[10][4] ;
 wire \scanline[10][5] ;
 wire \scanline[10][6] ;
 wire \scanline[110][0] ;
 wire \scanline[110][1] ;
 wire \scanline[110][2] ;
 wire \scanline[110][3] ;
 wire \scanline[110][4] ;
 wire \scanline[110][5] ;
 wire \scanline[110][6] ;
 wire \scanline[111][0] ;
 wire \scanline[111][1] ;
 wire \scanline[111][2] ;
 wire \scanline[111][3] ;
 wire \scanline[111][4] ;
 wire \scanline[111][5] ;
 wire \scanline[111][6] ;
 wire \scanline[112][0] ;
 wire \scanline[112][1] ;
 wire \scanline[112][2] ;
 wire \scanline[112][3] ;
 wire \scanline[112][4] ;
 wire \scanline[112][5] ;
 wire \scanline[112][6] ;
 wire \scanline[113][0] ;
 wire \scanline[113][1] ;
 wire \scanline[113][2] ;
 wire \scanline[113][3] ;
 wire \scanline[113][4] ;
 wire \scanline[113][5] ;
 wire \scanline[113][6] ;
 wire \scanline[114][0] ;
 wire \scanline[114][1] ;
 wire \scanline[114][2] ;
 wire \scanline[114][3] ;
 wire \scanline[114][4] ;
 wire \scanline[114][5] ;
 wire \scanline[114][6] ;
 wire \scanline[115][0] ;
 wire \scanline[115][1] ;
 wire \scanline[115][2] ;
 wire \scanline[115][3] ;
 wire \scanline[115][4] ;
 wire \scanline[115][5] ;
 wire \scanline[115][6] ;
 wire \scanline[116][0] ;
 wire \scanline[116][1] ;
 wire \scanline[116][2] ;
 wire \scanline[116][3] ;
 wire \scanline[116][4] ;
 wire \scanline[116][5] ;
 wire \scanline[116][6] ;
 wire \scanline[117][0] ;
 wire \scanline[117][1] ;
 wire \scanline[117][2] ;
 wire \scanline[117][3] ;
 wire \scanline[117][4] ;
 wire \scanline[117][5] ;
 wire \scanline[117][6] ;
 wire \scanline[118][0] ;
 wire \scanline[118][1] ;
 wire \scanline[118][2] ;
 wire \scanline[118][3] ;
 wire \scanline[118][4] ;
 wire \scanline[118][5] ;
 wire \scanline[118][6] ;
 wire \scanline[119][0] ;
 wire \scanline[119][1] ;
 wire \scanline[119][2] ;
 wire \scanline[119][3] ;
 wire \scanline[119][4] ;
 wire \scanline[119][5] ;
 wire \scanline[119][6] ;
 wire \scanline[11][0] ;
 wire \scanline[11][1] ;
 wire \scanline[11][2] ;
 wire \scanline[11][3] ;
 wire \scanline[11][4] ;
 wire \scanline[11][5] ;
 wire \scanline[11][6] ;
 wire \scanline[120][0] ;
 wire \scanline[120][1] ;
 wire \scanline[120][2] ;
 wire \scanline[120][3] ;
 wire \scanline[120][4] ;
 wire \scanline[120][5] ;
 wire \scanline[120][6] ;
 wire \scanline[121][0] ;
 wire \scanline[121][1] ;
 wire \scanline[121][2] ;
 wire \scanline[121][3] ;
 wire \scanline[121][4] ;
 wire \scanline[121][5] ;
 wire \scanline[121][6] ;
 wire \scanline[122][0] ;
 wire \scanline[122][1] ;
 wire \scanline[122][2] ;
 wire \scanline[122][3] ;
 wire \scanline[122][4] ;
 wire \scanline[122][5] ;
 wire \scanline[122][6] ;
 wire \scanline[123][0] ;
 wire \scanline[123][1] ;
 wire \scanline[123][2] ;
 wire \scanline[123][3] ;
 wire \scanline[123][4] ;
 wire \scanline[123][5] ;
 wire \scanline[123][6] ;
 wire \scanline[124][0] ;
 wire \scanline[124][1] ;
 wire \scanline[124][2] ;
 wire \scanline[124][3] ;
 wire \scanline[124][4] ;
 wire \scanline[124][5] ;
 wire \scanline[124][6] ;
 wire \scanline[125][0] ;
 wire \scanline[125][1] ;
 wire \scanline[125][2] ;
 wire \scanline[125][3] ;
 wire \scanline[125][4] ;
 wire \scanline[125][5] ;
 wire \scanline[125][6] ;
 wire \scanline[126][0] ;
 wire \scanline[126][1] ;
 wire \scanline[126][2] ;
 wire \scanline[126][3] ;
 wire \scanline[126][4] ;
 wire \scanline[126][5] ;
 wire \scanline[126][6] ;
 wire \scanline[127][0] ;
 wire \scanline[127][1] ;
 wire \scanline[127][2] ;
 wire \scanline[127][3] ;
 wire \scanline[127][4] ;
 wire \scanline[127][5] ;
 wire \scanline[127][6] ;
 wire \scanline[128][0] ;
 wire \scanline[128][1] ;
 wire \scanline[128][2] ;
 wire \scanline[128][3] ;
 wire \scanline[128][4] ;
 wire \scanline[128][5] ;
 wire \scanline[128][6] ;
 wire \scanline[129][0] ;
 wire \scanline[129][1] ;
 wire \scanline[129][2] ;
 wire \scanline[129][3] ;
 wire \scanline[129][4] ;
 wire \scanline[129][5] ;
 wire \scanline[129][6] ;
 wire \scanline[12][0] ;
 wire \scanline[12][1] ;
 wire \scanline[12][2] ;
 wire \scanline[12][3] ;
 wire \scanline[12][4] ;
 wire \scanline[12][5] ;
 wire \scanline[12][6] ;
 wire \scanline[130][0] ;
 wire \scanline[130][1] ;
 wire \scanline[130][2] ;
 wire \scanline[130][3] ;
 wire \scanline[130][4] ;
 wire \scanline[130][5] ;
 wire \scanline[130][6] ;
 wire \scanline[131][0] ;
 wire \scanline[131][1] ;
 wire \scanline[131][2] ;
 wire \scanline[131][3] ;
 wire \scanline[131][4] ;
 wire \scanline[131][5] ;
 wire \scanline[131][6] ;
 wire \scanline[132][0] ;
 wire \scanline[132][1] ;
 wire \scanline[132][2] ;
 wire \scanline[132][3] ;
 wire \scanline[132][4] ;
 wire \scanline[132][5] ;
 wire \scanline[132][6] ;
 wire \scanline[133][0] ;
 wire \scanline[133][1] ;
 wire \scanline[133][2] ;
 wire \scanline[133][3] ;
 wire \scanline[133][4] ;
 wire \scanline[133][5] ;
 wire \scanline[133][6] ;
 wire \scanline[134][0] ;
 wire \scanline[134][1] ;
 wire \scanline[134][2] ;
 wire \scanline[134][3] ;
 wire \scanline[134][4] ;
 wire \scanline[134][5] ;
 wire \scanline[134][6] ;
 wire \scanline[135][0] ;
 wire \scanline[135][1] ;
 wire \scanline[135][2] ;
 wire \scanline[135][3] ;
 wire \scanline[135][4] ;
 wire \scanline[135][5] ;
 wire \scanline[135][6] ;
 wire \scanline[136][0] ;
 wire \scanline[136][1] ;
 wire \scanline[136][2] ;
 wire \scanline[136][3] ;
 wire \scanline[136][4] ;
 wire \scanline[136][5] ;
 wire \scanline[136][6] ;
 wire \scanline[137][0] ;
 wire \scanline[137][1] ;
 wire \scanline[137][2] ;
 wire \scanline[137][3] ;
 wire \scanline[137][4] ;
 wire \scanline[137][5] ;
 wire \scanline[137][6] ;
 wire \scanline[138][0] ;
 wire \scanline[138][1] ;
 wire \scanline[138][2] ;
 wire \scanline[138][3] ;
 wire \scanline[138][4] ;
 wire \scanline[138][5] ;
 wire \scanline[138][6] ;
 wire \scanline[139][0] ;
 wire \scanline[139][1] ;
 wire \scanline[139][2] ;
 wire \scanline[139][3] ;
 wire \scanline[139][4] ;
 wire \scanline[139][5] ;
 wire \scanline[139][6] ;
 wire \scanline[13][0] ;
 wire \scanline[13][1] ;
 wire \scanline[13][2] ;
 wire \scanline[13][3] ;
 wire \scanline[13][4] ;
 wire \scanline[13][5] ;
 wire \scanline[13][6] ;
 wire \scanline[140][0] ;
 wire \scanline[140][1] ;
 wire \scanline[140][2] ;
 wire \scanline[140][3] ;
 wire \scanline[140][4] ;
 wire \scanline[140][5] ;
 wire \scanline[140][6] ;
 wire \scanline[141][0] ;
 wire \scanline[141][1] ;
 wire \scanline[141][2] ;
 wire \scanline[141][3] ;
 wire \scanline[141][4] ;
 wire \scanline[141][5] ;
 wire \scanline[141][6] ;
 wire \scanline[142][0] ;
 wire \scanline[142][1] ;
 wire \scanline[142][2] ;
 wire \scanline[142][3] ;
 wire \scanline[142][4] ;
 wire \scanline[142][5] ;
 wire \scanline[142][6] ;
 wire \scanline[143][0] ;
 wire \scanline[143][1] ;
 wire \scanline[143][2] ;
 wire \scanline[143][3] ;
 wire \scanline[143][4] ;
 wire \scanline[143][5] ;
 wire \scanline[143][6] ;
 wire \scanline[144][0] ;
 wire \scanline[144][1] ;
 wire \scanline[144][2] ;
 wire \scanline[144][3] ;
 wire \scanline[144][4] ;
 wire \scanline[144][5] ;
 wire \scanline[144][6] ;
 wire \scanline[145][0] ;
 wire \scanline[145][1] ;
 wire \scanline[145][2] ;
 wire \scanline[145][3] ;
 wire \scanline[145][4] ;
 wire \scanline[145][5] ;
 wire \scanline[145][6] ;
 wire \scanline[146][0] ;
 wire \scanline[146][1] ;
 wire \scanline[146][2] ;
 wire \scanline[146][3] ;
 wire \scanline[146][4] ;
 wire \scanline[146][5] ;
 wire \scanline[146][6] ;
 wire \scanline[147][0] ;
 wire \scanline[147][1] ;
 wire \scanline[147][2] ;
 wire \scanline[147][3] ;
 wire \scanline[147][4] ;
 wire \scanline[147][5] ;
 wire \scanline[147][6] ;
 wire \scanline[148][0] ;
 wire \scanline[148][1] ;
 wire \scanline[148][2] ;
 wire \scanline[148][3] ;
 wire \scanline[148][4] ;
 wire \scanline[148][5] ;
 wire \scanline[148][6] ;
 wire \scanline[149][0] ;
 wire \scanline[149][1] ;
 wire \scanline[149][2] ;
 wire \scanline[149][3] ;
 wire \scanline[149][4] ;
 wire \scanline[149][5] ;
 wire \scanline[149][6] ;
 wire \scanline[14][0] ;
 wire \scanline[14][1] ;
 wire \scanline[14][2] ;
 wire \scanline[14][3] ;
 wire \scanline[14][4] ;
 wire \scanline[14][5] ;
 wire \scanline[14][6] ;
 wire \scanline[150][0] ;
 wire \scanline[150][1] ;
 wire \scanline[150][2] ;
 wire \scanline[150][3] ;
 wire \scanline[150][4] ;
 wire \scanline[150][5] ;
 wire \scanline[150][6] ;
 wire \scanline[151][0] ;
 wire \scanline[151][1] ;
 wire \scanline[151][2] ;
 wire \scanline[151][3] ;
 wire \scanline[151][4] ;
 wire \scanline[151][5] ;
 wire \scanline[151][6] ;
 wire \scanline[152][0] ;
 wire \scanline[152][1] ;
 wire \scanline[152][2] ;
 wire \scanline[152][3] ;
 wire \scanline[152][4] ;
 wire \scanline[152][5] ;
 wire \scanline[152][6] ;
 wire \scanline[153][0] ;
 wire \scanline[153][1] ;
 wire \scanline[153][2] ;
 wire \scanline[153][3] ;
 wire \scanline[153][4] ;
 wire \scanline[153][5] ;
 wire \scanline[153][6] ;
 wire \scanline[154][0] ;
 wire \scanline[154][1] ;
 wire \scanline[154][2] ;
 wire \scanline[154][3] ;
 wire \scanline[154][4] ;
 wire \scanline[154][5] ;
 wire \scanline[154][6] ;
 wire \scanline[155][0] ;
 wire \scanline[155][1] ;
 wire \scanline[155][2] ;
 wire \scanline[155][3] ;
 wire \scanline[155][4] ;
 wire \scanline[155][5] ;
 wire \scanline[155][6] ;
 wire \scanline[156][0] ;
 wire \scanline[156][1] ;
 wire \scanline[156][2] ;
 wire \scanline[156][3] ;
 wire \scanline[156][4] ;
 wire \scanline[156][5] ;
 wire \scanline[156][6] ;
 wire \scanline[157][0] ;
 wire \scanline[157][1] ;
 wire \scanline[157][2] ;
 wire \scanline[157][3] ;
 wire \scanline[157][4] ;
 wire \scanline[157][5] ;
 wire \scanline[157][6] ;
 wire \scanline[158][0] ;
 wire \scanline[158][1] ;
 wire \scanline[158][2] ;
 wire \scanline[158][3] ;
 wire \scanline[158][4] ;
 wire \scanline[158][5] ;
 wire \scanline[158][6] ;
 wire \scanline[159][0] ;
 wire \scanline[159][1] ;
 wire \scanline[159][2] ;
 wire \scanline[159][3] ;
 wire \scanline[159][4] ;
 wire \scanline[159][5] ;
 wire \scanline[159][6] ;
 wire \scanline[15][0] ;
 wire \scanline[15][1] ;
 wire \scanline[15][2] ;
 wire \scanline[15][3] ;
 wire \scanline[15][4] ;
 wire \scanline[15][5] ;
 wire \scanline[15][6] ;
 wire \scanline[16][0] ;
 wire \scanline[16][1] ;
 wire \scanline[16][2] ;
 wire \scanline[16][3] ;
 wire \scanline[16][4] ;
 wire \scanline[16][5] ;
 wire \scanline[16][6] ;
 wire \scanline[17][0] ;
 wire \scanline[17][1] ;
 wire \scanline[17][2] ;
 wire \scanline[17][3] ;
 wire \scanline[17][4] ;
 wire \scanline[17][5] ;
 wire \scanline[17][6] ;
 wire \scanline[18][0] ;
 wire \scanline[18][1] ;
 wire \scanline[18][2] ;
 wire \scanline[18][3] ;
 wire \scanline[18][4] ;
 wire \scanline[18][5] ;
 wire \scanline[18][6] ;
 wire \scanline[19][0] ;
 wire \scanline[19][1] ;
 wire \scanline[19][2] ;
 wire \scanline[19][3] ;
 wire \scanline[19][4] ;
 wire \scanline[19][5] ;
 wire \scanline[19][6] ;
 wire \scanline[1][0] ;
 wire \scanline[1][1] ;
 wire \scanline[1][2] ;
 wire \scanline[1][3] ;
 wire \scanline[1][4] ;
 wire \scanline[1][5] ;
 wire \scanline[1][6] ;
 wire \scanline[20][0] ;
 wire \scanline[20][1] ;
 wire \scanline[20][2] ;
 wire \scanline[20][3] ;
 wire \scanline[20][4] ;
 wire \scanline[20][5] ;
 wire \scanline[20][6] ;
 wire \scanline[21][0] ;
 wire \scanline[21][1] ;
 wire \scanline[21][2] ;
 wire \scanline[21][3] ;
 wire \scanline[21][4] ;
 wire \scanline[21][5] ;
 wire \scanline[21][6] ;
 wire \scanline[22][0] ;
 wire \scanline[22][1] ;
 wire \scanline[22][2] ;
 wire \scanline[22][3] ;
 wire \scanline[22][4] ;
 wire \scanline[22][5] ;
 wire \scanline[22][6] ;
 wire \scanline[23][0] ;
 wire \scanline[23][1] ;
 wire \scanline[23][2] ;
 wire \scanline[23][3] ;
 wire \scanline[23][4] ;
 wire \scanline[23][5] ;
 wire \scanline[23][6] ;
 wire \scanline[24][0] ;
 wire \scanline[24][1] ;
 wire \scanline[24][2] ;
 wire \scanline[24][3] ;
 wire \scanline[24][4] ;
 wire \scanline[24][5] ;
 wire \scanline[24][6] ;
 wire \scanline[25][0] ;
 wire \scanline[25][1] ;
 wire \scanline[25][2] ;
 wire \scanline[25][3] ;
 wire \scanline[25][4] ;
 wire \scanline[25][5] ;
 wire \scanline[25][6] ;
 wire \scanline[26][0] ;
 wire \scanline[26][1] ;
 wire \scanline[26][2] ;
 wire \scanline[26][3] ;
 wire \scanline[26][4] ;
 wire \scanline[26][5] ;
 wire \scanline[26][6] ;
 wire \scanline[27][0] ;
 wire \scanline[27][1] ;
 wire \scanline[27][2] ;
 wire \scanline[27][3] ;
 wire \scanline[27][4] ;
 wire \scanline[27][5] ;
 wire \scanline[27][6] ;
 wire \scanline[28][0] ;
 wire \scanline[28][1] ;
 wire \scanline[28][2] ;
 wire \scanline[28][3] ;
 wire \scanline[28][4] ;
 wire \scanline[28][5] ;
 wire \scanline[28][6] ;
 wire \scanline[29][0] ;
 wire \scanline[29][1] ;
 wire \scanline[29][2] ;
 wire \scanline[29][3] ;
 wire \scanline[29][4] ;
 wire \scanline[29][5] ;
 wire \scanline[29][6] ;
 wire \scanline[2][0] ;
 wire \scanline[2][1] ;
 wire \scanline[2][2] ;
 wire \scanline[2][3] ;
 wire \scanline[2][4] ;
 wire \scanline[2][5] ;
 wire \scanline[2][6] ;
 wire \scanline[30][0] ;
 wire \scanline[30][1] ;
 wire \scanline[30][2] ;
 wire \scanline[30][3] ;
 wire \scanline[30][4] ;
 wire \scanline[30][5] ;
 wire \scanline[30][6] ;
 wire \scanline[31][0] ;
 wire \scanline[31][1] ;
 wire \scanline[31][2] ;
 wire \scanline[31][3] ;
 wire \scanline[31][4] ;
 wire \scanline[31][5] ;
 wire \scanline[31][6] ;
 wire \scanline[32][0] ;
 wire \scanline[32][1] ;
 wire \scanline[32][2] ;
 wire \scanline[32][3] ;
 wire \scanline[32][4] ;
 wire \scanline[32][5] ;
 wire \scanline[32][6] ;
 wire \scanline[33][0] ;
 wire \scanline[33][1] ;
 wire \scanline[33][2] ;
 wire \scanline[33][3] ;
 wire \scanline[33][4] ;
 wire \scanline[33][5] ;
 wire \scanline[33][6] ;
 wire \scanline[34][0] ;
 wire \scanline[34][1] ;
 wire \scanline[34][2] ;
 wire \scanline[34][3] ;
 wire \scanline[34][4] ;
 wire \scanline[34][5] ;
 wire \scanline[34][6] ;
 wire \scanline[35][0] ;
 wire \scanline[35][1] ;
 wire \scanline[35][2] ;
 wire \scanline[35][3] ;
 wire \scanline[35][4] ;
 wire \scanline[35][5] ;
 wire \scanline[35][6] ;
 wire \scanline[36][0] ;
 wire \scanline[36][1] ;
 wire \scanline[36][2] ;
 wire \scanline[36][3] ;
 wire \scanline[36][4] ;
 wire \scanline[36][5] ;
 wire \scanline[36][6] ;
 wire \scanline[37][0] ;
 wire \scanline[37][1] ;
 wire \scanline[37][2] ;
 wire \scanline[37][3] ;
 wire \scanline[37][4] ;
 wire \scanline[37][5] ;
 wire \scanline[37][6] ;
 wire \scanline[38][0] ;
 wire \scanline[38][1] ;
 wire \scanline[38][2] ;
 wire \scanline[38][3] ;
 wire \scanline[38][4] ;
 wire \scanline[38][5] ;
 wire \scanline[38][6] ;
 wire \scanline[39][0] ;
 wire \scanline[39][1] ;
 wire \scanline[39][2] ;
 wire \scanline[39][3] ;
 wire \scanline[39][4] ;
 wire \scanline[39][5] ;
 wire \scanline[39][6] ;
 wire \scanline[3][0] ;
 wire \scanline[3][1] ;
 wire \scanline[3][2] ;
 wire \scanline[3][3] ;
 wire \scanline[3][4] ;
 wire \scanline[3][5] ;
 wire \scanline[3][6] ;
 wire \scanline[40][0] ;
 wire \scanline[40][1] ;
 wire \scanline[40][2] ;
 wire \scanline[40][3] ;
 wire \scanline[40][4] ;
 wire \scanline[40][5] ;
 wire \scanline[40][6] ;
 wire \scanline[41][0] ;
 wire \scanline[41][1] ;
 wire \scanline[41][2] ;
 wire \scanline[41][3] ;
 wire \scanline[41][4] ;
 wire \scanline[41][5] ;
 wire \scanline[41][6] ;
 wire \scanline[42][0] ;
 wire \scanline[42][1] ;
 wire \scanline[42][2] ;
 wire \scanline[42][3] ;
 wire \scanline[42][4] ;
 wire \scanline[42][5] ;
 wire \scanline[42][6] ;
 wire \scanline[43][0] ;
 wire \scanline[43][1] ;
 wire \scanline[43][2] ;
 wire \scanline[43][3] ;
 wire \scanline[43][4] ;
 wire \scanline[43][5] ;
 wire \scanline[43][6] ;
 wire \scanline[44][0] ;
 wire \scanline[44][1] ;
 wire \scanline[44][2] ;
 wire \scanline[44][3] ;
 wire \scanline[44][4] ;
 wire \scanline[44][5] ;
 wire \scanline[44][6] ;
 wire \scanline[45][0] ;
 wire \scanline[45][1] ;
 wire \scanline[45][2] ;
 wire \scanline[45][3] ;
 wire \scanline[45][4] ;
 wire \scanline[45][5] ;
 wire \scanline[45][6] ;
 wire \scanline[46][0] ;
 wire \scanline[46][1] ;
 wire \scanline[46][2] ;
 wire \scanline[46][3] ;
 wire \scanline[46][4] ;
 wire \scanline[46][5] ;
 wire \scanline[46][6] ;
 wire \scanline[47][0] ;
 wire \scanline[47][1] ;
 wire \scanline[47][2] ;
 wire \scanline[47][3] ;
 wire \scanline[47][4] ;
 wire \scanline[47][5] ;
 wire \scanline[47][6] ;
 wire \scanline[48][0] ;
 wire \scanline[48][1] ;
 wire \scanline[48][2] ;
 wire \scanline[48][3] ;
 wire \scanline[48][4] ;
 wire \scanline[48][5] ;
 wire \scanline[48][6] ;
 wire \scanline[49][0] ;
 wire \scanline[49][1] ;
 wire \scanline[49][2] ;
 wire \scanline[49][3] ;
 wire \scanline[49][4] ;
 wire \scanline[49][5] ;
 wire \scanline[49][6] ;
 wire \scanline[4][0] ;
 wire \scanline[4][1] ;
 wire \scanline[4][2] ;
 wire \scanline[4][3] ;
 wire \scanline[4][4] ;
 wire \scanline[4][5] ;
 wire \scanline[4][6] ;
 wire \scanline[50][0] ;
 wire \scanline[50][1] ;
 wire \scanline[50][2] ;
 wire \scanline[50][3] ;
 wire \scanline[50][4] ;
 wire \scanline[50][5] ;
 wire \scanline[50][6] ;
 wire \scanline[51][0] ;
 wire \scanline[51][1] ;
 wire \scanline[51][2] ;
 wire \scanline[51][3] ;
 wire \scanline[51][4] ;
 wire \scanline[51][5] ;
 wire \scanline[51][6] ;
 wire \scanline[52][0] ;
 wire \scanline[52][1] ;
 wire \scanline[52][2] ;
 wire \scanline[52][3] ;
 wire \scanline[52][4] ;
 wire \scanline[52][5] ;
 wire \scanline[52][6] ;
 wire \scanline[53][0] ;
 wire \scanline[53][1] ;
 wire \scanline[53][2] ;
 wire \scanline[53][3] ;
 wire \scanline[53][4] ;
 wire \scanline[53][5] ;
 wire \scanline[53][6] ;
 wire \scanline[54][0] ;
 wire \scanline[54][1] ;
 wire \scanline[54][2] ;
 wire \scanline[54][3] ;
 wire \scanline[54][4] ;
 wire \scanline[54][5] ;
 wire \scanline[54][6] ;
 wire \scanline[55][0] ;
 wire \scanline[55][1] ;
 wire \scanline[55][2] ;
 wire \scanline[55][3] ;
 wire \scanline[55][4] ;
 wire \scanline[55][5] ;
 wire \scanline[55][6] ;
 wire \scanline[56][0] ;
 wire \scanline[56][1] ;
 wire \scanline[56][2] ;
 wire \scanline[56][3] ;
 wire \scanline[56][4] ;
 wire \scanline[56][5] ;
 wire \scanline[56][6] ;
 wire \scanline[57][0] ;
 wire \scanline[57][1] ;
 wire \scanline[57][2] ;
 wire \scanline[57][3] ;
 wire \scanline[57][4] ;
 wire \scanline[57][5] ;
 wire \scanline[57][6] ;
 wire \scanline[58][0] ;
 wire \scanline[58][1] ;
 wire \scanline[58][2] ;
 wire \scanline[58][3] ;
 wire \scanline[58][4] ;
 wire \scanline[58][5] ;
 wire \scanline[58][6] ;
 wire \scanline[59][0] ;
 wire \scanline[59][1] ;
 wire \scanline[59][2] ;
 wire \scanline[59][3] ;
 wire \scanline[59][4] ;
 wire \scanline[59][5] ;
 wire \scanline[59][6] ;
 wire \scanline[5][0] ;
 wire \scanline[5][1] ;
 wire \scanline[5][2] ;
 wire \scanline[5][3] ;
 wire \scanline[5][4] ;
 wire \scanline[5][5] ;
 wire \scanline[5][6] ;
 wire \scanline[60][0] ;
 wire \scanline[60][1] ;
 wire \scanline[60][2] ;
 wire \scanline[60][3] ;
 wire \scanline[60][4] ;
 wire \scanline[60][5] ;
 wire \scanline[60][6] ;
 wire \scanline[61][0] ;
 wire \scanline[61][1] ;
 wire \scanline[61][2] ;
 wire \scanline[61][3] ;
 wire \scanline[61][4] ;
 wire \scanline[61][5] ;
 wire \scanline[61][6] ;
 wire \scanline[62][0] ;
 wire \scanline[62][1] ;
 wire \scanline[62][2] ;
 wire \scanline[62][3] ;
 wire \scanline[62][4] ;
 wire \scanline[62][5] ;
 wire \scanline[62][6] ;
 wire \scanline[63][0] ;
 wire \scanline[63][1] ;
 wire \scanline[63][2] ;
 wire \scanline[63][3] ;
 wire \scanline[63][4] ;
 wire \scanline[63][5] ;
 wire \scanline[63][6] ;
 wire \scanline[64][0] ;
 wire \scanline[64][1] ;
 wire \scanline[64][2] ;
 wire \scanline[64][3] ;
 wire \scanline[64][4] ;
 wire \scanline[64][5] ;
 wire \scanline[64][6] ;
 wire \scanline[65][0] ;
 wire \scanline[65][1] ;
 wire \scanline[65][2] ;
 wire \scanline[65][3] ;
 wire \scanline[65][4] ;
 wire \scanline[65][5] ;
 wire \scanline[65][6] ;
 wire \scanline[66][0] ;
 wire \scanline[66][1] ;
 wire \scanline[66][2] ;
 wire \scanline[66][3] ;
 wire \scanline[66][4] ;
 wire \scanline[66][5] ;
 wire \scanline[66][6] ;
 wire \scanline[67][0] ;
 wire \scanline[67][1] ;
 wire \scanline[67][2] ;
 wire \scanline[67][3] ;
 wire \scanline[67][4] ;
 wire \scanline[67][5] ;
 wire \scanline[67][6] ;
 wire \scanline[68][0] ;
 wire \scanline[68][1] ;
 wire \scanline[68][2] ;
 wire \scanline[68][3] ;
 wire \scanline[68][4] ;
 wire \scanline[68][5] ;
 wire \scanline[68][6] ;
 wire \scanline[69][0] ;
 wire \scanline[69][1] ;
 wire \scanline[69][2] ;
 wire \scanline[69][3] ;
 wire \scanline[69][4] ;
 wire \scanline[69][5] ;
 wire \scanline[69][6] ;
 wire \scanline[6][0] ;
 wire \scanline[6][1] ;
 wire \scanline[6][2] ;
 wire \scanline[6][3] ;
 wire \scanline[6][4] ;
 wire \scanline[6][5] ;
 wire \scanline[6][6] ;
 wire \scanline[70][0] ;
 wire \scanline[70][1] ;
 wire \scanline[70][2] ;
 wire \scanline[70][3] ;
 wire \scanline[70][4] ;
 wire \scanline[70][5] ;
 wire \scanline[70][6] ;
 wire \scanline[71][0] ;
 wire \scanline[71][1] ;
 wire \scanline[71][2] ;
 wire \scanline[71][3] ;
 wire \scanline[71][4] ;
 wire \scanline[71][5] ;
 wire \scanline[71][6] ;
 wire \scanline[72][0] ;
 wire \scanline[72][1] ;
 wire \scanline[72][2] ;
 wire \scanline[72][3] ;
 wire \scanline[72][4] ;
 wire \scanline[72][5] ;
 wire \scanline[72][6] ;
 wire \scanline[73][0] ;
 wire \scanline[73][1] ;
 wire \scanline[73][2] ;
 wire \scanline[73][3] ;
 wire \scanline[73][4] ;
 wire \scanline[73][5] ;
 wire \scanline[73][6] ;
 wire \scanline[74][0] ;
 wire \scanline[74][1] ;
 wire \scanline[74][2] ;
 wire \scanline[74][3] ;
 wire \scanline[74][4] ;
 wire \scanline[74][5] ;
 wire \scanline[74][6] ;
 wire \scanline[75][0] ;
 wire \scanline[75][1] ;
 wire \scanline[75][2] ;
 wire \scanline[75][3] ;
 wire \scanline[75][4] ;
 wire \scanline[75][5] ;
 wire \scanline[75][6] ;
 wire \scanline[76][0] ;
 wire \scanline[76][1] ;
 wire \scanline[76][2] ;
 wire \scanline[76][3] ;
 wire \scanline[76][4] ;
 wire \scanline[76][5] ;
 wire \scanline[76][6] ;
 wire \scanline[77][0] ;
 wire \scanline[77][1] ;
 wire \scanline[77][2] ;
 wire \scanline[77][3] ;
 wire \scanline[77][4] ;
 wire \scanline[77][5] ;
 wire \scanline[77][6] ;
 wire \scanline[78][0] ;
 wire \scanline[78][1] ;
 wire \scanline[78][2] ;
 wire \scanline[78][3] ;
 wire \scanline[78][4] ;
 wire \scanline[78][5] ;
 wire \scanline[78][6] ;
 wire \scanline[79][0] ;
 wire \scanline[79][1] ;
 wire \scanline[79][2] ;
 wire \scanline[79][3] ;
 wire \scanline[79][4] ;
 wire \scanline[79][5] ;
 wire \scanline[79][6] ;
 wire \scanline[7][0] ;
 wire \scanline[7][1] ;
 wire \scanline[7][2] ;
 wire \scanline[7][3] ;
 wire \scanline[7][4] ;
 wire \scanline[7][5] ;
 wire \scanline[7][6] ;
 wire \scanline[80][0] ;
 wire \scanline[80][1] ;
 wire \scanline[80][2] ;
 wire \scanline[80][3] ;
 wire \scanline[80][4] ;
 wire \scanline[80][5] ;
 wire \scanline[80][6] ;
 wire \scanline[81][0] ;
 wire \scanline[81][1] ;
 wire \scanline[81][2] ;
 wire \scanline[81][3] ;
 wire \scanline[81][4] ;
 wire \scanline[81][5] ;
 wire \scanline[81][6] ;
 wire \scanline[82][0] ;
 wire \scanline[82][1] ;
 wire \scanline[82][2] ;
 wire \scanline[82][3] ;
 wire \scanline[82][4] ;
 wire \scanline[82][5] ;
 wire \scanline[82][6] ;
 wire \scanline[83][0] ;
 wire \scanline[83][1] ;
 wire \scanline[83][2] ;
 wire \scanline[83][3] ;
 wire \scanline[83][4] ;
 wire \scanline[83][5] ;
 wire \scanline[83][6] ;
 wire \scanline[84][0] ;
 wire \scanline[84][1] ;
 wire \scanline[84][2] ;
 wire \scanline[84][3] ;
 wire \scanline[84][4] ;
 wire \scanline[84][5] ;
 wire \scanline[84][6] ;
 wire \scanline[85][0] ;
 wire \scanline[85][1] ;
 wire \scanline[85][2] ;
 wire \scanline[85][3] ;
 wire \scanline[85][4] ;
 wire \scanline[85][5] ;
 wire \scanline[85][6] ;
 wire \scanline[86][0] ;
 wire \scanline[86][1] ;
 wire \scanline[86][2] ;
 wire \scanline[86][3] ;
 wire \scanline[86][4] ;
 wire \scanline[86][5] ;
 wire \scanline[86][6] ;
 wire \scanline[87][0] ;
 wire \scanline[87][1] ;
 wire \scanline[87][2] ;
 wire \scanline[87][3] ;
 wire \scanline[87][4] ;
 wire \scanline[87][5] ;
 wire \scanline[87][6] ;
 wire \scanline[88][0] ;
 wire \scanline[88][1] ;
 wire \scanline[88][2] ;
 wire \scanline[88][3] ;
 wire \scanline[88][4] ;
 wire \scanline[88][5] ;
 wire \scanline[88][6] ;
 wire \scanline[89][0] ;
 wire \scanline[89][1] ;
 wire \scanline[89][2] ;
 wire \scanline[89][3] ;
 wire \scanline[89][4] ;
 wire \scanline[89][5] ;
 wire \scanline[89][6] ;
 wire \scanline[8][0] ;
 wire \scanline[8][1] ;
 wire \scanline[8][2] ;
 wire \scanline[8][3] ;
 wire \scanline[8][4] ;
 wire \scanline[8][5] ;
 wire \scanline[8][6] ;
 wire \scanline[90][0] ;
 wire \scanline[90][1] ;
 wire \scanline[90][2] ;
 wire \scanline[90][3] ;
 wire \scanline[90][4] ;
 wire \scanline[90][5] ;
 wire \scanline[90][6] ;
 wire \scanline[91][0] ;
 wire \scanline[91][1] ;
 wire \scanline[91][2] ;
 wire \scanline[91][3] ;
 wire \scanline[91][4] ;
 wire \scanline[91][5] ;
 wire \scanline[91][6] ;
 wire \scanline[92][0] ;
 wire \scanline[92][1] ;
 wire \scanline[92][2] ;
 wire \scanline[92][3] ;
 wire \scanline[92][4] ;
 wire \scanline[92][5] ;
 wire \scanline[92][6] ;
 wire \scanline[93][0] ;
 wire \scanline[93][1] ;
 wire \scanline[93][2] ;
 wire \scanline[93][3] ;
 wire \scanline[93][4] ;
 wire \scanline[93][5] ;
 wire \scanline[93][6] ;
 wire \scanline[94][0] ;
 wire \scanline[94][1] ;
 wire \scanline[94][2] ;
 wire \scanline[94][3] ;
 wire \scanline[94][4] ;
 wire \scanline[94][5] ;
 wire \scanline[94][6] ;
 wire \scanline[95][0] ;
 wire \scanline[95][1] ;
 wire \scanline[95][2] ;
 wire \scanline[95][3] ;
 wire \scanline[95][4] ;
 wire \scanline[95][5] ;
 wire \scanline[95][6] ;
 wire \scanline[96][0] ;
 wire \scanline[96][1] ;
 wire \scanline[96][2] ;
 wire \scanline[96][3] ;
 wire \scanline[96][4] ;
 wire \scanline[96][5] ;
 wire \scanline[96][6] ;
 wire \scanline[97][0] ;
 wire \scanline[97][1] ;
 wire \scanline[97][2] ;
 wire \scanline[97][3] ;
 wire \scanline[97][4] ;
 wire \scanline[97][5] ;
 wire \scanline[97][6] ;
 wire \scanline[98][0] ;
 wire \scanline[98][1] ;
 wire \scanline[98][2] ;
 wire \scanline[98][3] ;
 wire \scanline[98][4] ;
 wire \scanline[98][5] ;
 wire \scanline[98][6] ;
 wire \scanline[99][0] ;
 wire \scanline[99][1] ;
 wire \scanline[99][2] ;
 wire \scanline[99][3] ;
 wire \scanline[99][4] ;
 wire \scanline[99][5] ;
 wire \scanline[99][6] ;
 wire \scanline[9][0] ;
 wire \scanline[9][1] ;
 wire \scanline[9][2] ;
 wire \scanline[9][3] ;
 wire \scanline[9][4] ;
 wire \scanline[9][5] ;
 wire \scanline[9][6] ;
 wire spi_data_ready_last;
 wire spi_restart;
 wire tia_vsync_last;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire clknet_leaf_0_clk;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_338_clk;
 wire clknet_leaf_339_clk;
 wire clknet_leaf_340_clk;
 wire clknet_leaf_341_clk;
 wire clknet_leaf_342_clk;
 wire clknet_leaf_343_clk;
 wire clknet_leaf_344_clk;
 wire clknet_leaf_345_clk;
 wire clknet_leaf_346_clk;
 wire clknet_leaf_347_clk;
 wire clknet_leaf_348_clk;
 wire clknet_leaf_349_clk;
 wire clknet_leaf_350_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_353_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_356_clk;
 wire clknet_leaf_357_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_359_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_361_clk;
 wire clknet_leaf_362_clk;
 wire clknet_leaf_363_clk;
 wire clknet_leaf_364_clk;
 wire clknet_leaf_365_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net7570;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7574;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net7578;
 wire net7579;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7584;
 wire net7585;
 wire net7586;
 wire net7587;
 wire net7588;
 wire net7589;
 wire net7590;
 wire net7591;
 wire net7592;
 wire net7593;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7597;
 wire net7598;
 wire net7599;
 wire net7600;
 wire net7601;

 sg13g2_inv_1 _16791_ (.Y(_08473_),
    .A(\flash_rom.fsm_state[0] ));
 sg13g2_inv_1 _16792_ (.Y(_08474_),
    .A(\flash_rom.nibbles_remaining[0] ));
 sg13g2_inv_1 _16793_ (.Y(_08475_),
    .A(net4534));
 sg13g2_inv_1 _16794_ (.Y(_08476_),
    .A(net6809));
 sg13g2_inv_1 _16795_ (.Y(_08477_),
    .A(net7227));
 sg13g2_inv_1 _16796_ (.Y(_08478_),
    .A(net7083));
 sg13g2_inv_1 _16797_ (.Y(_08479_),
    .A(net7147));
 sg13g2_inv_1 _16798_ (.Y(_08480_),
    .A(net6716));
 sg13g2_inv_1 _16799_ (.Y(_08481_),
    .A(net6678));
 sg13g2_inv_1 _16800_ (.Y(_08482_),
    .A(net6709));
 sg13g2_inv_1 _16801_ (.Y(_08483_),
    .A(net7231));
 sg13g2_inv_1 _16802_ (.Y(_08484_),
    .A(net7094));
 sg13g2_inv_1 _16803_ (.Y(_08485_),
    .A(net6924));
 sg13g2_inv_1 _16804_ (.Y(_08486_),
    .A(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_inv_1 _16805_ (.Y(_08487_),
    .A(net2935));
 sg13g2_inv_1 _16806_ (.Y(_08488_),
    .A(net2955));
 sg13g2_inv_1 _16807_ (.Y(_08489_),
    .A(\atari2600.clk_counter[0] ));
 sg13g2_inv_1 _16808_ (.Y(_08490_),
    .A(net2946));
 sg13g2_inv_1 _16809_ (.Y(_08491_),
    .A(\atari2600.tia.poly9_r.x[4] ));
 sg13g2_inv_1 _16810_ (.Y(_08492_),
    .A(\atari2600.tia.p9_r ));
 sg13g2_inv_1 _16811_ (.Y(_08493_),
    .A(net7201));
 sg13g2_inv_1 _16812_ (.Y(_08494_),
    .A(\atari2600.tia.p5_r ));
 sg13g2_inv_1 _16813_ (.Y(_08495_),
    .A(\atari2600.tia.poly4_r.x[1] ));
 sg13g2_inv_1 _16814_ (.Y(_08496_),
    .A(\atari2600.tia.poly9_l.x[4] ));
 sg13g2_inv_2 _16815_ (.Y(_08497_),
    .A(\atari2600.tia.p9_l ));
 sg13g2_inv_1 _16816_ (.Y(_08498_),
    .A(net6916));
 sg13g2_inv_1 _16817_ (.Y(_08499_),
    .A(\atari2600.tia.p5_l ));
 sg13g2_inv_1 _16818_ (.Y(_08500_),
    .A(\atari2600.tia.poly4_l.x[1] ));
 sg13g2_inv_1 _16819_ (.Y(_08501_),
    .A(\atari2600.tia.audf1[2] ));
 sg13g2_inv_2 _16820_ (.Y(_08502_),
    .A(\atari2600.tia.audf0[3] ));
 sg13g2_inv_1 _16821_ (.Y(_08503_),
    .A(\atari2600.tia.audf0[1] ));
 sg13g2_inv_1 _16822_ (.Y(_08504_),
    .A(\atari2600.tia.audf0[0] ));
 sg13g2_inv_1 _16823_ (.Y(_08505_),
    .A(\atari2600.tia.audc1[3] ));
 sg13g2_inv_1 _16824_ (.Y(_08506_),
    .A(\atari2600.tia.audc1[2] ));
 sg13g2_inv_1 _16825_ (.Y(_08507_),
    .A(\atari2600.tia.audc1[1] ));
 sg13g2_inv_1 _16826_ (.Y(_08508_),
    .A(\atari2600.tia.audc1[0] ));
 sg13g2_inv_1 _16827_ (.Y(_08509_),
    .A(\atari2600.tia.audc0[1] ));
 sg13g2_inv_1 _16828_ (.Y(_08510_),
    .A(\atari2600.tia.audc0[0] ));
 sg13g2_inv_1 _16829_ (.Y(_08511_),
    .A(\atari2600.tia.hmbl[3] ));
 sg13g2_inv_1 _16830_ (.Y(_08512_),
    .A(\atari2600.tia.hmbl[2] ));
 sg13g2_inv_1 _16831_ (.Y(_08513_),
    .A(\atari2600.tia.hmm0[3] ));
 sg13g2_inv_1 _16832_ (.Y(_08514_),
    .A(\atari2600.tia.hmm0[2] ));
 sg13g2_inv_1 _16833_ (.Y(_08515_),
    .A(net6266));
 sg13g2_inv_1 _16834_ (.Y(_08516_),
    .A(\atari2600.tia.hmp1[2] ));
 sg13g2_inv_1 _16835_ (.Y(_08517_),
    .A(net6267));
 sg13g2_inv_1 _16836_ (.Y(_08518_),
    .A(\atari2600.tia.hmp0[2] ));
 sg13g2_inv_1 _16837_ (.Y(_08519_),
    .A(\atari2600.tia.diag[38] ));
 sg13g2_inv_1 _16838_ (.Y(_08520_),
    .A(\atari2600.tia.diag[37] ));
 sg13g2_inv_1 _16839_ (.Y(_08521_),
    .A(\atari2600.tia.diag[36] ));
 sg13g2_inv_1 _16840_ (.Y(_08522_),
    .A(net7492));
 sg13g2_inv_1 _16841_ (.Y(_08523_),
    .A(net7494));
 sg13g2_inv_1 _16842_ (.Y(_08524_),
    .A(net7535));
 sg13g2_inv_2 _16843_ (.Y(_08525_),
    .A(net7459));
 sg13g2_inv_1 _16844_ (.Y(_08526_),
    .A(net7508));
 sg13g2_inv_1 _16845_ (.Y(_08527_),
    .A(net7545));
 sg13g2_inv_1 _16846_ (.Y(_08528_),
    .A(net7505));
 sg13g2_inv_1 _16847_ (.Y(_08529_),
    .A(net7507));
 sg13g2_inv_1 _16848_ (.Y(_08530_),
    .A(net7520));
 sg13g2_inv_2 _16849_ (.Y(_08531_),
    .A(\atari2600.tia.diag[62] ));
 sg13g2_inv_1 _16850_ (.Y(_08532_),
    .A(\atari2600.tia.diag[61] ));
 sg13g2_inv_1 _16851_ (.Y(_08533_),
    .A(net6270));
 sg13g2_inv_1 _16852_ (.Y(_08534_),
    .A(net6271));
 sg13g2_inv_1 _16853_ (.Y(_08535_),
    .A(\atari2600.tia.diag[58] ));
 sg13g2_inv_2 _16854_ (.Y(_08536_),
    .A(\atari2600.tia.diag[57] ));
 sg13g2_inv_2 _16855_ (.Y(_08537_),
    .A(\atari2600.tia.diag[70] ));
 sg13g2_inv_1 _16856_ (.Y(_08538_),
    .A(net6273));
 sg13g2_inv_1 _16857_ (.Y(_08539_),
    .A(net6275));
 sg13g2_inv_1 _16858_ (.Y(_08540_),
    .A(\atari2600.tia.diag[64] ));
 sg13g2_inv_2 _16859_ (.Y(_08541_),
    .A(\atari2600.tia.scorepf ));
 sg13g2_inv_1 _16860_ (.Y(_08542_),
    .A(\atari2600.tia.colupf[6] ));
 sg13g2_inv_1 _16861_ (.Y(_08543_),
    .A(\atari2600.tia.colupf[5] ));
 sg13g2_inv_1 _16862_ (.Y(_08544_),
    .A(\atari2600.tia.colupf[4] ));
 sg13g2_inv_1 _16863_ (.Y(_08545_),
    .A(net7341));
 sg13g2_inv_1 _16864_ (.Y(_08546_),
    .A(\atari2600.tia.colupf[2] ));
 sg13g2_inv_1 _16865_ (.Y(_08547_),
    .A(net7600));
 sg13g2_inv_1 _16866_ (.Y(_08548_),
    .A(\atari2600.tia.colup1[5] ));
 sg13g2_inv_1 _16867_ (.Y(_08549_),
    .A(\atari2600.tia.colup1[4] ));
 sg13g2_inv_1 _16868_ (.Y(_08550_),
    .A(\atari2600.tia.colup1[3] ));
 sg13g2_inv_1 _16869_ (.Y(_08551_),
    .A(\atari2600.tia.colubk[6] ));
 sg13g2_inv_1 _16870_ (.Y(_08552_),
    .A(\atari2600.tia.colubk[5] ));
 sg13g2_inv_1 _16871_ (.Y(_08553_),
    .A(\atari2600.tia.colubk[4] ));
 sg13g2_inv_1 _16872_ (.Y(_08554_),
    .A(\atari2600.tia.colubk[3] ));
 sg13g2_inv_1 _16873_ (.Y(_08555_),
    .A(\atari2600.tia.colubk[2] ));
 sg13g2_inv_1 _16874_ (.Y(_08556_),
    .A(\atari2600.tia.colubk[1] ));
 sg13g2_inv_1 _16875_ (.Y(_08557_),
    .A(net7461));
 sg13g2_inv_1 _16876_ (.Y(_08558_),
    .A(\flash_rom.addr[20] ));
 sg13g2_inv_1 _16877_ (.Y(_08559_),
    .A(\atari2600.tia.p0_w[4] ));
 sg13g2_inv_1 _16878_ (.Y(_08560_),
    .A(\atari2600.tia.p0_scale[1] ));
 sg13g2_inv_1 _16879_ (.Y(_08561_),
    .A(\atari2600.tia.p0_scale[0] ));
 sg13g2_inv_1 _16880_ (.Y(_08562_),
    .A(\atari2600.tia.p1_w[4] ));
 sg13g2_inv_1 _16881_ (.Y(_08563_),
    .A(net4324));
 sg13g2_inv_1 _16882_ (.Y(_08564_),
    .A(net7024));
 sg13g2_inv_1 _16883_ (.Y(_08565_),
    .A(net6597));
 sg13g2_inv_1 _16884_ (.Y(_08566_),
    .A(net7487));
 sg13g2_inv_1 _16885_ (.Y(_08567_),
    .A(net7159));
 sg13g2_inv_1 _16886_ (.Y(_08568_),
    .A(net4758));
 sg13g2_inv_1 _16887_ (.Y(_08569_),
    .A(net2933));
 sg13g2_inv_1 _16888_ (.Y(_08570_),
    .A(\atari2600.tia.vid_ypos[5] ));
 sg13g2_inv_1 _16889_ (.Y(_08571_),
    .A(\atari2600.tia.vid_ypos[4] ));
 sg13g2_inv_1 _16890_ (.Y(_08572_),
    .A(net7131));
 sg13g2_inv_1 _16891_ (.Y(_08573_),
    .A(\hvsync_gen.vga.vpos[4] ));
 sg13g2_inv_1 _16892_ (.Y(_08574_),
    .A(net3469));
 sg13g2_inv_1 _16893_ (.Y(_08575_),
    .A(_00071_));
 sg13g2_inv_1 _16894_ (.Y(_08576_),
    .A(net3154));
 sg13g2_inv_1 _16895_ (.Y(_08577_),
    .A(net7386));
 sg13g2_inv_1 _16896_ (.Y(_08578_),
    .A(net7119));
 sg13g2_inv_1 _16897_ (.Y(_08579_),
    .A(net7261));
 sg13g2_inv_1 _16898_ (.Y(_08580_),
    .A(net6251));
 sg13g2_inv_1 _16899_ (.Y(_08581_),
    .A(net4480));
 sg13g2_inv_1 _16900_ (.Y(_08582_),
    .A(\atari2600.cpu.C ));
 sg13g2_inv_1 _16901_ (.Y(_08583_),
    .A(_00077_));
 sg13g2_inv_1 _16902_ (.Y(_08584_),
    .A(net6864));
 sg13g2_inv_1 _16903_ (.Y(_08585_),
    .A(_00078_));
 sg13g2_inv_2 _16904_ (.Y(_08586_),
    .A(net7420));
 sg13g2_inv_2 _16905_ (.Y(_08587_),
    .A(net7238));
 sg13g2_inv_1 _16906_ (.Y(_08588_),
    .A(net7438));
 sg13g2_inv_1 _16907_ (.Y(_08589_),
    .A(net7455));
 sg13g2_inv_1 _16908_ (.Y(_08590_),
    .A(net7477));
 sg13g2_inv_1 _16909_ (.Y(_08591_),
    .A(\atari2600.cpu.rotate ));
 sg13g2_inv_1 _16910_ (.Y(_08592_),
    .A(net6247));
 sg13g2_inv_1 _16911_ (.Y(_08593_),
    .A(net7145));
 sg13g2_inv_1 _16912_ (.Y(_08594_),
    .A(net6248));
 sg13g2_inv_1 _16913_ (.Y(_08595_),
    .A(net7241));
 sg13g2_inv_2 _16914_ (.Y(_08596_),
    .A(_00086_));
 sg13g2_inv_1 _16915_ (.Y(_08597_),
    .A(_00090_));
 sg13g2_inv_1 _16916_ (.Y(_08598_),
    .A(net7175));
 sg13g2_inv_2 _16917_ (.Y(_08599_),
    .A(_00091_));
 sg13g2_inv_1 _16918_ (.Y(_08600_),
    .A(net7233));
 sg13g2_inv_1 _16919_ (.Y(_08601_),
    .A(net7246));
 sg13g2_inv_1 _16920_ (.Y(_08602_),
    .A(net7113));
 sg13g2_inv_1 _16921_ (.Y(_08603_),
    .A(\atari2600.address_bus_r[9] ));
 sg13g2_inv_1 _16922_ (.Y(_08604_),
    .A(net7329));
 sg13g2_inv_1 _16923_ (.Y(_08605_),
    .A(net7116));
 sg13g2_inv_1 _16924_ (.Y(_08606_),
    .A(net6964));
 sg13g2_inv_1 _16925_ (.Y(_08607_),
    .A(net7165));
 sg13g2_inv_1 _16926_ (.Y(_08608_),
    .A(_00093_));
 sg13g2_inv_1 _16927_ (.Y(_08609_),
    .A(net7369));
 sg13g2_inv_1 _16928_ (.Y(_08610_),
    .A(net7365));
 sg13g2_inv_1 _16929_ (.Y(_08611_),
    .A(net7281));
 sg13g2_inv_1 _16930_ (.Y(_08612_),
    .A(net7336));
 sg13g2_inv_1 _16931_ (.Y(_08613_),
    .A(net7422));
 sg13g2_inv_1 _16932_ (.Y(_08614_),
    .A(net7316));
 sg13g2_inv_1 _16933_ (.Y(_08615_),
    .A(net7323));
 sg13g2_inv_1 _16934_ (.Y(_08616_),
    .A(net7406));
 sg13g2_inv_2 _16935_ (.Y(_08617_),
    .A(net6549));
 sg13g2_inv_1 _16936_ (.Y(_08618_),
    .A(_00096_));
 sg13g2_inv_1 _16937_ (.Y(_08619_),
    .A(_00111_));
 sg13g2_inv_1 _16938_ (.Y(_08620_),
    .A(_00115_));
 sg13g2_inv_1 _16939_ (.Y(_08621_),
    .A(_00116_));
 sg13g2_inv_1 _16940_ (.Y(_08622_),
    .A(_00118_));
 sg13g2_inv_1 _16941_ (.Y(_08623_),
    .A(_00120_));
 sg13g2_inv_1 _16942_ (.Y(_08624_),
    .A(_00125_));
 sg13g2_inv_1 _16943_ (.Y(_08625_),
    .A(\flash_rom.data_ready ));
 sg13g2_inv_4 _16944_ (.A(net6501),
    .Y(_08626_));
 sg13g2_inv_1 _16945_ (.Y(_08627_),
    .A(net6502));
 sg13g2_inv_2 _16946_ (.Y(_08628_),
    .A(net6504));
 sg13g2_inv_4 _16947_ (.A(net6506),
    .Y(_08629_));
 sg13g2_inv_2 _16948_ (.Y(_08630_),
    .A(net6495));
 sg13g2_inv_1 _16949_ (.Y(_08631_),
    .A(net6490));
 sg13g2_inv_1 _16950_ (.Y(_08632_),
    .A(net6488));
 sg13g2_inv_4 _16951_ (.A(net6482),
    .Y(_08633_));
 sg13g2_inv_1 _16952_ (.Y(_08634_),
    .A(net3065));
 sg13g2_inv_1 _16953_ (.Y(_08635_),
    .A(net4321));
 sg13g2_inv_1 _16954_ (.Y(_08636_),
    .A(net6824));
 sg13g2_inv_1 _16955_ (.Y(_08637_),
    .A(net7170));
 sg13g2_inv_1 _16956_ (.Y(_08638_),
    .A(net7212));
 sg13g2_inv_2 _16957_ (.Y(_08639_),
    .A(net7523));
 sg13g2_inv_1 _16958_ (.Y(_08640_),
    .A(net3225));
 sg13g2_inv_1 _16959_ (.Y(_08641_),
    .A(net7204));
 sg13g2_inv_1 _16960_ (.Y(_08642_),
    .A(net4807));
 sg13g2_inv_1 _16961_ (.Y(_08643_),
    .A(net4421));
 sg13g2_inv_1 _16962_ (.Y(_08644_),
    .A(net3786));
 sg13g2_inv_1 _16963_ (.Y(_08645_),
    .A(net4450));
 sg13g2_inv_1 _16964_ (.Y(_08646_),
    .A(net4103));
 sg13g2_inv_1 _16965_ (.Y(_08647_),
    .A(net4350));
 sg13g2_inv_1 _16966_ (.Y(_08648_),
    .A(net4483));
 sg13g2_inv_1 _16967_ (.Y(_08649_),
    .A(net6845));
 sg13g2_inv_1 _16968_ (.Y(_08650_),
    .A(net4431));
 sg13g2_inv_1 _16969_ (.Y(_08651_),
    .A(net3422));
 sg13g2_inv_4 _16970_ (.A(net6160),
    .Y(_08652_));
 sg13g2_inv_2 _16971_ (.Y(_08653_),
    .A(net6128));
 sg13g2_inv_2 _16972_ (.Y(_08654_),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_inv_4 _16973_ (.A(net6125),
    .Y(_08655_));
 sg13g2_inv_4 _16974_ (.A(net6127),
    .Y(_08656_));
 sg13g2_inv_1 _16975_ (.Y(_08657_),
    .A(net7));
 sg13g2_inv_1 _16976_ (.Y(_08658_),
    .A(\atari2600.cpu.PC[13] ));
 sg13g2_inv_1 _16977_ (.Y(_08659_),
    .A(net7413));
 sg13g2_inv_1 _16978_ (.Y(_08660_),
    .A(_00138_));
 sg13g2_inv_2 _16979_ (.Y(_08661_),
    .A(_00142_));
 sg13g2_inv_1 _16980_ (.Y(_08662_),
    .A(_00150_));
 sg13g2_inv_1 _16981_ (.Y(_08663_),
    .A(net4492));
 sg13g2_inv_1 _16982_ (.Y(_08664_),
    .A(net4643));
 sg13g2_inv_1 _16983_ (.Y(_08665_),
    .A(net7128));
 sg13g2_inv_1 _16984_ (.Y(_08666_),
    .A(net7167));
 sg13g2_inv_1 _16985_ (.Y(_08667_),
    .A(net7157));
 sg13g2_inv_1 _16986_ (.Y(_08668_),
    .A(net4459));
 sg13g2_inv_1 _16987_ (.Y(_08669_),
    .A(net4779));
 sg13g2_inv_1 _16988_ (.Y(_08670_),
    .A(_00056_));
 sg13g2_inv_1 _16989_ (.Y(_08671_),
    .A(\scanline[157][1] ));
 sg13g2_inv_1 _16990_ (.Y(_08672_),
    .A(_00065_));
 sg13g2_inv_1 _16991_ (.Y(_08673_),
    .A(_00066_));
 sg13g2_inv_1 _16992_ (.Y(_08674_),
    .A(net7556));
 sg13g2_nor2_1 _16993_ (.A(\atari2600.clk_counter[7] ),
    .B(\atari2600.clk_counter[6] ),
    .Y(_08675_));
 sg13g2_nor4_1 _16994_ (.A(\atari2600.clk_counter[5] ),
    .B(\atari2600.clk_counter[4] ),
    .C(\atari2600.clk_counter[3] ),
    .D(\atari2600.clk_counter[2] ),
    .Y(_08676_));
 sg13g2_nand2_1 _16995_ (.Y(_08677_),
    .A(_08675_),
    .B(_08676_));
 sg13g2_nor2_1 _16996_ (.A(\atari2600.clk_counter[8] ),
    .B(_08677_),
    .Y(_08678_));
 sg13g2_or2_2 _16997_ (.X(_08679_),
    .B(_08677_),
    .A(\atari2600.clk_counter[8] ));
 sg13g2_nor3_2 _16998_ (.A(\atari2600.clk_counter[1] ),
    .B(_08489_),
    .C(_08679_),
    .Y(_08680_));
 sg13g2_nand2_1 _16999_ (.Y(_08681_),
    .A(_08570_),
    .B(\hvsync_gen.vga.vpos[6] ));
 sg13g2_nand2b_1 _17000_ (.Y(_08682_),
    .B(\atari2600.tia.vid_ypos[4] ),
    .A_N(\hvsync_gen.vga.vpos[5] ));
 sg13g2_nand2b_1 _17001_ (.Y(_08683_),
    .B(\hvsync_gen.vga.vpos[3] ),
    .A_N(\atari2600.tia.vid_ypos[2] ));
 sg13g2_nor2b_1 _17002_ (.A(\atari2600.tia.vid_ypos[1] ),
    .B_N(\hvsync_gen.vga.vpos[2] ),
    .Y(_08684_));
 sg13g2_nand2b_1 _17003_ (.Y(_08685_),
    .B(\atari2600.tia.vid_ypos[0] ),
    .A_N(\hvsync_gen.vga.vpos[1] ));
 sg13g2_nand2b_1 _17004_ (.Y(_08686_),
    .B(\atari2600.tia.vid_ypos[1] ),
    .A_N(\hvsync_gen.vga.vpos[2] ));
 sg13g2_o21ai_1 _17005_ (.B1(_08686_),
    .Y(_08687_),
    .A1(_08684_),
    .A2(_08685_));
 sg13g2_nor2b_1 _17006_ (.A(\hvsync_gen.vga.vpos[3] ),
    .B_N(\atari2600.tia.vid_ypos[2] ),
    .Y(_08688_));
 sg13g2_a221oi_1 _17007_ (.B2(_08687_),
    .C1(_08688_),
    .B1(_08683_),
    .A1(\atari2600.tia.vid_ypos[3] ),
    .Y(_08689_),
    .A2(_08573_));
 sg13g2_nand2_1 _17008_ (.Y(_08690_),
    .A(_08571_),
    .B(\hvsync_gen.vga.vpos[5] ));
 sg13g2_o21ai_1 _17009_ (.B1(_08690_),
    .Y(_08691_),
    .A1(\atari2600.tia.vid_ypos[3] ),
    .A2(_08573_));
 sg13g2_o21ai_1 _17010_ (.B1(_08682_),
    .Y(_08692_),
    .A1(_08689_),
    .A2(_08691_));
 sg13g2_nor2b_1 _17011_ (.A(\atari2600.tia.vid_ypos[6] ),
    .B_N(\hvsync_gen.vga.vpos[7] ),
    .Y(_08693_));
 sg13g2_nor2b_1 _17012_ (.A(\hvsync_gen.vga.vpos[7] ),
    .B_N(\atari2600.tia.vid_ypos[6] ),
    .Y(_08694_));
 sg13g2_nand2b_1 _17013_ (.Y(_08695_),
    .B(\atari2600.tia.vid_ypos[7] ),
    .A_N(\hvsync_gen.vga.vpos[8] ));
 sg13g2_o21ai_1 _17014_ (.B1(_08695_),
    .Y(_08696_),
    .A1(_08570_),
    .A2(\hvsync_gen.vga.vpos[6] ));
 sg13g2_or3_1 _17015_ (.A(_08693_),
    .B(_08694_),
    .C(_08696_),
    .X(_08697_));
 sg13g2_a21oi_1 _17016_ (.A1(_08681_),
    .A2(_08692_),
    .Y(_08698_),
    .B1(_08697_));
 sg13g2_nor2b_1 _17017_ (.A(\atari2600.tia.vid_ypos[7] ),
    .B_N(\hvsync_gen.vga.vpos[8] ),
    .Y(_08699_));
 sg13g2_o21ai_1 _17018_ (.B1(_08695_),
    .Y(_08700_),
    .A1(_08693_),
    .A2(_08699_));
 sg13g2_nor2_2 _17019_ (.A(\atari2600.tia.vid_ypos[7] ),
    .B(\atari2600.tia.vid_ypos[6] ),
    .Y(_08701_));
 sg13g2_or2_1 _17020_ (.X(_08702_),
    .B(\atari2600.tia.vid_ypos[0] ),
    .A(\atari2600.tia.vid_ypos[1] ));
 sg13g2_nand2_1 _17021_ (.Y(_08703_),
    .A(\atari2600.tia.vid_ypos[2] ),
    .B(_08702_));
 sg13g2_nor3_1 _17022_ (.A(_08570_),
    .B(\atari2600.tia.vid_ypos[4] ),
    .C(\atari2600.tia.vid_ypos[3] ),
    .Y(_08704_));
 sg13g2_a21o_1 _17023_ (.A2(_08704_),
    .A1(_08703_),
    .B1(_00070_),
    .X(_08705_));
 sg13g2_a21oi_1 _17024_ (.A1(_08701_),
    .A2(_08705_),
    .Y(_08706_),
    .B1(\hvsync_gen.vga.vpos[9] ));
 sg13g2_o21ai_1 _17025_ (.B1(_08700_),
    .Y(_08707_),
    .A1(\atari2600.tia.vid_ypos[8] ),
    .A2(_08706_));
 sg13g2_a22oi_1 _17026_ (.Y(_08708_),
    .B1(rom_data_pending),
    .B2(_08680_),
    .A2(_08572_),
    .A1(\atari2600.tia.vid_ypos[8] ));
 sg13g2_o21ai_1 _17027_ (.B1(_08708_),
    .Y(_08709_),
    .A1(_08698_),
    .A2(_08707_));
 sg13g2_inv_1 _17028_ (.Y(_08710_),
    .A(net5929));
 sg13g2_nor4_2 _17029_ (.A(net6246),
    .B(_08489_),
    .C(_08679_),
    .Y(_08711_),
    .D(net5929));
 sg13g2_nand2_2 _17030_ (.Y(_08712_),
    .A(_08680_),
    .B(_08710_));
 sg13g2_nor2_1 _17031_ (.A(\atari2600.stall_cpu ),
    .B(net5868),
    .Y(_08713_));
 sg13g2_nand2b_1 _17032_ (.Y(_08714_),
    .B(net5911),
    .A_N(\atari2600.stall_cpu ));
 sg13g2_nor2b_2 _17033_ (.A(net6513),
    .B_N(net6515),
    .Y(_08715_));
 sg13g2_nand2b_1 _17034_ (.Y(_08716_),
    .B(net6516),
    .A_N(net6514));
 sg13g2_nor2_1 _17035_ (.A(net6520),
    .B(net6521),
    .Y(_08717_));
 sg13g2_or2_2 _17036_ (.X(_08718_),
    .B(net6521),
    .A(net6520));
 sg13g2_nor2b_2 _17037_ (.A(net6519),
    .B_N(net6517),
    .Y(_08719_));
 sg13g2_nand2b_1 _17038_ (.Y(_08720_),
    .B(net6517),
    .A_N(net6519));
 sg13g2_nor3_2 _17039_ (.A(net6112),
    .B(_08718_),
    .C(net6109),
    .Y(_08721_));
 sg13g2_or4_2 _17040_ (.A(\atari2600.clk_counter[1] ),
    .B(_08489_),
    .C(_08679_),
    .D(net5929),
    .X(_08722_));
 sg13g2_nor2_1 _17041_ (.A(\atari2600.stall_cpu ),
    .B(_08722_),
    .Y(_08723_));
 sg13g2_or2_1 _17042_ (.X(_08724_),
    .B(_08722_),
    .A(\atari2600.stall_cpu ));
 sg13g2_mux2_1 _17043_ (.A0(\atari2600.cpu.DI[2] ),
    .A1(net7311),
    .S(net5866),
    .X(\atari2600.cpu.DIMUX[2] ));
 sg13g2_nor2b_1 _17044_ (.A(net6256),
    .B_N(net5827),
    .Y(_08725_));
 sg13g2_a21o_1 _17045_ (.A2(\atari2600.cpu.IRHOLD[2] ),
    .A1(net6256),
    .B1(_08725_),
    .X(_08726_));
 sg13g2_a21oi_2 _17046_ (.B1(_08725_),
    .Y(_08727_),
    .A2(\atari2600.cpu.IRHOLD[2] ),
    .A1(net6256));
 sg13g2_mux2_1 _17047_ (.A0(net7267),
    .A1(\atari2600.cpu.DIHOLD[3] ),
    .S(net5866),
    .X(\atari2600.cpu.DIMUX[3] ));
 sg13g2_nor2b_1 _17048_ (.A(net6254),
    .B_N(net5826),
    .Y(_08728_));
 sg13g2_a21o_1 _17049_ (.A2(\atari2600.cpu.IRHOLD[3] ),
    .A1(net6254),
    .B1(_08728_),
    .X(_08729_));
 sg13g2_a21oi_2 _17050_ (.B1(_08728_),
    .Y(_08730_),
    .A2(\atari2600.cpu.IRHOLD[3] ),
    .A1(net6254));
 sg13g2_mux2_2 _17051_ (.A0(_00082_),
    .A1(net7516),
    .S(net5867),
    .X(_08731_));
 sg13g2_inv_2 _17052_ (.Y(\atari2600.cpu.DIMUX[0] ),
    .A(net7517));
 sg13g2_nor2_1 _17053_ (.A(\atari2600.cpu.IRHOLD_valid ),
    .B(_08731_),
    .Y(_08732_));
 sg13g2_a21oi_2 _17054_ (.B1(_08732_),
    .Y(_08733_),
    .A2(\atari2600.cpu.IRHOLD[0] ),
    .A1(\atari2600.cpu.IRHOLD_valid ));
 sg13g2_and2_1 _17055_ (.A(_00079_),
    .B(net5866),
    .X(_08734_));
 sg13g2_a21o_2 _17056_ (.A2(net5835),
    .A1(net7574),
    .B1(_08734_),
    .X(_08735_));
 sg13g2_inv_4 _17057_ (.A(net7575),
    .Y(\atari2600.cpu.DIMUX[1] ));
 sg13g2_nor2_1 _17058_ (.A(net6255),
    .B(_08735_),
    .Y(_08736_));
 sg13g2_a21o_1 _17059_ (.A2(\atari2600.cpu.IRHOLD[1] ),
    .A1(net6255),
    .B1(_08736_),
    .X(_08737_));
 sg13g2_a21oi_2 _17060_ (.B1(_08736_),
    .Y(_08738_),
    .A2(\atari2600.cpu.IRHOLD[1] ),
    .A1(net6255));
 sg13g2_and2_1 _17061_ (.A(net5754),
    .B(_08738_),
    .X(_08739_));
 sg13g2_nand2_2 _17062_ (.Y(_08740_),
    .A(net5754),
    .B(_08738_));
 sg13g2_nor2_1 _17063_ (.A(_08727_),
    .B(_08740_),
    .Y(_08741_));
 sg13g2_nor3_2 _17064_ (.A(_08727_),
    .B(_08730_),
    .C(_08740_),
    .Y(_08742_));
 sg13g2_and2_1 _17065_ (.A(\atari2600.cpu.DIHOLD[7] ),
    .B(net5866),
    .X(_08743_));
 sg13g2_a21oi_2 _17066_ (.B1(_08743_),
    .Y(_08744_),
    .A2(net5835),
    .A1(\atari2600.cpu.DI[7] ));
 sg13g2_inv_4 _17067_ (.A(_08744_),
    .Y(\atari2600.cpu.DIMUX[7] ));
 sg13g2_nor2_1 _17068_ (.A(net6255),
    .B(_08744_),
    .Y(_08745_));
 sg13g2_a21o_2 _17069_ (.A2(\atari2600.cpu.IRHOLD[7] ),
    .A1(net6255),
    .B1(_08745_),
    .X(_08746_));
 sg13g2_a21oi_2 _17070_ (.B1(_08745_),
    .Y(_08747_),
    .A2(\atari2600.cpu.IRHOLD[7] ),
    .A1(net6255));
 sg13g2_and2_1 _17071_ (.A(\atari2600.cpu.DIHOLD[4] ),
    .B(net5865),
    .X(_08748_));
 sg13g2_a21oi_2 _17072_ (.B1(_08748_),
    .Y(_08749_),
    .A2(net5835),
    .A1(\atari2600.cpu.DI[4] ));
 sg13g2_inv_4 _17073_ (.A(_08749_),
    .Y(\atari2600.cpu.DIMUX[4] ));
 sg13g2_nor2_1 _17074_ (.A(net6254),
    .B(_08749_),
    .Y(_08750_));
 sg13g2_a21o_1 _17075_ (.A2(\atari2600.cpu.IRHOLD[4] ),
    .A1(net6254),
    .B1(_08750_),
    .X(_08751_));
 sg13g2_a21oi_1 _17076_ (.A1(net6254),
    .A2(\atari2600.cpu.IRHOLD[4] ),
    .Y(_08752_),
    .B1(_08750_));
 sg13g2_nor2_2 _17077_ (.A(_08746_),
    .B(net5735),
    .Y(_08753_));
 sg13g2_nand2_2 _17078_ (.Y(_08754_),
    .A(net5736),
    .B(net5733));
 sg13g2_mux2_1 _17079_ (.A0(net7299),
    .A1(\atari2600.cpu.DIHOLD[6] ),
    .S(net5866),
    .X(\atari2600.cpu.DIMUX[6] ));
 sg13g2_nor2b_1 _17080_ (.A(net6256),
    .B_N(net5825),
    .Y(_08755_));
 sg13g2_a21o_2 _17081_ (.A2(\atari2600.cpu.IRHOLD[6] ),
    .A1(net6256),
    .B1(_08755_),
    .X(_08756_));
 sg13g2_a21oi_2 _17082_ (.B1(_08755_),
    .Y(_08757_),
    .A2(\atari2600.cpu.IRHOLD[6] ),
    .A1(net6256));
 sg13g2_and2_1 _17083_ (.A(\atari2600.cpu.DIHOLD[5] ),
    .B(net5865),
    .X(_08758_));
 sg13g2_a21oi_2 _17084_ (.B1(_08758_),
    .Y(_08759_),
    .A2(net5835),
    .A1(\atari2600.cpu.DI[5] ));
 sg13g2_inv_4 _17085_ (.A(_08759_),
    .Y(\atari2600.cpu.DIMUX[5] ));
 sg13g2_nor2_1 _17086_ (.A(net6254),
    .B(_08759_),
    .Y(_08760_));
 sg13g2_a21o_2 _17087_ (.A2(net7036),
    .A1(net6254),
    .B1(_08760_),
    .X(_08761_));
 sg13g2_a21oi_2 _17088_ (.B1(_08760_),
    .Y(_08762_),
    .A2(net7036),
    .A1(net6255));
 sg13g2_nor2_2 _17089_ (.A(_08757_),
    .B(net5731),
    .Y(_08763_));
 sg13g2_nor2_1 _17090_ (.A(_08754_),
    .B(net5732),
    .Y(_08764_));
 sg13g2_nand3_1 _17091_ (.B(_08753_),
    .C(_08763_),
    .A(_08742_),
    .Y(_08765_));
 sg13g2_inv_1 _17092_ (.Y(_08766_),
    .A(_08765_));
 sg13g2_nor2_1 _17093_ (.A(net6515),
    .B(net6513),
    .Y(_08767_));
 sg13g2_or2_1 _17094_ (.X(_08768_),
    .B(net6514),
    .A(net6516));
 sg13g2_nand2_2 _17095_ (.Y(_08769_),
    .A(net6517),
    .B(net6519));
 sg13g2_nor3_1 _17096_ (.A(_08718_),
    .B(net6107),
    .C(_08769_),
    .Y(_08770_));
 sg13g2_nand4_1 _17097_ (.B(net6519),
    .C(net6110),
    .A(net6517),
    .Y(_08771_),
    .D(net6108));
 sg13g2_nor2_1 _17098_ (.A(net5858),
    .B(_08771_),
    .Y(_08772_));
 sg13g2_nand2_1 _17099_ (.Y(_08773_),
    .A(net5856),
    .B(net6035));
 sg13g2_nor2b_2 _17100_ (.A(net6515),
    .B_N(net6513),
    .Y(_08774_));
 sg13g2_nand2b_1 _17101_ (.Y(_08775_),
    .B(net6514),
    .A_N(net6516));
 sg13g2_nor2b_1 _17102_ (.A(net6517),
    .B_N(net6519),
    .Y(_08776_));
 sg13g2_nand2_2 _17103_ (.Y(_08777_),
    .A(net6520),
    .B(net6521));
 sg13g2_nand3_1 _17104_ (.B(net6521),
    .C(_08776_),
    .A(net6520),
    .Y(_08778_));
 sg13g2_nor2_1 _17105_ (.A(net6104),
    .B(_08778_),
    .Y(_08779_));
 sg13g2_nor2_1 _17106_ (.A(net5863),
    .B(net5999),
    .Y(_08780_));
 sg13g2_nand3_1 _17107_ (.B(_08719_),
    .C(_08774_),
    .A(net6110),
    .Y(_08781_));
 sg13g2_a21oi_1 _17108_ (.A1(net5866),
    .A2(_08781_),
    .Y(_08782_),
    .B1(_08780_));
 sg13g2_a221oi_1 _17109_ (.B2(net5823),
    .C1(_08782_),
    .B1(_08766_),
    .A1(net5866),
    .Y(_08783_),
    .A2(_08721_));
 sg13g2_nor2b_1 _17110_ (.A(net6520),
    .B_N(\atari2600.cpu.state[0] ),
    .Y(_08784_));
 sg13g2_nand2b_1 _17111_ (.Y(_08785_),
    .B(net6521),
    .A_N(net6520));
 sg13g2_nor2_1 _17112_ (.A(_08769_),
    .B(_08785_),
    .Y(_08786_));
 sg13g2_nand2b_1 _17113_ (.Y(_08787_),
    .B(net6102),
    .A_N(_08769_));
 sg13g2_nor2_1 _17114_ (.A(net6515),
    .B(_08787_),
    .Y(_08788_));
 sg13g2_a21oi_1 _17115_ (.A1(net6513),
    .A2(_08788_),
    .Y(_08789_),
    .B1(net5836));
 sg13g2_nand4_1 _17116_ (.B(net6519),
    .C(net6110),
    .A(net6517),
    .Y(_08790_),
    .D(_08774_));
 sg13g2_a21oi_1 _17117_ (.A1(net5836),
    .A2(_08790_),
    .Y(_08791_),
    .B1(_08789_));
 sg13g2_nand4_1 _17118_ (.B(net6519),
    .C(_08715_),
    .A(net6517),
    .Y(_08792_),
    .D(_08717_));
 sg13g2_nand3_1 _17119_ (.B(net5852),
    .C(_08786_),
    .A(_08715_),
    .Y(_08793_));
 sg13g2_o21ai_1 _17120_ (.B1(_08793_),
    .Y(_08794_),
    .A1(net5852),
    .A2(_08792_));
 sg13g2_nor2_2 _17121_ (.A(net6106),
    .B(_08787_),
    .Y(_08795_));
 sg13g2_nand2_2 _17122_ (.Y(_08796_),
    .A(net6108),
    .B(_08786_));
 sg13g2_nor2_2 _17123_ (.A(net6518),
    .B(net6519),
    .Y(_08797_));
 sg13g2_nand2_2 _17124_ (.Y(_08798_),
    .A(net6102),
    .B(_08797_));
 sg13g2_nand2_1 _17125_ (.Y(_08799_),
    .A(net6516),
    .B(net6513));
 sg13g2_nor2_2 _17126_ (.A(_08798_),
    .B(_08799_),
    .Y(_08800_));
 sg13g2_nor2_2 _17127_ (.A(_08769_),
    .B(_08777_),
    .Y(_08801_));
 sg13g2_nor3_2 _17128_ (.A(_08769_),
    .B(net6104),
    .C(_08777_),
    .Y(_08802_));
 sg13g2_nand2_1 _17129_ (.Y(_08803_),
    .A(_08774_),
    .B(_08801_));
 sg13g2_nand2_2 _17130_ (.Y(_08804_),
    .A(net6110),
    .B(net6103));
 sg13g2_nor2_2 _17131_ (.A(net6106),
    .B(_08804_),
    .Y(_08805_));
 sg13g2_nor2_2 _17132_ (.A(net6106),
    .B(_08798_),
    .Y(_08806_));
 sg13g2_nor4_2 _17133_ (.A(_08800_),
    .B(_08802_),
    .C(_08805_),
    .Y(_08807_),
    .D(_08806_));
 sg13g2_inv_1 _17134_ (.Y(_08808_),
    .A(_08807_));
 sg13g2_nor2b_1 _17135_ (.A(_08807_),
    .B_N(_00133_),
    .Y(_08809_));
 sg13g2_o21ai_1 _17136_ (.B1(_08786_),
    .Y(_08810_),
    .A1(_08715_),
    .A2(_08774_));
 sg13g2_nor2b_2 _17137_ (.A(net6521),
    .B_N(net6520),
    .Y(_08811_));
 sg13g2_nand2b_2 _17138_ (.Y(_08812_),
    .B(\atari2600.cpu.state[1] ),
    .A_N(\atari2600.cpu.state[0] ));
 sg13g2_nand2b_2 _17139_ (.Y(_08813_),
    .B(_08811_),
    .A_N(_08769_));
 sg13g2_nor2_2 _17140_ (.A(net6104),
    .B(_08813_),
    .Y(_08814_));
 sg13g2_or2_2 _17141_ (.X(_08815_),
    .B(_08813_),
    .A(net6104));
 sg13g2_nand2_1 _17142_ (.Y(_08816_),
    .A(net6103),
    .B(net6102));
 sg13g2_nand3_1 _17143_ (.B(net6103),
    .C(net6102),
    .A(_08715_),
    .Y(_08817_));
 sg13g2_nand3_1 _17144_ (.B(_08815_),
    .C(_08817_),
    .A(_08810_),
    .Y(_08818_));
 sg13g2_nor2_2 _17145_ (.A(net6111),
    .B(_08804_),
    .Y(_08819_));
 sg13g2_nor2_1 _17146_ (.A(net6247),
    .B(\atari2600.cpu.store ),
    .Y(_08820_));
 sg13g2_nand2b_1 _17147_ (.Y(_08821_),
    .B(_08797_),
    .A_N(_08777_));
 sg13g2_nor2_1 _17148_ (.A(net6106),
    .B(_08821_),
    .Y(_08822_));
 sg13g2_or2_1 _17149_ (.X(_08823_),
    .B(_08821_),
    .A(net6106));
 sg13g2_nor3_1 _17150_ (.A(\atari2600.cpu.ALU.CO ),
    .B(\atari2600.cpu.store ),
    .C(\atari2600.cpu.write_back ),
    .Y(_08824_));
 sg13g2_a22oi_1 _17151_ (.Y(_08825_),
    .B1(_08822_),
    .B2(_08824_),
    .A2(_08820_),
    .A1(_08819_));
 sg13g2_o21ai_1 _17152_ (.B1(_08825_),
    .Y(_08826_),
    .A1(net6111),
    .A2(_08798_));
 sg13g2_nor4_1 _17153_ (.A(net5861),
    .B(_08809_),
    .C(_08818_),
    .D(_08826_),
    .Y(_08827_));
 sg13g2_a21oi_1 _17154_ (.A1(net5852),
    .A2(_08796_),
    .Y(_08828_),
    .B1(_08827_));
 sg13g2_nor3_1 _17155_ (.A(_08791_),
    .B(_08794_),
    .C(_08828_),
    .Y(_08829_));
 sg13g2_nor2_2 _17156_ (.A(net5754),
    .B(_08737_),
    .Y(_08830_));
 sg13g2_nand2b_2 _17157_ (.Y(_08831_),
    .B(_08738_),
    .A_N(net5754));
 sg13g2_nand2_1 _17158_ (.Y(_08832_),
    .A(_08727_),
    .B(_08729_));
 sg13g2_nor2_1 _17159_ (.A(_08831_),
    .B(net5730),
    .Y(_08833_));
 sg13g2_nand2_1 _17160_ (.Y(_08834_),
    .A(net5754),
    .B(_08746_));
 sg13g2_nor2_1 _17161_ (.A(net5755),
    .B(_08729_),
    .Y(_08835_));
 sg13g2_nand2_2 _17162_ (.Y(_08836_),
    .A(_08727_),
    .B(_08730_));
 sg13g2_nor2_1 _17163_ (.A(_08834_),
    .B(_08836_),
    .Y(_08837_));
 sg13g2_nor2_1 _17164_ (.A(net5735),
    .B(net5818),
    .Y(_08838_));
 sg13g2_o21ai_1 _17165_ (.B1(net5733),
    .Y(_08839_),
    .A1(_08833_),
    .A2(_08837_));
 sg13g2_o21ai_1 _17166_ (.B1(_08829_),
    .Y(_08840_),
    .A1(net5821),
    .A2(_08839_));
 sg13g2_nor2_1 _17167_ (.A(_08727_),
    .B(_08729_),
    .Y(_08841_));
 sg13g2_a22oi_1 _17168_ (.Y(_08842_),
    .B1(_08838_),
    .B2(_08841_),
    .A2(_08802_),
    .A1(net5850));
 sg13g2_or2_1 _17169_ (.X(_08843_),
    .B(_08813_),
    .A(net6106));
 sg13g2_nand2_2 _17170_ (.Y(_08844_),
    .A(net6108),
    .B(_08801_));
 sg13g2_mux2_1 _17171_ (.A0(_08843_),
    .A1(_08844_),
    .S(net5862),
    .X(_08845_));
 sg13g2_nand2_1 _17172_ (.Y(_08846_),
    .A(_08842_),
    .B(_08845_));
 sg13g2_nand4_1 _17173_ (.B(\atari2600.cpu.state[0] ),
    .C(_08719_),
    .A(net6520),
    .Y(_08847_),
    .D(net6108));
 sg13g2_nor3_2 _17174_ (.A(net6514),
    .B(_08720_),
    .C(_08812_),
    .Y(_08848_));
 sg13g2_nor3_2 _17175_ (.A(net6109),
    .B(net6107),
    .C(_08812_),
    .Y(_08849_));
 sg13g2_nand3_1 _17176_ (.B(_08767_),
    .C(_08811_),
    .A(_08719_),
    .Y(_08850_));
 sg13g2_nor2_1 _17177_ (.A(net5864),
    .B(_08849_),
    .Y(_08851_));
 sg13g2_a21oi_1 _17178_ (.A1(net5864),
    .A2(_08847_),
    .Y(_08852_),
    .B1(_08851_));
 sg13g2_nor3_2 _17179_ (.A(net6112),
    .B(net6109),
    .C(_08812_),
    .Y(_08853_));
 sg13g2_nand2_1 _17180_ (.Y(_08854_),
    .A(net6516),
    .B(_08848_));
 sg13g2_nor3_2 _17181_ (.A(net6112),
    .B(net6109),
    .C(_08777_),
    .Y(_08855_));
 sg13g2_nor2_1 _17182_ (.A(net5836),
    .B(_08855_),
    .Y(_08856_));
 sg13g2_a21oi_1 _17183_ (.A1(net5836),
    .A2(_08854_),
    .Y(_08857_),
    .B1(_08856_));
 sg13g2_nor3_2 _17184_ (.A(net6109),
    .B(net6105),
    .C(_08812_),
    .Y(_08858_));
 sg13g2_nor3_2 _17185_ (.A(net6109),
    .B(net6105),
    .C(_08777_),
    .Y(_08859_));
 sg13g2_mux2_1 _17186_ (.A0(_08858_),
    .A1(_08859_),
    .S(net5863),
    .X(_08860_));
 sg13g2_nor3_1 _17187_ (.A(_08852_),
    .B(_08857_),
    .C(_08860_),
    .Y(_08861_));
 sg13g2_nand2_1 _17188_ (.Y(_08862_),
    .A(_08719_),
    .B(net6102));
 sg13g2_nor2_1 _17189_ (.A(net6105),
    .B(_08862_),
    .Y(_08863_));
 sg13g2_nor2_1 _17190_ (.A(net5836),
    .B(_08863_),
    .Y(_08864_));
 sg13g2_a21oi_1 _17191_ (.A1(net5834),
    .A2(_08781_),
    .Y(_08865_),
    .B1(_08864_));
 sg13g2_nand3_1 _17192_ (.B(_08719_),
    .C(net6102),
    .A(_08715_),
    .Y(_08866_));
 sg13g2_nand2_1 _17193_ (.Y(_08867_),
    .A(net5834),
    .B(_08721_));
 sg13g2_o21ai_1 _17194_ (.B1(_08867_),
    .Y(_08868_),
    .A1(net5834),
    .A2(_08866_));
 sg13g2_nor2_1 _17195_ (.A(net6107),
    .B(_08862_),
    .Y(_08869_));
 sg13g2_nand3_1 _17196_ (.B(net6108),
    .C(_08784_),
    .A(_08719_),
    .Y(_08870_));
 sg13g2_nand2_1 _17197_ (.Y(_08871_),
    .A(net5864),
    .B(_08869_));
 sg13g2_nor3_2 _17198_ (.A(_08718_),
    .B(net6109),
    .C(_08768_),
    .Y(_08872_));
 sg13g2_nand3_1 _17199_ (.B(_08719_),
    .C(net6108),
    .A(net6110),
    .Y(_08873_));
 sg13g2_o21ai_1 _17200_ (.B1(_08871_),
    .Y(_08874_),
    .A1(net5864),
    .A2(_08873_));
 sg13g2_nor3_1 _17201_ (.A(_08865_),
    .B(_08868_),
    .C(_08874_),
    .Y(_08875_));
 sg13g2_nand2_1 _17202_ (.Y(_08876_),
    .A(net5864),
    .B(_08850_));
 sg13g2_o21ai_1 _17203_ (.B1(_08876_),
    .Y(_08877_),
    .A1(net5864),
    .A2(_08869_));
 sg13g2_nor2_2 _17204_ (.A(net6111),
    .B(_08813_),
    .Y(_08878_));
 sg13g2_or2_1 _17205_ (.X(_08879_),
    .B(_08813_),
    .A(net6111));
 sg13g2_nor2_1 _17206_ (.A(net5862),
    .B(_08878_),
    .Y(_08880_));
 sg13g2_nand2_2 _17207_ (.Y(_08881_),
    .A(_08715_),
    .B(_08801_));
 sg13g2_a21oi_1 _17208_ (.A1(net5860),
    .A2(_08881_),
    .Y(_08882_),
    .B1(_08880_));
 sg13g2_inv_1 _17209_ (.Y(_08883_),
    .A(_08882_));
 sg13g2_nand4_1 _17210_ (.B(_08875_),
    .C(_08877_),
    .A(_08861_),
    .Y(_08884_),
    .D(_08883_));
 sg13g2_nor3_1 _17211_ (.A(_08840_),
    .B(_08846_),
    .C(_08884_),
    .Y(_08885_));
 sg13g2_nor2_2 _17212_ (.A(_08740_),
    .B(net5730),
    .Y(_08886_));
 sg13g2_or2_1 _17213_ (.X(_08887_),
    .B(net5730),
    .A(_08740_));
 sg13g2_nor2_2 _17214_ (.A(net5818),
    .B(_08887_),
    .Y(_08888_));
 sg13g2_a22oi_1 _17215_ (.Y(_08889_),
    .B1(_08888_),
    .B2(_08764_),
    .A2(_08878_),
    .A1(net5850));
 sg13g2_nor4_1 _17216_ (.A(net5735),
    .B(net5818),
    .C(_08831_),
    .D(_08836_),
    .Y(_08890_));
 sg13g2_or2_2 _17217_ (.X(_08891_),
    .B(_08821_),
    .A(net6104));
 sg13g2_nor2_1 _17218_ (.A(net5833),
    .B(_08814_),
    .Y(_08892_));
 sg13g2_a21oi_2 _17219_ (.B1(_08892_),
    .Y(_08893_),
    .A2(_08891_),
    .A1(net5833));
 sg13g2_o21ai_1 _17220_ (.B1(_08889_),
    .Y(_08894_),
    .A1(net5856),
    .A2(_08843_));
 sg13g2_nor3_1 _17221_ (.A(_08890_),
    .B(_08893_),
    .C(_08894_),
    .Y(_08895_));
 sg13g2_nor3_2 _17222_ (.A(_08754_),
    .B(_08756_),
    .C(net5732),
    .Y(_08896_));
 sg13g2_nor2_1 _17223_ (.A(_08740_),
    .B(_08836_),
    .Y(_08897_));
 sg13g2_nor3_1 _17224_ (.A(_08740_),
    .B(net5818),
    .C(_08836_),
    .Y(_08898_));
 sg13g2_a22oi_1 _17225_ (.Y(_08899_),
    .B1(_08896_),
    .B2(_08898_),
    .A2(_08853_),
    .A1(net5851));
 sg13g2_and3_1 _17226_ (.X(_08900_),
    .A(_08753_),
    .B(_08763_),
    .C(_08897_));
 sg13g2_a22oi_1 _17227_ (.Y(_08901_),
    .B1(_08900_),
    .B2(net5823),
    .A2(_08858_),
    .A1(net5850));
 sg13g2_and2_1 _17228_ (.A(_08899_),
    .B(_08901_),
    .X(_08902_));
 sg13g2_nand2_1 _17229_ (.Y(_08903_),
    .A(_08899_),
    .B(_08901_));
 sg13g2_nand4_1 _17230_ (.B(_08885_),
    .C(_08895_),
    .A(_08783_),
    .Y(_08904_),
    .D(_08902_));
 sg13g2_nor3_2 _17231_ (.A(_08754_),
    .B(_08757_),
    .C(_08761_),
    .Y(_08905_));
 sg13g2_nand2_1 _17232_ (.Y(_08906_),
    .A(_08742_),
    .B(_08905_));
 sg13g2_nand3_1 _17233_ (.B(net6035),
    .C(_08905_),
    .A(_08742_),
    .Y(_08907_));
 sg13g2_nand4_1 _17234_ (.B(_08847_),
    .C(_08866_),
    .A(net5835),
    .Y(_08908_),
    .D(_08907_));
 sg13g2_and2_1 _17235_ (.A(net6103),
    .B(_08811_),
    .X(_08909_));
 sg13g2_nand2_1 _17236_ (.Y(_08910_),
    .A(net6103),
    .B(_08811_));
 sg13g2_nor2_1 _17237_ (.A(net6112),
    .B(_08910_),
    .Y(_08911_));
 sg13g2_o21ai_1 _17238_ (.B1(_08908_),
    .Y(_08912_),
    .A1(net5834),
    .A2(_08911_));
 sg13g2_nor2_2 _17239_ (.A(net6104),
    .B(_08816_),
    .Y(_08913_));
 sg13g2_nand2_2 _17240_ (.Y(_08914_),
    .A(_08774_),
    .B(_08909_));
 sg13g2_nand2_1 _17241_ (.Y(_08915_),
    .A(net5862),
    .B(_08914_));
 sg13g2_o21ai_1 _17242_ (.B1(_08915_),
    .Y(_08916_),
    .A1(net5862),
    .A2(_08913_));
 sg13g2_nor2_1 _17243_ (.A(net6107),
    .B(_08910_),
    .Y(_08917_));
 sg13g2_nand2_1 _17244_ (.Y(_08918_),
    .A(_08767_),
    .B(_08909_));
 sg13g2_nor2_1 _17245_ (.A(net6107),
    .B(_08816_),
    .Y(_08919_));
 sg13g2_nand3_1 _17246_ (.B(net6103),
    .C(net6102),
    .A(net6108),
    .Y(_08920_));
 sg13g2_o21ai_1 _17247_ (.B1(_00056_),
    .Y(_08921_),
    .A1(\atari2600.cpu.cond_code[1] ),
    .A2(\atari2600.cpu.cond_code[0] ));
 sg13g2_nor2_1 _17248_ (.A(\atari2600.cpu.N ),
    .B(\atari2600.cpu.cond_code[2] ),
    .Y(_08922_));
 sg13g2_a21oi_1 _17249_ (.A1(_08582_),
    .A2(\atari2600.cpu.cond_code[2] ),
    .Y(_08923_),
    .B1(\atari2600.cpu.cond_code[1] ));
 sg13g2_o21ai_1 _17250_ (.B1(\atari2600.cpu.cond_code[1] ),
    .Y(_08924_),
    .A1(\atari2600.cpu.V ),
    .A2(_08670_));
 sg13g2_a21oi_1 _17251_ (.A1(_08578_),
    .A2(\atari2600.cpu.cond_code[2] ),
    .Y(_08925_),
    .B1(_08924_));
 sg13g2_nor3_1 _17252_ (.A(\atari2600.cpu.cond_code[0] ),
    .B(_08923_),
    .C(_08925_),
    .Y(_08926_));
 sg13g2_a22oi_1 _17253_ (.Y(_08927_),
    .B1(_00056_),
    .B2(\atari2600.cpu.V ),
    .A2(\atari2600.cpu.cond_code[2] ),
    .A1(\atari2600.cpu.Z ));
 sg13g2_nand2_1 _17254_ (.Y(_08928_),
    .A(\atari2600.cpu.cond_code[1] ),
    .B(_08927_));
 sg13g2_a221oi_1 _17255_ (.B2(_08660_),
    .C1(\atari2600.cpu.cond_code[1] ),
    .B1(_00056_),
    .A1(\atari2600.cpu.C ),
    .Y(_08929_),
    .A2(\atari2600.cpu.cond_code[2] ));
 sg13g2_nor2b_1 _17256_ (.A(_08929_),
    .B_N(\atari2600.cpu.cond_code[0] ),
    .Y(_08930_));
 sg13g2_a221oi_1 _17257_ (.B2(_08930_),
    .C1(_08926_),
    .B1(_08928_),
    .A1(_08921_),
    .Y(_08931_),
    .A2(_08922_));
 sg13g2_nor3_1 _17258_ (.A(net5861),
    .B(_08920_),
    .C(_08931_),
    .Y(_08932_));
 sg13g2_a21oi_2 _17259_ (.B1(_08932_),
    .Y(_08933_),
    .A2(net5995),
    .A1(net5861));
 sg13g2_nand4_1 _17260_ (.B(_08912_),
    .C(_08916_),
    .A(_08895_),
    .Y(_08934_),
    .D(_08933_));
 sg13g2_nor2_2 _17261_ (.A(net5733),
    .B(net5817),
    .Y(_08935_));
 sg13g2_nand3_1 _17262_ (.B(_08835_),
    .C(_08935_),
    .A(_08830_),
    .Y(_08936_));
 sg13g2_nand3_1 _17263_ (.B(_08797_),
    .C(_08811_),
    .A(_08715_),
    .Y(_08937_));
 sg13g2_o21ai_1 _17264_ (.B1(_08936_),
    .Y(_08938_),
    .A1(net5856),
    .A2(_08937_));
 sg13g2_nand3_1 _17265_ (.B(net6102),
    .C(_08797_),
    .A(_08774_),
    .Y(_08939_));
 sg13g2_nor4_2 _17266_ (.A(net6517),
    .B(\atari2600.cpu.state[2] ),
    .C(net6105),
    .Y(_08940_),
    .D(_08812_));
 sg13g2_nor2_1 _17267_ (.A(net5851),
    .B(_08939_),
    .Y(_08941_));
 sg13g2_a21oi_1 _17268_ (.A1(net5851),
    .A2(_08940_),
    .Y(_08942_),
    .B1(_08941_));
 sg13g2_nand3_1 _17269_ (.B(_08797_),
    .C(_08811_),
    .A(net6108),
    .Y(_08943_));
 sg13g2_a21o_1 _17270_ (.A2(_08870_),
    .A1(net5836),
    .B1(_08943_),
    .X(_08944_));
 sg13g2_a21oi_1 _17271_ (.A1(_08727_),
    .A2(_08831_),
    .Y(_08945_),
    .B1(_08730_));
 sg13g2_nand2_1 _17272_ (.Y(_08946_),
    .A(_08935_),
    .B(_08945_));
 sg13g2_nand4_1 _17273_ (.B(_08942_),
    .C(_08944_),
    .A(_08877_),
    .Y(_08947_),
    .D(_08946_));
 sg13g2_nor4_1 _17274_ (.A(_08903_),
    .B(_08934_),
    .C(_08938_),
    .D(_08947_),
    .Y(_08948_));
 sg13g2_a22oi_1 _17275_ (.Y(_08949_),
    .B1(_08913_),
    .B2(net5850),
    .A2(_08905_),
    .A1(_08898_));
 sg13g2_inv_1 _17276_ (.Y(_08950_),
    .A(_08949_));
 sg13g2_nand3b_1 _17277_ (.B(_08819_),
    .C(net5856),
    .Y(_08951_),
    .A_N(_08820_));
 sg13g2_o21ai_1 _17278_ (.B1(_08951_),
    .Y(_08952_),
    .A1(net5837),
    .A2(_08817_));
 sg13g2_nor3_1 _17279_ (.A(_08840_),
    .B(_08950_),
    .C(_08952_),
    .Y(_08953_));
 sg13g2_nand3_1 _17280_ (.B(net5732),
    .C(_08888_),
    .A(_08753_),
    .Y(_08954_));
 sg13g2_o21ai_1 _17281_ (.B1(_08954_),
    .Y(_08955_),
    .A1(net5856),
    .A2(_08939_));
 sg13g2_a22oi_1 _17282_ (.Y(_08956_),
    .B1(_08935_),
    .B2(_08897_),
    .A2(_08919_),
    .A1(net5850));
 sg13g2_nand2_2 _17283_ (.Y(_08957_),
    .A(net6110),
    .B(_08797_));
 sg13g2_nor2_2 _17284_ (.A(_08799_),
    .B(_08957_),
    .Y(_08958_));
 sg13g2_nand2b_1 _17285_ (.Y(_08959_),
    .B(net5857),
    .A_N(_08958_));
 sg13g2_o21ai_1 _17286_ (.B1(_08959_),
    .Y(_08960_),
    .A1(net5856),
    .A2(_08800_));
 sg13g2_nor2_2 _17287_ (.A(net6111),
    .B(_08957_),
    .Y(_08961_));
 sg13g2_o21ai_1 _17288_ (.B1(net5852),
    .Y(_08962_),
    .A1(net6111),
    .A2(_08798_));
 sg13g2_o21ai_1 _17289_ (.B1(_08962_),
    .Y(_08963_),
    .A1(net5852),
    .A2(_08961_));
 sg13g2_and2_1 _17290_ (.A(_08960_),
    .B(_08963_),
    .X(_08964_));
 sg13g2_nor3_1 _17291_ (.A(net5860),
    .B(net6106),
    .C(_08957_),
    .Y(_08965_));
 sg13g2_a21oi_1 _17292_ (.A1(net5860),
    .A2(_08806_),
    .Y(_08966_),
    .B1(_08965_));
 sg13g2_nand4_1 _17293_ (.B(_08956_),
    .C(_08964_),
    .A(_08875_),
    .Y(_08967_),
    .D(_08966_));
 sg13g2_nor2_1 _17294_ (.A(_08955_),
    .B(_08967_),
    .Y(_08968_));
 sg13g2_nor2_1 _17295_ (.A(net5834),
    .B(net5999),
    .Y(_08969_));
 sg13g2_a21oi_1 _17296_ (.A1(net5834),
    .A2(_08914_),
    .Y(_08970_),
    .B1(_08969_));
 sg13g2_nor2_1 _17297_ (.A(net6112),
    .B(_08778_),
    .Y(_08971_));
 sg13g2_mux2_1 _17298_ (.A0(_08911_),
    .A1(_08971_),
    .S(net5864),
    .X(_08972_));
 sg13g2_nor3_1 _17299_ (.A(_08846_),
    .B(_08970_),
    .C(_08972_),
    .Y(_08973_));
 sg13g2_nor2_2 _17300_ (.A(net6107),
    .B(_08778_),
    .Y(_08974_));
 sg13g2_or2_1 _17301_ (.X(_08975_),
    .B(_08778_),
    .A(net6107));
 sg13g2_xor2_1 _17302_ (.B(net6247),
    .A(\atari2600.cpu.backwards ),
    .X(_08976_));
 sg13g2_a21oi_1 _17303_ (.A1(net5995),
    .A2(_08976_),
    .Y(_08977_),
    .B1(net5865));
 sg13g2_a21oi_1 _17304_ (.A1(net5852),
    .A2(net5990),
    .Y(_08978_),
    .B1(_08977_));
 sg13g2_nor2_1 _17305_ (.A(_08882_),
    .B(_08978_),
    .Y(_08979_));
 sg13g2_or2_2 _17306_ (.X(_08980_),
    .B(_08821_),
    .A(net6111));
 sg13g2_and2_1 _17307_ (.A(net5860),
    .B(_08980_),
    .X(_08981_));
 sg13g2_a21oi_1 _17308_ (.A1(net5834),
    .A2(_08937_),
    .Y(_08982_),
    .B1(_08981_));
 sg13g2_or3_1 _17309_ (.A(_00133_),
    .B(net5860),
    .C(_08807_),
    .X(_08983_));
 sg13g2_o21ai_1 _17310_ (.B1(_08983_),
    .Y(_08984_),
    .A1(net5837),
    .A2(_08891_));
 sg13g2_nand2_1 _17311_ (.Y(_08985_),
    .A(net5860),
    .B(_08822_));
 sg13g2_o21ai_1 _17312_ (.B1(_08985_),
    .Y(_08986_),
    .A1(net5860),
    .A2(_08943_));
 sg13g2_nor3_1 _17313_ (.A(_08982_),
    .B(_08984_),
    .C(_08986_),
    .Y(_08987_));
 sg13g2_and4_1 _17314_ (.A(_08861_),
    .B(_08973_),
    .C(_08979_),
    .D(_08987_),
    .X(_08988_));
 sg13g2_nand3_1 _17315_ (.B(_08968_),
    .C(_08988_),
    .A(_08953_),
    .Y(_00171_));
 sg13g2_and2_2 _17316_ (.A(_08733_),
    .B(_08737_),
    .X(_08989_));
 sg13g2_nand2_1 _17317_ (.Y(_08990_),
    .A(net5754),
    .B(_08737_));
 sg13g2_nand2b_2 _17318_ (.Y(_08991_),
    .B(_08989_),
    .A_N(net5730));
 sg13g2_inv_1 _17319_ (.Y(_08992_),
    .A(_08991_));
 sg13g2_o21ai_1 _17320_ (.B1(_08991_),
    .Y(_08993_),
    .A1(_08753_),
    .A2(_08887_));
 sg13g2_nor2_2 _17321_ (.A(net6104),
    .B(_08804_),
    .Y(_08994_));
 sg13g2_nand3_1 _17322_ (.B(_08774_),
    .C(net6103),
    .A(net6110),
    .Y(_08995_));
 sg13g2_a22oi_1 _17323_ (.Y(_08996_),
    .B1(_08994_),
    .B2(net5850),
    .A2(_08993_),
    .A1(net5823));
 sg13g2_nor2_1 _17324_ (.A(net5852),
    .B(_08980_),
    .Y(_08997_));
 sg13g2_a21oi_1 _17325_ (.A1(net5852),
    .A2(_08819_),
    .Y(_08998_),
    .B1(_08997_));
 sg13g2_nor3_1 _17326_ (.A(net5860),
    .B(_08823_),
    .C(_08824_),
    .Y(_08999_));
 sg13g2_a21oi_1 _17327_ (.A1(net5861),
    .A2(_08805_),
    .Y(_09000_),
    .B1(_08999_));
 sg13g2_nand3_1 _17328_ (.B(_08998_),
    .C(_09000_),
    .A(_08996_),
    .Y(_09001_));
 sg13g2_nand3_1 _17329_ (.B(_08834_),
    .C(_08990_),
    .A(_08831_),
    .Y(_09002_));
 sg13g2_nand4_1 _17330_ (.B(_08729_),
    .C(net5733),
    .A(net5755),
    .Y(_09003_),
    .D(_09002_));
 sg13g2_nand2_2 _17331_ (.Y(_09004_),
    .A(_08741_),
    .B(_08896_));
 sg13g2_o21ai_1 _17332_ (.B1(_09003_),
    .Y(_09005_),
    .A1(_08730_),
    .A2(_09004_));
 sg13g2_a22oi_1 _17333_ (.Y(_09006_),
    .B1(_08958_),
    .B2(net5850),
    .A2(_08935_),
    .A1(_08841_));
 sg13g2_nor2_1 _17334_ (.A(net5862),
    .B(_08844_),
    .Y(_09007_));
 sg13g2_a21oi_1 _17335_ (.A1(net5850),
    .A2(_08961_),
    .Y(_09008_),
    .B1(_09007_));
 sg13g2_nand2_1 _17336_ (.Y(_09009_),
    .A(_09006_),
    .B(_09008_));
 sg13g2_nand2_1 _17337_ (.Y(_09010_),
    .A(net5834),
    .B(_08881_));
 sg13g2_nand3_1 _17338_ (.B(_08774_),
    .C(_08797_),
    .A(net6110),
    .Y(_09011_));
 sg13g2_nand2_1 _17339_ (.Y(_09012_),
    .A(net5863),
    .B(_09011_));
 sg13g2_o21ai_1 _17340_ (.B1(net5851),
    .Y(_09013_),
    .A1(net6516),
    .A2(_08957_));
 sg13g2_nand2_1 _17341_ (.Y(_09014_),
    .A(_09010_),
    .B(_09012_));
 sg13g2_a221oi_1 _17342_ (.B2(_09013_),
    .C1(_09009_),
    .B1(_09010_),
    .A1(net5823),
    .Y(_09015_),
    .A2(_09005_));
 sg13g2_nand2_1 _17343_ (.Y(_09016_),
    .A(_08783_),
    .B(_09015_));
 sg13g2_nor3_1 _17344_ (.A(_00171_),
    .B(_09001_),
    .C(_09016_),
    .Y(_09017_));
 sg13g2_nand2_1 _17345_ (.Y(_09018_),
    .A(net5734),
    .B(_08886_));
 sg13g2_nand4_1 _17346_ (.B(_08887_),
    .C(_08906_),
    .A(_08839_),
    .Y(_09019_),
    .D(_08991_));
 sg13g2_o21ai_1 _17347_ (.B1(_08730_),
    .Y(_09020_),
    .A1(net5755),
    .A2(_08830_));
 sg13g2_a21o_1 _17348_ (.A2(_08945_),
    .A1(net5735),
    .B1(_08900_),
    .X(_09021_));
 sg13g2_o21ai_1 _17349_ (.B1(net5733),
    .Y(_09022_),
    .A1(_08746_),
    .A2(_08763_));
 sg13g2_nand2_1 _17350_ (.Y(_09023_),
    .A(_08897_),
    .B(_09022_));
 sg13g2_nand3_1 _17351_ (.B(_09020_),
    .C(_09023_),
    .A(_08765_),
    .Y(_09024_));
 sg13g2_nor4_1 _17352_ (.A(_09005_),
    .B(_09019_),
    .C(_09021_),
    .D(_09024_),
    .Y(_09025_));
 sg13g2_o21ai_1 _17353_ (.B1(net6034),
    .Y(_09026_),
    .A1(net5862),
    .A2(_09025_));
 sg13g2_nand2_1 _17354_ (.Y(_09027_),
    .A(net5863),
    .B(_08792_));
 sg13g2_o21ai_1 _17355_ (.B1(_09027_),
    .Y(_09028_),
    .A1(net5863),
    .A2(_08855_));
 sg13g2_nand2_1 _17356_ (.Y(_09029_),
    .A(net5863),
    .B(_08790_));
 sg13g2_o21ai_1 _17357_ (.B1(_09029_),
    .Y(_09030_),
    .A1(net5863),
    .A2(_08859_));
 sg13g2_and2_1 _17358_ (.A(net5991),
    .B(_08931_),
    .X(_09031_));
 sg13g2_o21ai_1 _17359_ (.B1(_09011_),
    .Y(_09032_),
    .A1(net6513),
    .A2(_08778_));
 sg13g2_nor2_1 _17360_ (.A(net5992),
    .B(_08976_),
    .Y(_09033_));
 sg13g2_nor3_1 _17361_ (.A(_08795_),
    .B(_09032_),
    .C(_09033_),
    .Y(_09034_));
 sg13g2_nor4_1 _17362_ (.A(_08863_),
    .B(net6031),
    .C(_08994_),
    .D(_09031_),
    .Y(_09035_));
 sg13g2_a21o_1 _17363_ (.A2(_09035_),
    .A1(_09034_),
    .B1(net5863),
    .X(_09036_));
 sg13g2_nand4_1 _17364_ (.B(_09028_),
    .C(_09030_),
    .A(_09026_),
    .Y(_09037_),
    .D(_09036_));
 sg13g2_a21oi_1 _17365_ (.A1(_08948_),
    .A2(_09017_),
    .Y(_00176_),
    .B1(_08904_));
 sg13g2_or3_2 _17366_ (.A(net2983),
    .B(\flash_rom.fsm_state[1] ),
    .C(\flash_rom.fsm_state[0] ),
    .X(_09038_));
 sg13g2_inv_2 _17367_ (.Y(\flash_rom.spi_select ),
    .A(net2984));
 sg13g2_or2_1 _17368_ (.X(_09039_),
    .B(\hvsync_gen.vga.vpos[4] ),
    .A(\hvsync_gen.vga.vpos[5] ));
 sg13g2_nor4_1 _17369_ (.A(\hvsync_gen.vga.vpos[7] ),
    .B(\hvsync_gen.vga.vpos[6] ),
    .C(\hvsync_gen.vga.vpos[1] ),
    .D(_09039_),
    .Y(_09040_));
 sg13g2_nor4_1 _17370_ (.A(net7595),
    .B(\hvsync_gen.vga.vpos[8] ),
    .C(\hvsync_gen.vga.vpos[3] ),
    .D(\hvsync_gen.vga.vpos[2] ),
    .Y(_09041_));
 sg13g2_and2_2 _17371_ (.A(_09040_),
    .B(_09041_),
    .X(_00021_));
 sg13g2_nor2_1 _17372_ (.A(_08872_),
    .B(net6031),
    .Y(_09042_));
 sg13g2_nor2_2 _17373_ (.A(_08858_),
    .B(_08913_),
    .Y(_09043_));
 sg13g2_nand2_1 _17374_ (.Y(_09044_),
    .A(net5997),
    .B(_09043_));
 sg13g2_nand3_1 _17375_ (.B(_09042_),
    .C(_09043_),
    .A(net5997),
    .Y(_09045_));
 sg13g2_and3_1 _17376_ (.X(_09046_),
    .A(_08781_),
    .B(_08790_),
    .C(_08881_));
 sg13g2_nand4_1 _17377_ (.B(_08847_),
    .C(net5997),
    .A(_08792_),
    .Y(_09047_),
    .D(_09046_));
 sg13g2_or2_1 _17378_ (.X(_09048_),
    .B(_09047_),
    .A(net5940));
 sg13g2_nor4_1 _17379_ (.A(_00072_),
    .B(net6034),
    .C(_08878_),
    .D(_09048_),
    .Y(_09049_));
 sg13g2_nor2b_1 _17380_ (.A(_08958_),
    .B_N(_08980_),
    .Y(_09050_));
 sg13g2_nand3_1 _17381_ (.B(_08943_),
    .C(_09050_),
    .A(_08843_),
    .Y(_09051_));
 sg13g2_nor2_1 _17382_ (.A(_08577_),
    .B(_08771_),
    .Y(_09052_));
 sg13g2_nor3_2 _17383_ (.A(_09049_),
    .B(_09051_),
    .C(_09052_),
    .Y(_09053_));
 sg13g2_nor4_1 _17384_ (.A(net6035),
    .B(_08878_),
    .C(_09048_),
    .D(_09051_),
    .Y(_09054_));
 sg13g2_a22oi_1 _17385_ (.Y(_09055_),
    .B1(_09051_),
    .B2(\atari2600.cpu.index_y ),
    .A2(net6035),
    .A1(\atari2600.cpu.dst_reg[0] ));
 sg13g2_nand3b_1 _17386_ (.B(_09055_),
    .C(_08879_),
    .Y(_09056_),
    .A_N(_09048_));
 sg13g2_a21o_2 _17387_ (.A2(_09054_),
    .A1(_08575_),
    .B1(_09056_),
    .X(_09057_));
 sg13g2_nor2b_2 _17388_ (.A(_09053_),
    .B_N(_09057_),
    .Y(_09058_));
 sg13g2_nor2_2 _17389_ (.A(_09053_),
    .B(_09057_),
    .Y(_09059_));
 sg13g2_a22oi_1 _17390_ (.Y(_09060_),
    .B1(_09059_),
    .B2(\atari2600.cpu.AXYS[2][4] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][4] ));
 sg13g2_nor2b_2 _17391_ (.A(_09057_),
    .B_N(_09053_),
    .Y(_09061_));
 sg13g2_and2_2 _17392_ (.A(_09053_),
    .B(_09057_),
    .X(_09062_));
 sg13g2_a22oi_1 _17393_ (.Y(_09063_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][4] ),
    .A2(_09061_),
    .A1(\atari2600.cpu.AXYS[0][4] ));
 sg13g2_nand2_2 _17394_ (.Y(_09064_),
    .A(_09060_),
    .B(_09063_));
 sg13g2_nand2_1 _17395_ (.Y(_09065_),
    .A(_08803_),
    .B(_08937_));
 sg13g2_and2_2 _17396_ (.A(_08891_),
    .B(_08995_),
    .X(_09066_));
 sg13g2_nand3_1 _17397_ (.B(net5992),
    .C(_09066_),
    .A(_08815_),
    .Y(_09067_));
 sg13g2_nor2_1 _17398_ (.A(_08855_),
    .B(_08859_),
    .Y(_09068_));
 sg13g2_nor2b_1 _17399_ (.A(net5999),
    .B_N(_08844_),
    .Y(_09069_));
 sg13g2_nand2_1 _17400_ (.Y(_09070_),
    .A(_09068_),
    .B(_09069_));
 sg13g2_nand3_1 _17401_ (.B(_08870_),
    .C(_08914_),
    .A(_08850_),
    .Y(_09071_));
 sg13g2_or2_1 _17402_ (.X(_09072_),
    .B(_09071_),
    .A(_09070_));
 sg13g2_a21oi_1 _17403_ (.A1(net6112),
    .A2(net6104),
    .Y(_09073_),
    .B1(_08862_));
 sg13g2_nor2_2 _17404_ (.A(_08971_),
    .B(_09073_),
    .Y(_09074_));
 sg13g2_nand2b_1 _17405_ (.Y(_09075_),
    .B(_08823_),
    .A_N(_08819_));
 sg13g2_o21ai_1 _17406_ (.B1(_09074_),
    .Y(_09076_),
    .A1(net6513),
    .A2(_08798_));
 sg13g2_or2_1 _17407_ (.X(_09077_),
    .B(_09076_),
    .A(_09075_));
 sg13g2_inv_1 _17408_ (.Y(_09078_),
    .A(net5927));
 sg13g2_nor3_1 _17409_ (.A(_08800_),
    .B(_08961_),
    .C(net5928),
    .Y(_09079_));
 sg13g2_nand4_1 _17410_ (.B(_09046_),
    .C(_09078_),
    .A(_08980_),
    .Y(_09080_),
    .D(_09079_));
 sg13g2_nand3b_1 _17411_ (.B(_08817_),
    .C(net5990),
    .Y(_09081_),
    .A_N(_08805_));
 sg13g2_nor4_2 _17412_ (.A(net5940),
    .B(net5949),
    .C(_09080_),
    .Y(_09082_),
    .D(net5948));
 sg13g2_inv_1 _17413_ (.Y(_09083_),
    .A(_09082_));
 sg13g2_nor2_1 _17414_ (.A(net5939),
    .B(_09083_),
    .Y(_09084_));
 sg13g2_nand2b_2 _17415_ (.Y(_09085_),
    .B(_09082_),
    .A_N(net5939));
 sg13g2_nand3b_1 _17416_ (.B(_08815_),
    .C(_09066_),
    .Y(_09086_),
    .A_N(_09081_));
 sg13g2_nand2b_1 _17417_ (.Y(_09087_),
    .B(net5992),
    .A_N(_09080_));
 sg13g2_a221oi_1 _17418_ (.B2(net6250),
    .C1(net5751),
    .B1(_09087_),
    .A1(\atari2600.cpu.ABL[4] ),
    .Y(_09088_),
    .A2(_09086_));
 sg13g2_inv_1 _17419_ (.Y(_09089_),
    .A(_09088_));
 sg13g2_a221oi_1 _17420_ (.B2(\atari2600.cpu.DIMUX[4] ),
    .C1(_09089_),
    .B1(net5949),
    .A1(net5940),
    .Y(_09090_),
    .A2(_09064_));
 sg13g2_a21oi_2 _17421_ (.B1(_09090_),
    .Y(_09091_),
    .A2(net5750),
    .A1(_00085_));
 sg13g2_and2_1 _17422_ (.A(net5910),
    .B(_09091_),
    .X(_09092_));
 sg13g2_a21oi_2 _17423_ (.B1(_09092_),
    .Y(_09093_),
    .A2(_08722_),
    .A1(\atari2600.address_bus_r[4] ));
 sg13g2_a21o_1 _17424_ (.A2(_08722_),
    .A1(\atari2600.address_bus_r[4] ),
    .B1(_09092_),
    .X(_09094_));
 sg13g2_or2_1 _17425_ (.X(_09095_),
    .B(net5910),
    .A(\atari2600.address_bus_r[5] ));
 sg13g2_a22oi_1 _17426_ (.Y(_09096_),
    .B1(_09059_),
    .B2(\atari2600.cpu.AXYS[2][5] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][5] ));
 sg13g2_a22oi_1 _17427_ (.Y(_09097_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][5] ),
    .A2(_09061_),
    .A1(\atari2600.cpu.AXYS[0][5] ));
 sg13g2_nand2_2 _17428_ (.Y(_09098_),
    .A(_09096_),
    .B(_09097_));
 sg13g2_nand2_1 _17429_ (.Y(_09099_),
    .A(net5940),
    .B(_09098_));
 sg13g2_a22oi_1 _17430_ (.Y(_09100_),
    .B1(_09086_),
    .B2(\atari2600.cpu.ABL[5] ),
    .A2(net5994),
    .A1(_08596_));
 sg13g2_nand2_1 _17431_ (.Y(_09101_),
    .A(_09085_),
    .B(_09100_));
 sg13g2_a221oi_1 _17432_ (.B2(net6249),
    .C1(_09101_),
    .B1(_09080_),
    .A1(\atari2600.cpu.DIMUX[5] ),
    .Y(_09102_),
    .A2(net5949));
 sg13g2_a22oi_1 _17433_ (.Y(_09103_),
    .B1(_09099_),
    .B2(_09102_),
    .A2(net5750),
    .A1(_08595_));
 sg13g2_o21ai_1 _17434_ (.B1(_09095_),
    .Y(_09104_),
    .A1(net5868),
    .A2(_09103_));
 sg13g2_and2_2 _17435_ (.A(net5282),
    .B(net5572),
    .X(_09105_));
 sg13g2_nand2_1 _17436_ (.Y(_09106_),
    .A(net5279),
    .B(net5569));
 sg13g2_nand2b_1 _17437_ (.Y(_09107_),
    .B(_08870_),
    .A_N(_08855_));
 sg13g2_or4_1 _17438_ (.A(_08848_),
    .B(_08872_),
    .C(net6031),
    .D(net5989),
    .X(_09108_));
 sg13g2_nand2b_1 _17439_ (.Y(_09109_),
    .B(_08815_),
    .A_N(_09108_));
 sg13g2_inv_2 _17440_ (.Y(_09110_),
    .A(net5938));
 sg13g2_nor3_1 _17441_ (.A(net6518),
    .B(net6111),
    .C(_08785_),
    .Y(_09111_));
 sg13g2_o21ai_1 _17442_ (.B1(\atari2600.cpu.store ),
    .Y(_09112_),
    .A1(_08808_),
    .A2(_09111_));
 sg13g2_o21ai_1 _17443_ (.B1(_09112_),
    .Y(_09113_),
    .A1(\atari2600.cpu.res ),
    .A2(_09110_));
 sg13g2_a22oi_1 _17444_ (.Y(_09114_),
    .B1(_09061_),
    .B2(\atari2600.cpu.AXYS[0][7] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][7] ));
 sg13g2_a22oi_1 _17445_ (.Y(_09115_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][7] ),
    .A2(_09059_),
    .A1(\atari2600.cpu.AXYS[2][7] ));
 sg13g2_nand2_1 _17446_ (.Y(_09116_),
    .A(_09114_),
    .B(_09115_));
 sg13g2_nand2_1 _17447_ (.Y(_09117_),
    .A(net5940),
    .B(_09116_));
 sg13g2_a22oi_1 _17448_ (.Y(_09118_),
    .B1(_09086_),
    .B2(\atari2600.cpu.ABL[7] ),
    .A2(net5994),
    .A1(_08599_));
 sg13g2_a22oi_1 _17449_ (.Y(_09119_),
    .B1(_09080_),
    .B2(\atari2600.cpu.ADD[7] ),
    .A2(net5949),
    .A1(\atari2600.cpu.DIMUX[7] ));
 sg13g2_nand4_1 _17450_ (.B(_09117_),
    .C(_09118_),
    .A(_09085_),
    .Y(_09120_),
    .D(_09119_));
 sg13g2_o21ai_1 _17451_ (.B1(_09120_),
    .Y(_09121_),
    .A1(\atari2600.cpu.PC[7] ),
    .A2(_09085_));
 sg13g2_nand2_1 _17452_ (.Y(_09122_),
    .A(\atari2600.cpu.DIMUX[4] ),
    .B(net5927));
 sg13g2_a221oi_1 _17453_ (.B2(net6250),
    .C1(net5751),
    .B1(net5948),
    .A1(\atari2600.cpu.ABH[4] ),
    .Y(_09123_),
    .A2(net5939));
 sg13g2_a22oi_1 _17454_ (.Y(_09124_),
    .B1(_09122_),
    .B2(_09123_),
    .A2(net5750),
    .A1(_08598_));
 sg13g2_nor2_2 _17455_ (.A(net5869),
    .B(_09124_),
    .Y(_09125_));
 sg13g2_nand3_1 _17456_ (.B(_09121_),
    .C(_09125_),
    .A(_09113_),
    .Y(_09126_));
 sg13g2_nor2_2 _17457_ (.A(net5272),
    .B(_09126_),
    .Y(_09127_));
 sg13g2_or2_2 _17458_ (.X(_09128_),
    .B(_09126_),
    .A(net5271));
 sg13g2_mux4_1 _17459_ (.S0(_09057_),
    .A0(\atari2600.cpu.AXYS[2][1] ),
    .A1(\atari2600.cpu.AXYS[3][1] ),
    .A2(\atari2600.cpu.AXYS[0][1] ),
    .A3(\atari2600.cpu.AXYS[1][1] ),
    .S1(_09053_),
    .X(_09129_));
 sg13g2_nor2_1 _17460_ (.A(_00074_),
    .B(_08918_),
    .Y(_09130_));
 sg13g2_a221oi_1 _17461_ (.B2(\atari2600.cpu.ABL[1] ),
    .C1(_09130_),
    .B1(_09086_),
    .A1(net6252),
    .Y(_09131_),
    .A2(_09080_));
 sg13g2_nand2_1 _17462_ (.Y(_09132_),
    .A(_09085_),
    .B(_09131_));
 sg13g2_a221oi_1 _17463_ (.B2(_09045_),
    .C1(_09132_),
    .B1(_09129_),
    .A1(\atari2600.cpu.DIMUX[1] ),
    .Y(_09133_),
    .A2(_09065_));
 sg13g2_a21oi_2 _17464_ (.B1(_09133_),
    .Y(_09134_),
    .A2(net5752),
    .A1(_00088_));
 sg13g2_mux2_2 _17465_ (.A0(\atari2600.address_bus_r[1] ),
    .A1(_09134_),
    .S(net5911),
    .X(_09135_));
 sg13g2_or2_1 _17466_ (.X(_09136_),
    .B(net5911),
    .A(\atari2600.address_bus_r[2] ));
 sg13g2_a22oi_1 _17467_ (.Y(_09137_),
    .B1(_09061_),
    .B2(\atari2600.cpu.AXYS[0][2] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][2] ));
 sg13g2_a22oi_1 _17468_ (.Y(_09138_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][2] ),
    .A2(_09059_),
    .A1(\atari2600.cpu.AXYS[2][2] ));
 sg13g2_nand2_2 _17469_ (.Y(_09139_),
    .A(_09137_),
    .B(_09138_));
 sg13g2_nor2_1 _17470_ (.A(_00076_),
    .B(net5992),
    .Y(_09140_));
 sg13g2_a221oi_1 _17471_ (.B2(\atari2600.cpu.ABL[2] ),
    .C1(_09140_),
    .B1(_09086_),
    .A1(net6251),
    .Y(_09141_),
    .A2(_09080_));
 sg13g2_nand2_1 _17472_ (.Y(_09142_),
    .A(_09085_),
    .B(_09141_));
 sg13g2_a221oi_1 _17473_ (.B2(net5940),
    .C1(_09142_),
    .B1(_09139_),
    .A1(net5827),
    .Y(_09143_),
    .A2(net5949));
 sg13g2_a21oi_2 _17474_ (.B1(_09143_),
    .Y(_09144_),
    .A2(net5752),
    .A1(_00078_));
 sg13g2_mux2_1 _17475_ (.A0(\atari2600.address_bus_r[2] ),
    .A1(_09144_),
    .S(net5911),
    .X(_09145_));
 sg13g2_o21ai_1 _17476_ (.B1(_09136_),
    .Y(_09146_),
    .A1(net5868),
    .A2(_09144_));
 sg13g2_nor2_2 _17477_ (.A(net5566),
    .B(net5558),
    .Y(_09147_));
 sg13g2_mux4_1 _17478_ (.S0(_09057_),
    .A0(\atari2600.cpu.AXYS[2][0] ),
    .A1(\atari2600.cpu.AXYS[3][0] ),
    .A2(\atari2600.cpu.AXYS[0][0] ),
    .A3(\atari2600.cpu.AXYS[1][0] ),
    .S1(_09053_),
    .X(_09148_));
 sg13g2_a22oi_1 _17479_ (.Y(_09149_),
    .B1(_09087_),
    .B2(\atari2600.cpu.ADD[0] ),
    .A2(_09086_),
    .A1(\atari2600.cpu.ABL[0] ));
 sg13g2_nand2_1 _17480_ (.Y(_09150_),
    .A(_09085_),
    .B(_09149_));
 sg13g2_a221oi_1 _17481_ (.B2(_09045_),
    .C1(_09150_),
    .B1(_09148_),
    .A1(\atari2600.cpu.DIMUX[0] ),
    .Y(_09151_),
    .A2(net5949));
 sg13g2_a21oi_2 _17482_ (.B1(_09151_),
    .Y(_09152_),
    .A2(net5752),
    .A1(_00087_));
 sg13g2_and2_1 _17483_ (.A(net5911),
    .B(_09152_),
    .X(_09153_));
 sg13g2_a21oi_1 _17484_ (.A1(net7579),
    .A2(_08722_),
    .Y(_09154_),
    .B1(_09153_));
 sg13g2_a21o_1 _17485_ (.A2(_08722_),
    .A1(\atari2600.address_bus_r[0] ),
    .B1(_09153_),
    .X(_09155_));
 sg13g2_or2_1 _17486_ (.X(_09156_),
    .B(net5910),
    .A(\atari2600.address_bus_r[3] ));
 sg13g2_a22oi_1 _17487_ (.Y(_09157_),
    .B1(_09061_),
    .B2(\atari2600.cpu.AXYS[0][3] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][3] ));
 sg13g2_a22oi_1 _17488_ (.Y(_09158_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][3] ),
    .A2(_09059_),
    .A1(\atari2600.cpu.AXYS[2][3] ));
 sg13g2_nand2_2 _17489_ (.Y(_09159_),
    .A(_09157_),
    .B(_09158_));
 sg13g2_nor2_1 _17490_ (.A(_00090_),
    .B(net5992),
    .Y(_09160_));
 sg13g2_a221oi_1 _17491_ (.B2(\atari2600.cpu.ABL[3] ),
    .C1(_09160_),
    .B1(_09086_),
    .A1(\atari2600.cpu.ADD[3] ),
    .Y(_09161_),
    .A2(_09080_));
 sg13g2_nand2_1 _17492_ (.Y(_09162_),
    .A(_09085_),
    .B(_09161_));
 sg13g2_a221oi_1 _17493_ (.B2(net5940),
    .C1(_09162_),
    .B1(_09159_),
    .A1(net5826),
    .Y(_09163_),
    .A2(net5949));
 sg13g2_a21oi_2 _17494_ (.B1(_09163_),
    .Y(_09164_),
    .A2(net5750),
    .A1(_00089_));
 sg13g2_mux2_1 _17495_ (.A0(\atari2600.address_bus_r[3] ),
    .A1(_09164_),
    .S(net5910),
    .X(_09165_));
 sg13g2_o21ai_1 _17496_ (.B1(_09156_),
    .Y(_09166_),
    .A1(net5868),
    .A2(_09164_));
 sg13g2_nand2_1 _17497_ (.Y(_09167_),
    .A(net5528),
    .B(net5550));
 sg13g2_nor2_2 _17498_ (.A(net5567),
    .B(net5532),
    .Y(_09168_));
 sg13g2_nand2b_2 _17499_ (.Y(_09169_),
    .B(net5527),
    .A_N(net5565));
 sg13g2_nor2_2 _17500_ (.A(net5558),
    .B(net5553),
    .Y(_09170_));
 sg13g2_nand2_2 _17501_ (.Y(_09171_),
    .A(net5563),
    .B(net5548));
 sg13g2_nor2_2 _17502_ (.A(_09169_),
    .B(net5524),
    .Y(_09172_));
 sg13g2_and2_2 _17503_ (.A(_09127_),
    .B(_09172_),
    .X(_09173_));
 sg13g2_nand2_2 _17504_ (.Y(_09174_),
    .A(net6563),
    .B(_09173_));
 sg13g2_nor2_1 _17505_ (.A(_09109_),
    .B(_09129_),
    .Y(_09175_));
 sg13g2_nand2b_1 _17506_ (.Y(_09176_),
    .B(net6031),
    .A_N(\atari2600.cpu.php ));
 sg13g2_nand2_2 _17507_ (.Y(_09177_),
    .A(_08815_),
    .B(_09176_));
 sg13g2_nand2b_1 _17508_ (.Y(_09178_),
    .B(_09177_),
    .A_N(_00074_));
 sg13g2_a21oi_2 _17509_ (.B1(_08849_),
    .Y(_09179_),
    .A2(net6031),
    .A1(\atari2600.cpu.php ));
 sg13g2_or2_1 _17510_ (.X(_09180_),
    .B(_09179_),
    .A(_00073_));
 sg13g2_nand2_2 _17511_ (.Y(_09181_),
    .A(net5997),
    .B(_08873_));
 sg13g2_a22oi_1 _17512_ (.Y(_09182_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[9] ),
    .A2(_09107_),
    .A1(\atari2600.cpu.PC[1] ));
 sg13g2_nand4_1 _17513_ (.B(_09178_),
    .C(_09180_),
    .A(net5938),
    .Y(_09183_),
    .D(_09182_));
 sg13g2_nor2b_1 _17514_ (.A(_09175_),
    .B_N(_09183_),
    .Y(_09184_));
 sg13g2_o21ai_1 _17515_ (.B1(_09183_),
    .Y(_09185_),
    .A1(net5938),
    .A2(_09129_));
 sg13g2_nor2_1 _17516_ (.A(net5937),
    .B(_09139_),
    .Y(_09186_));
 sg13g2_or2_1 _17517_ (.X(_09187_),
    .B(_09179_),
    .A(_00075_));
 sg13g2_nand2b_1 _17518_ (.Y(_09188_),
    .B(_09177_),
    .A_N(_00076_));
 sg13g2_a22oi_1 _17519_ (.Y(_09189_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[10] ),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[2] ));
 sg13g2_nand4_1 _17520_ (.B(_09187_),
    .C(_09188_),
    .A(net5938),
    .Y(_09190_),
    .D(_09189_));
 sg13g2_nor2b_1 _17521_ (.A(_09186_),
    .B_N(_09190_),
    .Y(_09191_));
 sg13g2_o21ai_1 _17522_ (.B1(_09190_),
    .Y(_09192_),
    .A1(net5936),
    .A2(_09139_));
 sg13g2_nor2_1 _17523_ (.A(net5938),
    .B(_09148_),
    .Y(_09193_));
 sg13g2_nand3_1 _17524_ (.B(\atari2600.cpu.C ),
    .C(net6031),
    .A(\atari2600.cpu.php ),
    .Y(_09194_));
 sg13g2_o21ai_1 _17525_ (.B1(_09194_),
    .Y(_09195_),
    .A1(_00077_),
    .A2(_08850_));
 sg13g2_a21oi_1 _17526_ (.A1(\atari2600.cpu.PC[0] ),
    .A2(net5989),
    .Y(_09196_),
    .B1(_09195_));
 sg13g2_a22oi_1 _17527_ (.Y(_09197_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[8] ),
    .A2(_09177_),
    .A1(\atari2600.cpu.ADD[0] ));
 sg13g2_nand3_1 _17528_ (.B(_09196_),
    .C(_09197_),
    .A(net5938),
    .Y(_09198_));
 sg13g2_nor2b_2 _17529_ (.A(_09193_),
    .B_N(_09198_),
    .Y(_09199_));
 sg13g2_o21ai_1 _17530_ (.B1(_09198_),
    .Y(_09200_),
    .A1(net5938),
    .A2(_09148_));
 sg13g2_nand2_1 _17531_ (.Y(_09201_),
    .A(net5728),
    .B(net5743));
 sg13g2_xnor2_1 _17532_ (.Y(_09202_),
    .A(net5726),
    .B(net5743));
 sg13g2_nor2_2 _17533_ (.A(net5797),
    .B(net5743),
    .Y(_09203_));
 sg13g2_a22oi_1 _17534_ (.Y(_09204_),
    .B1(_09203_),
    .B2(net5726),
    .A2(_09202_),
    .A1(net5797));
 sg13g2_nor2_1 _17535_ (.A(net6535),
    .B(_09173_),
    .Y(_09205_));
 sg13g2_nand2_1 _17536_ (.Y(_09206_),
    .A(net4293),
    .B(net5079));
 sg13g2_o21ai_1 _17537_ (.B1(_09206_),
    .Y(_00020_),
    .A1(net5080),
    .A2(_09204_));
 sg13g2_nand2_1 _17538_ (.Y(_09207_),
    .A(net5748),
    .B(_09202_));
 sg13g2_nand2_1 _17539_ (.Y(_09208_),
    .A(net4429),
    .B(net5079));
 sg13g2_o21ai_1 _17540_ (.B1(_09208_),
    .Y(_00019_),
    .A1(net5080),
    .A2(_09207_));
 sg13g2_nor2_1 _17541_ (.A(net5564),
    .B(net5529),
    .Y(_09209_));
 sg13g2_nand2b_2 _17542_ (.Y(_09210_),
    .B(net5530),
    .A_N(net5566));
 sg13g2_nor2_2 _17543_ (.A(net5524),
    .B(_09210_),
    .Y(_09211_));
 sg13g2_nand2_2 _17544_ (.Y(_09212_),
    .A(_09170_),
    .B(net5402));
 sg13g2_nor2_2 _17545_ (.A(_09128_),
    .B(_09212_),
    .Y(_09213_));
 sg13g2_nand2_2 _17546_ (.Y(_09214_),
    .A(_09127_),
    .B(_09211_));
 sg13g2_nand2_2 _17547_ (.Y(_09215_),
    .A(net6561),
    .B(_09213_));
 sg13g2_nor2_2 _17548_ (.A(net6533),
    .B(_09213_),
    .Y(_09216_));
 sg13g2_nand2_1 _17549_ (.Y(_09217_),
    .A(net2979),
    .B(_09216_));
 sg13g2_o21ai_1 _17550_ (.B1(_09217_),
    .Y(_00018_),
    .A1(_09204_),
    .A2(_09215_));
 sg13g2_nand2_1 _17551_ (.Y(_09218_),
    .A(net3439),
    .B(_09216_));
 sg13g2_o21ai_1 _17552_ (.B1(_09218_),
    .Y(_00017_),
    .A1(_09207_),
    .A2(_09215_));
 sg13g2_nor2_1 _17553_ (.A(net2932),
    .B(\flash_rom.spi_select ),
    .Y(_00000_));
 sg13g2_nor2_2 _17554_ (.A(_08655_),
    .B(net6126),
    .Y(_09219_));
 sg13g2_nand2_2 _17555_ (.Y(_09220_),
    .A(net6125),
    .B(_08656_));
 sg13g2_and2_1 _17556_ (.A(\hvsync_gen.hpos[5] ),
    .B(net6134),
    .X(_09221_));
 sg13g2_nand2_1 _17557_ (.Y(_09222_),
    .A(net6133),
    .B(net6134));
 sg13g2_nand2_2 _17558_ (.Y(_09223_),
    .A(net6132),
    .B(\hvsync_gen.hpos[7] ));
 sg13g2_or2_1 _17559_ (.X(_09224_),
    .B(_09223_),
    .A(_09222_));
 sg13g2_a21oi_1 _17560_ (.A1(_09219_),
    .A2(_09224_),
    .Y(_09225_),
    .B1(net7569));
 sg13g2_nor2_2 _17561_ (.A(\hvsync_gen.hpos[7] ),
    .B(net6126),
    .Y(_09226_));
 sg13g2_nor2_2 _17562_ (.A(_08655_),
    .B(_09226_),
    .Y(_09227_));
 sg13g2_o21ai_1 _17563_ (.B1(net6125),
    .Y(_09228_),
    .A1(\hvsync_gen.hpos[7] ),
    .A2(net6126));
 sg13g2_nor2_1 _17564_ (.A(net6133),
    .B(net6134),
    .Y(_09229_));
 sg13g2_or2_1 _17565_ (.X(_09230_),
    .B(\hvsync_gen.hpos[4] ),
    .A(net6133));
 sg13g2_nor2_1 _17566_ (.A(net6129),
    .B(net6075),
    .Y(_09231_));
 sg13g2_nor3_1 _17567_ (.A(net6129),
    .B(net6126),
    .C(net6075),
    .Y(_09232_));
 sg13g2_nor3_2 _17568_ (.A(_09225_),
    .B(net6087),
    .C(_09232_),
    .Y(_00055_));
 sg13g2_nand4_1 _17569_ (.B(\hvsync_gen.vga.vpos[7] ),
    .C(\hvsync_gen.vga.vpos[6] ),
    .A(\hvsync_gen.vga.vpos[8] ),
    .Y(_09233_),
    .D(\hvsync_gen.vga.vpos[5] ));
 sg13g2_nor2_1 _17570_ (.A(\atari2600.tia.vblank ),
    .B(\hvsync_gen.vga.vpos[9] ),
    .Y(_09234_));
 sg13g2_nand3_1 _17571_ (.B(_09233_),
    .C(_09234_),
    .A(_09228_),
    .Y(_09235_));
 sg13g2_xor2_1 _17572_ (.B(\hvsync_gen.vga.vpos[0] ),
    .A(\frame_counter[0] ),
    .X(_09236_));
 sg13g2_xnor2_1 _17573_ (.Y(_09237_),
    .A(\frame_counter[0] ),
    .B(\hvsync_gen.vga.vpos[0] ));
 sg13g2_nand2_1 _17574_ (.Y(_09238_),
    .A(\b_pwm_odd[8] ),
    .B(_09237_));
 sg13g2_nand2_1 _17575_ (.Y(_09239_),
    .A(\b_pwm_even[8] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17576_ (.B1(_09235_),
    .Y(uo_out[6]),
    .A2(_09239_),
    .A1(_09238_));
 sg13g2_nand2_1 _17577_ (.Y(_09240_),
    .A(\b_pwm_odd[9] ),
    .B(_09237_));
 sg13g2_nand2_1 _17578_ (.Y(_09241_),
    .A(\b_pwm_even[9] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17579_ (.B1(_09235_),
    .Y(uo_out[2]),
    .A2(_09241_),
    .A1(_09240_));
 sg13g2_nand2_1 _17580_ (.Y(_09242_),
    .A(\g_pwm_odd[8] ),
    .B(_09237_));
 sg13g2_nand2_1 _17581_ (.Y(_09243_),
    .A(\g_pwm_even[8] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17582_ (.B1(_09235_),
    .Y(uo_out[5]),
    .A2(_09243_),
    .A1(_09242_));
 sg13g2_nand2_1 _17583_ (.Y(_09244_),
    .A(\g_pwm_odd[9] ),
    .B(_09237_));
 sg13g2_nand2_1 _17584_ (.Y(_09245_),
    .A(\g_pwm_even[9] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17585_ (.B1(_09235_),
    .Y(uo_out[1]),
    .A2(_09245_),
    .A1(_09244_));
 sg13g2_nand2_1 _17586_ (.Y(_09246_),
    .A(\r_pwm_odd[8] ),
    .B(_09237_));
 sg13g2_nand2_1 _17587_ (.Y(_09247_),
    .A(\r_pwm_even[8] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17588_ (.B1(_09235_),
    .Y(uo_out[4]),
    .A2(_09247_),
    .A1(_09246_));
 sg13g2_nand2_1 _17589_ (.Y(_09248_),
    .A(\r_pwm_odd[9] ),
    .B(_09237_));
 sg13g2_nand2_1 _17590_ (.Y(_09249_),
    .A(\r_pwm_even[9] ),
    .B(_09236_));
 sg13g2_a21oi_2 _17591_ (.B1(_09235_),
    .Y(uo_out[0]),
    .A2(_09249_),
    .A1(_09248_));
 sg13g2_or2_1 _17592_ (.X(_09250_),
    .B(net5910),
    .A(\atari2600.address_bus_r[6] ));
 sg13g2_a22oi_1 _17593_ (.Y(_09251_),
    .B1(_09062_),
    .B2(\atari2600.cpu.AXYS[1][6] ),
    .A2(_09058_),
    .A1(\atari2600.cpu.AXYS[3][6] ));
 sg13g2_a22oi_1 _17594_ (.Y(_09252_),
    .B1(_09061_),
    .B2(\atari2600.cpu.AXYS[0][6] ),
    .A2(_09059_),
    .A1(\atari2600.cpu.AXYS[2][6] ));
 sg13g2_nand2_2 _17595_ (.Y(_09253_),
    .A(_09251_),
    .B(_09252_));
 sg13g2_nor2_1 _17596_ (.A(_00092_),
    .B(net5992),
    .Y(_09254_));
 sg13g2_a221oi_1 _17597_ (.B2(\atari2600.cpu.ABL[6] ),
    .C1(_09254_),
    .B1(_09086_),
    .A1(net6248),
    .Y(_09255_),
    .A2(_09080_));
 sg13g2_nand2_1 _17598_ (.Y(_09256_),
    .A(_09085_),
    .B(_09255_));
 sg13g2_a221oi_1 _17599_ (.B2(net5940),
    .C1(_09256_),
    .B1(_09253_),
    .A1(net5825),
    .Y(_09257_),
    .A2(net5949));
 sg13g2_a21oi_2 _17600_ (.B1(_09257_),
    .Y(_09258_),
    .A2(net5750),
    .A1(_08593_));
 sg13g2_mux2_1 _17601_ (.A0(\atari2600.address_bus_r[6] ),
    .A1(_09258_),
    .S(net5910),
    .X(_09259_));
 sg13g2_o21ai_1 _17602_ (.B1(_09250_),
    .Y(_09260_),
    .A1(net5868),
    .A2(_09258_));
 sg13g2_nor2_2 _17603_ (.A(net5571),
    .B(_09260_),
    .Y(_09261_));
 sg13g2_nor2_2 _17604_ (.A(net5283),
    .B(net5551),
    .Y(_09262_));
 sg13g2_nand2_1 _17605_ (.Y(_09263_),
    .A(net5277),
    .B(net5553));
 sg13g2_and2_2 _17606_ (.A(_09261_),
    .B(_09262_),
    .X(_09264_));
 sg13g2_nand2_2 _17607_ (.Y(_09265_),
    .A(_09261_),
    .B(_09262_));
 sg13g2_nand2_1 _17608_ (.Y(_09266_),
    .A(\atari2600.address_bus_r[7] ),
    .B(net5868));
 sg13g2_o21ai_1 _17609_ (.B1(_09266_),
    .Y(_09267_),
    .A1(net5868),
    .A2(_09121_));
 sg13g2_nand2_1 _17610_ (.Y(_09268_),
    .A(\atari2600.cpu.DIMUX[0] ),
    .B(_09077_));
 sg13g2_a221oi_1 _17611_ (.B2(net6253),
    .C1(net5753),
    .B1(_09081_),
    .A1(\atari2600.cpu.ABH[0] ),
    .Y(_09269_),
    .A2(_09067_));
 sg13g2_a22oi_1 _17612_ (.Y(_09270_),
    .B1(_09268_),
    .B2(_09269_),
    .A2(net5752),
    .A1(_08584_));
 sg13g2_nor2b_1 _17613_ (.A(net5910),
    .B_N(net7585),
    .Y(_09271_));
 sg13g2_a21oi_2 _17614_ (.B1(_09271_),
    .Y(_09272_),
    .A2(_09270_),
    .A1(net5910));
 sg13g2_nand2_1 _17615_ (.Y(_09273_),
    .A(\atari2600.cpu.DIMUX[1] ),
    .B(net5927));
 sg13g2_a221oi_1 _17616_ (.B2(net6252),
    .C1(net5752),
    .B1(net5948),
    .A1(\atari2600.cpu.ABH[1] ),
    .Y(_09274_),
    .A2(_09067_));
 sg13g2_a22oi_1 _17617_ (.Y(_09275_),
    .B1(_09273_),
    .B2(_09274_),
    .A2(net5752),
    .A1(_08579_));
 sg13g2_nor2_2 _17618_ (.A(net5869),
    .B(_09275_),
    .Y(_09276_));
 sg13g2_a21oi_2 _17619_ (.B1(_09276_),
    .Y(_09277_),
    .A2(_08722_),
    .A1(_08603_));
 sg13g2_inv_2 _17620_ (.Y(_09278_),
    .A(_09277_));
 sg13g2_nand2_1 _17621_ (.Y(_09279_),
    .A(net5827),
    .B(net5927));
 sg13g2_a221oi_1 _17622_ (.B2(net6251),
    .C1(net5752),
    .B1(net5948),
    .A1(\atari2600.cpu.ABH[2] ),
    .Y(_09280_),
    .A2(net5939));
 sg13g2_a22oi_1 _17623_ (.Y(_09281_),
    .B1(_09279_),
    .B2(_09280_),
    .A2(net5752),
    .A1(_08581_));
 sg13g2_or2_1 _17624_ (.X(_09282_),
    .B(net5912),
    .A(\atari2600.address_bus_r[10] ));
 sg13g2_o21ai_1 _17625_ (.B1(_09282_),
    .Y(_09283_),
    .A1(net5868),
    .A2(_09281_));
 sg13g2_nor3_2 _17626_ (.A(_09272_),
    .B(_09278_),
    .C(_09283_),
    .Y(_09284_));
 sg13g2_nand4_1 _17627_ (.B(_09264_),
    .C(_09267_),
    .A(net5562),
    .Y(_09285_),
    .D(_09284_));
 sg13g2_nand2_1 _17628_ (.Y(_09286_),
    .A(net5826),
    .B(net5927));
 sg13g2_a221oi_1 _17629_ (.B2(\atari2600.cpu.ADD[3] ),
    .C1(net5751),
    .B1(net5948),
    .A1(\atari2600.cpu.ABH[3] ),
    .Y(_09287_),
    .A2(net5939));
 sg13g2_a22oi_1 _17630_ (.Y(_09288_),
    .B1(_09286_),
    .B2(_09287_),
    .A2(net5751),
    .A1(_08605_));
 sg13g2_mux2_1 _17631_ (.A0(\atari2600.address_bus_r[11] ),
    .A1(_09288_),
    .S(net5911),
    .X(_09289_));
 sg13g2_nand2_1 _17632_ (.Y(_09290_),
    .A(_09285_),
    .B(net5540));
 sg13g2_nor2_2 _17633_ (.A(net5561),
    .B(net5552),
    .Y(_09291_));
 sg13g2_nand2_1 _17634_ (.Y(_09292_),
    .A(net5560),
    .B(_09166_));
 sg13g2_nor2_2 _17635_ (.A(net5281),
    .B(_09291_),
    .Y(_09293_));
 sg13g2_o21ai_1 _17636_ (.B1(net5277),
    .Y(_09294_),
    .A1(net5530),
    .A2(net5504));
 sg13g2_nor2_2 _17637_ (.A(net5566),
    .B(net5561),
    .Y(_09295_));
 sg13g2_o21ai_1 _17638_ (.B1(net5553),
    .Y(_09296_),
    .A1(net5402),
    .A2(_09295_));
 sg13g2_a21oi_1 _17639_ (.A1(_09294_),
    .A2(_09296_),
    .Y(_09297_),
    .B1(net5572));
 sg13g2_and2_2 _17640_ (.A(net5564),
    .B(net5529),
    .X(_09298_));
 sg13g2_nand2_2 _17641_ (.Y(_09299_),
    .A(net5567),
    .B(net5528));
 sg13g2_nand3_1 _17642_ (.B(_09263_),
    .C(net5338),
    .A(net5572),
    .Y(_09300_));
 sg13g2_nor2_2 _17643_ (.A(net5276),
    .B(net5571),
    .Y(_09301_));
 sg13g2_or2_1 _17644_ (.X(_09302_),
    .B(net5572),
    .A(net5276));
 sg13g2_nand2_2 _17645_ (.Y(_09303_),
    .A(net5567),
    .B(net5562));
 sg13g2_and2_2 _17646_ (.A(net5564),
    .B(net5532),
    .X(_09304_));
 sg13g2_nand2_2 _17647_ (.Y(_09305_),
    .A(net5567),
    .B(net5532));
 sg13g2_nor2_2 _17648_ (.A(net5517),
    .B(_09305_),
    .Y(_09306_));
 sg13g2_nand2_2 _17649_ (.Y(_09307_),
    .A(_09170_),
    .B(net5309));
 sg13g2_o21ai_1 _17650_ (.B1(_09300_),
    .Y(_09308_),
    .A1(net5268),
    .A2(_09307_));
 sg13g2_o21ai_1 _17651_ (.B1(net5547),
    .Y(_09309_),
    .A1(_09297_),
    .A2(_09308_));
 sg13g2_nand2_1 _17652_ (.Y(_09310_),
    .A(_09293_),
    .B(net5338));
 sg13g2_nor2_2 _17653_ (.A(net5565),
    .B(net5549),
    .Y(_09311_));
 sg13g2_nor2_2 _17654_ (.A(net5557),
    .B(net5527),
    .Y(_09312_));
 sg13g2_nor3_1 _17655_ (.A(net5357),
    .B(_09311_),
    .C(_09312_),
    .Y(_09313_));
 sg13g2_nor2_2 _17656_ (.A(net5558),
    .B(net5549),
    .Y(_09314_));
 sg13g2_nand2_2 _17657_ (.Y(_09315_),
    .A(net5562),
    .B(net5556));
 sg13g2_o21ai_1 _17658_ (.B1(net5280),
    .Y(_09316_),
    .A1(net5309),
    .A2(net5491));
 sg13g2_o21ai_1 _17659_ (.B1(_09310_),
    .Y(_09317_),
    .A1(_09313_),
    .A2(_09316_));
 sg13g2_nor2_2 _17660_ (.A(net5569),
    .B(net5547),
    .Y(_09318_));
 sg13g2_and2_2 _17661_ (.A(net5277),
    .B(_09104_),
    .X(_09319_));
 sg13g2_nand2_1 _17662_ (.Y(_09320_),
    .A(net5277),
    .B(net5572));
 sg13g2_nor2_2 _17663_ (.A(net5546),
    .B(net5264),
    .Y(_09321_));
 sg13g2_nand2_2 _17664_ (.Y(_09322_),
    .A(net5542),
    .B(_09319_));
 sg13g2_and2_1 _17665_ (.A(net5567),
    .B(net5554),
    .X(_09323_));
 sg13g2_nand2_1 _17666_ (.Y(_09324_),
    .A(net5565),
    .B(_09314_));
 sg13g2_o21ai_1 _17667_ (.B1(_09324_),
    .Y(_09325_),
    .A1(net5530),
    .A2(_09314_));
 sg13g2_nand3_1 _17668_ (.B(_09278_),
    .C(_09283_),
    .A(_09272_),
    .Y(_09326_));
 sg13g2_nor2_2 _17669_ (.A(_09267_),
    .B(_09326_),
    .Y(_09327_));
 sg13g2_nor2_1 _17670_ (.A(net5270),
    .B(net5550),
    .Y(_09328_));
 sg13g2_nor2_2 _17671_ (.A(net5272),
    .B(net5544),
    .Y(_09329_));
 sg13g2_nand2_2 _17672_ (.Y(_09330_),
    .A(_09105_),
    .B(net5542));
 sg13g2_nand2_2 _17673_ (.Y(_09331_),
    .A(net5552),
    .B(_09329_));
 sg13g2_nor3_1 _17674_ (.A(net5404),
    .B(_09295_),
    .C(_09331_),
    .Y(_09332_));
 sg13g2_a21oi_1 _17675_ (.A1(_09321_),
    .A2(_09325_),
    .Y(_09333_),
    .B1(_09332_));
 sg13g2_nand3_1 _17676_ (.B(_09327_),
    .C(_09333_),
    .A(_09309_),
    .Y(_09334_));
 sg13g2_a21oi_1 _17677_ (.A1(_09317_),
    .A2(_09318_),
    .Y(_09335_),
    .B1(_09334_));
 sg13g2_o21ai_1 _17678_ (.B1(_09290_),
    .Y(_00009_),
    .A1(net5540),
    .A2(_09335_));
 sg13g2_a21oi_2 _17679_ (.B1(net5552),
    .Y(_09336_),
    .A2(net5356),
    .A1(net5561));
 sg13g2_nor2_2 _17680_ (.A(net5561),
    .B(net5384),
    .Y(_09337_));
 sg13g2_nand2_2 _17681_ (.Y(_09338_),
    .A(net5559),
    .B(net5405));
 sg13g2_nand2_2 _17682_ (.Y(_09339_),
    .A(net5530),
    .B(net5552));
 sg13g2_nor2_2 _17683_ (.A(net5561),
    .B(net5549),
    .Y(_09340_));
 sg13g2_nand2_1 _17684_ (.Y(_09341_),
    .A(net5559),
    .B(net5554));
 sg13g2_nor2_2 _17685_ (.A(net5561),
    .B(_09339_),
    .Y(_09342_));
 sg13g2_nand2_2 _17686_ (.Y(_09343_),
    .A(net5415),
    .B(_09340_));
 sg13g2_o21ai_1 _17687_ (.B1(net5278),
    .Y(_09344_),
    .A1(_09336_),
    .A2(_09337_));
 sg13g2_and2_2 _17688_ (.A(net5572),
    .B(net5545),
    .X(_09345_));
 sg13g2_inv_1 _17689_ (.Y(_09346_),
    .A(_09345_));
 sg13g2_a21oi_1 _17690_ (.A1(net5282),
    .A2(net5338),
    .Y(_09347_),
    .B1(_09346_));
 sg13g2_nand2_1 _17691_ (.Y(_09348_),
    .A(_09344_),
    .B(_09347_));
 sg13g2_nor2_2 _17692_ (.A(net5562),
    .B(_09305_),
    .Y(_09349_));
 sg13g2_nand2_2 _17693_ (.Y(_09350_),
    .A(net5559),
    .B(net5310));
 sg13g2_nor3_1 _17694_ (.A(net5558),
    .B(net5449),
    .C(_09323_),
    .Y(_09351_));
 sg13g2_o21ai_1 _17695_ (.B1(_09329_),
    .Y(_09352_),
    .A1(_09349_),
    .A2(_09351_));
 sg13g2_nor2_2 _17696_ (.A(net5559),
    .B(net5432),
    .Y(_09353_));
 sg13g2_and2_1 _17697_ (.A(net5565),
    .B(net5557),
    .X(_09354_));
 sg13g2_nand2_2 _17698_ (.Y(_09355_),
    .A(net5565),
    .B(net5557));
 sg13g2_a21oi_1 _17699_ (.A1(_09147_),
    .A2(net5552),
    .Y(_09356_),
    .B1(net5527));
 sg13g2_a22oi_1 _17700_ (.Y(_09357_),
    .B1(_09355_),
    .B2(_09356_),
    .A2(_09314_),
    .A1(net5449));
 sg13g2_nand2_2 _17701_ (.Y(_09358_),
    .A(_09167_),
    .B(_09339_));
 sg13g2_a21oi_1 _17702_ (.A1(net5566),
    .A2(_09358_),
    .Y(_09359_),
    .B1(_09353_));
 sg13g2_o21ai_1 _17703_ (.B1(_09294_),
    .Y(_09360_),
    .A1(net5278),
    .A2(_09359_));
 sg13g2_nand2b_2 _17704_ (.Y(_09361_),
    .B(net5276),
    .A_N(net5571));
 sg13g2_a221oi_1 _17705_ (.B2(_09350_),
    .C1(_09361_),
    .B1(_09336_),
    .A1(net5553),
    .Y(_09362_),
    .A2(net5338));
 sg13g2_nand2_2 _17706_ (.Y(_09363_),
    .A(net5303),
    .B(_09340_));
 sg13g2_nor2_2 _17707_ (.A(net5268),
    .B(_09363_),
    .Y(_09364_));
 sg13g2_or2_2 _17708_ (.X(_09365_),
    .B(_09363_),
    .A(net5269));
 sg13g2_nor3_1 _17709_ (.A(net5504),
    .B(net5268),
    .C(net5309),
    .Y(_09366_));
 sg13g2_nor3_1 _17710_ (.A(_09362_),
    .B(_09364_),
    .C(_09366_),
    .Y(_09367_));
 sg13g2_o21ai_1 _17711_ (.B1(_09367_),
    .Y(_09368_),
    .A1(net5264),
    .A2(_09357_));
 sg13g2_a22oi_1 _17712_ (.Y(_09369_),
    .B1(_09368_),
    .B2(net5542),
    .A2(_09360_),
    .A1(_09261_));
 sg13g2_and4_1 _17713_ (.A(_09327_),
    .B(_09348_),
    .C(_09352_),
    .D(_09369_),
    .X(_09370_));
 sg13g2_o21ai_1 _17714_ (.B1(_09290_),
    .Y(_00010_),
    .A1(net5540),
    .A2(_09370_));
 sg13g2_nor2_2 _17715_ (.A(net5402),
    .B(net5356),
    .Y(_09371_));
 sg13g2_nand2_1 _17716_ (.Y(_09372_),
    .A(net5384),
    .B(net5338));
 sg13g2_a21oi_1 _17717_ (.A1(_09291_),
    .A2(_09371_),
    .Y(_09373_),
    .B1(net5282));
 sg13g2_o21ai_1 _17718_ (.B1(_09373_),
    .Y(_09374_),
    .A1(net5384),
    .A2(_09291_));
 sg13g2_a21oi_1 _17719_ (.A1(net5531),
    .A2(_09311_),
    .Y(_09375_),
    .B1(net5278));
 sg13g2_nand2_2 _17720_ (.Y(_09376_),
    .A(net5566),
    .B(_09312_));
 sg13g2_a21oi_1 _17721_ (.A1(_09375_),
    .A2(_09376_),
    .Y(_09377_),
    .B1(net5570));
 sg13g2_nor3_1 _17722_ (.A(net5531),
    .B(_09311_),
    .C(net5264),
    .Y(_09378_));
 sg13g2_a221oi_1 _17723_ (.B2(_09377_),
    .C1(_09378_),
    .B1(_09374_),
    .A1(_09328_),
    .Y(_09379_),
    .A2(_09353_));
 sg13g2_nor2_1 _17724_ (.A(net5544),
    .B(_09379_),
    .Y(_09380_));
 sg13g2_o21ai_1 _17725_ (.B1(net5550),
    .Y(_09381_),
    .A1(_09147_),
    .A2(net5404));
 sg13g2_o21ai_1 _17726_ (.B1(_09375_),
    .Y(_09382_),
    .A1(_09312_),
    .A2(_09381_));
 sg13g2_nor3_1 _17727_ (.A(net5282),
    .B(net5552),
    .C(net5449),
    .Y(_09383_));
 sg13g2_and2_1 _17728_ (.A(net5557),
    .B(_09383_),
    .X(_09384_));
 sg13g2_nor2_1 _17729_ (.A(net5569),
    .B(_09384_),
    .Y(_09385_));
 sg13g2_nand4_1 _17730_ (.B(net5550),
    .C(_09319_),
    .A(net5531),
    .Y(_09386_),
    .D(_09355_));
 sg13g2_a22oi_1 _17731_ (.Y(_09387_),
    .B1(_09382_),
    .B2(_09385_),
    .A2(net5404),
    .A1(_09105_));
 sg13g2_a21oi_1 _17732_ (.A1(_09386_),
    .A2(_09387_),
    .Y(_09388_),
    .B1(net5543));
 sg13g2_nor4_1 _17733_ (.A(net5514),
    .B(_09326_),
    .C(_09380_),
    .D(_09388_),
    .Y(_09389_));
 sg13g2_o21ai_1 _17734_ (.B1(_09290_),
    .Y(_00011_),
    .A1(net5540),
    .A2(_09389_));
 sg13g2_nor3_1 _17735_ (.A(net5561),
    .B(net5531),
    .C(_09323_),
    .Y(_09390_));
 sg13g2_nor2_1 _17736_ (.A(net5268),
    .B(_09390_),
    .Y(_09391_));
 sg13g2_nor3_1 _17737_ (.A(net5552),
    .B(_09301_),
    .C(_09355_),
    .Y(_09392_));
 sg13g2_nand3_1 _17738_ (.B(net5553),
    .C(net5338),
    .A(net5571),
    .Y(_09393_));
 sg13g2_a21oi_1 _17739_ (.A1(net5557),
    .A2(net5530),
    .Y(_09394_),
    .B1(_09393_));
 sg13g2_nor4_1 _17740_ (.A(net5546),
    .B(_09319_),
    .C(_09392_),
    .D(_09394_),
    .Y(_09395_));
 sg13g2_a22oi_1 _17741_ (.Y(_09396_),
    .B1(_09391_),
    .B2(_09212_),
    .A2(_09372_),
    .A1(_09293_));
 sg13g2_nand2_2 _17742_ (.Y(_09397_),
    .A(net5281),
    .B(_09261_));
 sg13g2_nor2_2 _17743_ (.A(_09305_),
    .B(net5493),
    .Y(_09398_));
 sg13g2_a221oi_1 _17744_ (.B2(_09170_),
    .C1(_09398_),
    .B1(_09371_),
    .A1(net5565),
    .Y(_09399_),
    .A2(_09291_));
 sg13g2_a22oi_1 _17745_ (.Y(_09400_),
    .B1(_09383_),
    .B2(_09350_),
    .A2(_09372_),
    .A1(net5282));
 sg13g2_nor2_2 _17746_ (.A(net5508),
    .B(net5338),
    .Y(_09401_));
 sg13g2_nor2_1 _17747_ (.A(_09361_),
    .B(_09401_),
    .Y(_09402_));
 sg13g2_nor2_1 _17748_ (.A(net5432),
    .B(net5485),
    .Y(_09403_));
 sg13g2_nand2_2 _17749_ (.Y(_09404_),
    .A(net5443),
    .B(_09340_));
 sg13g2_o21ai_1 _17750_ (.B1(_09327_),
    .Y(_09405_),
    .A1(_09322_),
    .A2(_09404_));
 sg13g2_a221oi_1 _17751_ (.B2(net5546),
    .C1(_09405_),
    .B1(_09402_),
    .A1(_09345_),
    .Y(_09406_),
    .A2(_09400_));
 sg13g2_o21ai_1 _17752_ (.B1(_09406_),
    .Y(_09407_),
    .A1(_09397_),
    .A2(_09399_));
 sg13g2_a21oi_1 _17753_ (.A1(_09395_),
    .A2(_09396_),
    .Y(_09408_),
    .B1(_09407_));
 sg13g2_o21ai_1 _17754_ (.B1(_09290_),
    .Y(_00012_),
    .A1(net5540),
    .A2(_09408_));
 sg13g2_o21ai_1 _17755_ (.B1(_09212_),
    .Y(_09409_),
    .A1(net5339),
    .A2(net5499));
 sg13g2_nor2_1 _17756_ (.A(net5267),
    .B(_09343_),
    .Y(_09410_));
 sg13g2_a21oi_2 _17757_ (.B1(_09410_),
    .Y(_09411_),
    .A2(_09409_),
    .A1(_09301_));
 sg13g2_nor2_2 _17758_ (.A(_09260_),
    .B(_09411_),
    .Y(_09412_));
 sg13g2_nor2_2 _17759_ (.A(net5554),
    .B(_09330_),
    .Y(_09413_));
 sg13g2_nand2_2 _17760_ (.Y(_09414_),
    .A(net5548),
    .B(_09329_));
 sg13g2_o21ai_1 _17761_ (.B1(_09329_),
    .Y(_09415_),
    .A1(net5549),
    .A2(_09371_));
 sg13g2_nor2b_1 _17762_ (.A(_09295_),
    .B_N(_09336_),
    .Y(_09416_));
 sg13g2_nor3_1 _17763_ (.A(_09314_),
    .B(_09415_),
    .C(_09416_),
    .Y(_09417_));
 sg13g2_nand2_1 _17764_ (.Y(_09418_),
    .A(_09261_),
    .B(_09373_));
 sg13g2_nand2_2 _17765_ (.Y(_09419_),
    .A(_09327_),
    .B(_09418_));
 sg13g2_nand2_2 _17766_ (.Y(_09420_),
    .A(net5279),
    .B(_09318_));
 sg13g2_inv_4 _17767_ (.A(_09420_),
    .Y(_09421_));
 sg13g2_nand2_2 _17768_ (.Y(_09422_),
    .A(net5549),
    .B(_09421_));
 sg13g2_nand2_1 _17769_ (.Y(_09423_),
    .A(_09318_),
    .B(_09384_));
 sg13g2_o21ai_1 _17770_ (.B1(_09423_),
    .Y(_09424_),
    .A1(_09355_),
    .A2(_09422_));
 sg13g2_nor4_2 _17771_ (.A(_09412_),
    .B(_09417_),
    .C(_09419_),
    .Y(_09425_),
    .D(_09424_));
 sg13g2_o21ai_1 _17772_ (.B1(net5540),
    .Y(_09426_),
    .A1(net5527),
    .A2(_09285_));
 sg13g2_o21ai_1 _17773_ (.B1(_09426_),
    .Y(_00013_),
    .A1(net5541),
    .A2(_09425_));
 sg13g2_nor3_1 _17774_ (.A(_09147_),
    .B(net5552),
    .C(_09354_),
    .Y(_09427_));
 sg13g2_a22oi_1 _17775_ (.Y(_09428_),
    .B1(_09427_),
    .B2(net5530),
    .A2(_09340_),
    .A1(net5309));
 sg13g2_o21ai_1 _17776_ (.B1(_09355_),
    .Y(_09429_),
    .A1(net5557),
    .A2(net5527));
 sg13g2_nand3_1 _17777_ (.B(_09305_),
    .C(_09429_),
    .A(net5549),
    .Y(_09430_));
 sg13g2_o21ai_1 _17778_ (.B1(_09430_),
    .Y(_09431_),
    .A1(_09295_),
    .A2(_09339_));
 sg13g2_nand2_2 _17779_ (.Y(_09432_),
    .A(_09262_),
    .B(_09318_));
 sg13g2_o21ai_1 _17780_ (.B1(_09432_),
    .Y(_09433_),
    .A1(_09293_),
    .A2(_09346_));
 sg13g2_a22oi_1 _17781_ (.Y(_09434_),
    .B1(_09433_),
    .B2(net5309),
    .A2(_09431_),
    .A1(_09421_));
 sg13g2_o21ai_1 _17782_ (.B1(_09434_),
    .Y(_09435_),
    .A1(_09397_),
    .A2(_09428_));
 sg13g2_nand3_1 _17783_ (.B(net5549),
    .C(_09318_),
    .A(net5275),
    .Y(_09436_));
 sg13g2_nand2_2 _17784_ (.Y(_09437_),
    .A(net5527),
    .B(_09354_));
 sg13g2_a21oi_1 _17785_ (.A1(_09376_),
    .A2(_09437_),
    .Y(_09438_),
    .B1(_09436_));
 sg13g2_nor3_1 _17786_ (.A(_09311_),
    .B(_09312_),
    .C(_09330_),
    .Y(_09439_));
 sg13g2_o21ai_1 _17787_ (.B1(_09439_),
    .Y(_09440_),
    .A1(_09147_),
    .A2(_09167_));
 sg13g2_nand2_2 _17788_ (.Y(_09441_),
    .A(net5554),
    .B(_09321_));
 sg13g2_o21ai_1 _17789_ (.B1(_09440_),
    .Y(_09442_),
    .A1(net5432),
    .A2(_09441_));
 sg13g2_nor4_1 _17790_ (.A(_09419_),
    .B(_09435_),
    .C(_09438_),
    .D(_09442_),
    .Y(_09443_));
 sg13g2_o21ai_1 _17791_ (.B1(_09426_),
    .Y(_00014_),
    .A1(net5541),
    .A2(_09443_));
 sg13g2_nor2_2 _17792_ (.A(net5504),
    .B(_09305_),
    .Y(_09444_));
 sg13g2_nor2_1 _17793_ (.A(_09361_),
    .B(_09444_),
    .Y(_09445_));
 sg13g2_nor2_1 _17794_ (.A(net5264),
    .B(net5480),
    .Y(_09446_));
 sg13g2_a221oi_1 _17795_ (.B2(net5384),
    .C1(_09445_),
    .B1(_09446_),
    .A1(_09105_),
    .Y(_09447_),
    .A2(net5309));
 sg13g2_nor4_2 _17796_ (.A(_09311_),
    .B(_09342_),
    .C(_09397_),
    .Y(_09448_),
    .D(_09427_));
 sg13g2_nor2_1 _17797_ (.A(_09295_),
    .B(_09306_),
    .Y(_09449_));
 sg13g2_a21oi_1 _17798_ (.A1(_09363_),
    .A2(_09449_),
    .Y(_09450_),
    .B1(_09330_));
 sg13g2_o21ai_1 _17799_ (.B1(net5504),
    .Y(_09451_),
    .A1(net5282),
    .A2(net5528));
 sg13g2_nand3_1 _17800_ (.B(_09318_),
    .C(_09451_),
    .A(net5384),
    .Y(_09452_));
 sg13g2_o21ai_1 _17801_ (.B1(_09327_),
    .Y(_09453_),
    .A1(_09376_),
    .A2(_09441_));
 sg13g2_o21ai_1 _17802_ (.B1(_09452_),
    .Y(_09454_),
    .A1(net5542),
    .A2(_09447_));
 sg13g2_nor4_1 _17803_ (.A(_09448_),
    .B(_09450_),
    .C(_09453_),
    .D(_09454_),
    .Y(_09455_));
 sg13g2_o21ai_1 _17804_ (.B1(_09426_),
    .Y(_00015_),
    .A1(net5540),
    .A2(_09455_));
 sg13g2_nand3_1 _17805_ (.B(net5553),
    .C(_09355_),
    .A(net5530),
    .Y(_09456_));
 sg13g2_a21oi_1 _17806_ (.A1(_09291_),
    .A2(_09372_),
    .Y(_09457_),
    .B1(net5272));
 sg13g2_o21ai_1 _17807_ (.B1(_09430_),
    .Y(_09458_),
    .A1(net5565),
    .A2(_09339_));
 sg13g2_nand2b_1 _17808_ (.Y(_09459_),
    .B(_09458_),
    .A_N(_09361_));
 sg13g2_a21oi_1 _17809_ (.A1(net5557),
    .A2(_09358_),
    .Y(_09460_),
    .B1(_09429_));
 sg13g2_nor2_1 _17810_ (.A(net5268),
    .B(_09460_),
    .Y(_09461_));
 sg13g2_a221oi_1 _17811_ (.B2(_09457_),
    .C1(_09461_),
    .B1(_09456_),
    .A1(net5527),
    .Y(_09462_),
    .A2(_09319_));
 sg13g2_a21oi_1 _17812_ (.A1(_09459_),
    .A2(_09462_),
    .Y(_09463_),
    .B1(net5544));
 sg13g2_a21oi_1 _17813_ (.A1(net5565),
    .A2(_09314_),
    .Y(_09464_),
    .B1(_09416_));
 sg13g2_a21oi_1 _17814_ (.A1(_09339_),
    .A2(_09464_),
    .Y(_09465_),
    .B1(_09397_));
 sg13g2_a21oi_1 _17815_ (.A1(net5531),
    .A2(net5550),
    .Y(_09466_),
    .B1(net5282));
 sg13g2_a221oi_1 _17816_ (.B2(_09466_),
    .C1(_09346_),
    .B1(_09338_),
    .A1(net5282),
    .Y(_09467_),
    .A2(net5384));
 sg13g2_nor4_2 _17817_ (.A(_09419_),
    .B(_09463_),
    .C(_09465_),
    .Y(_09468_),
    .D(_09467_));
 sg13g2_o21ai_1 _17818_ (.B1(_09426_),
    .Y(_00016_),
    .A1(net5540),
    .A2(_09468_));
 sg13g2_nor4_1 _17819_ (.A(net6246),
    .B(\atari2600.clk_counter[0] ),
    .C(_08634_),
    .D(_08677_),
    .Y(_09469_));
 sg13g2_a21oi_1 _17820_ (.A1(net6246),
    .A2(_08678_),
    .Y(_09470_),
    .B1(_09469_));
 sg13g2_nand2_1 _17821_ (.Y(_09471_),
    .A(net6571),
    .B(_08710_));
 sg13g2_or2_2 _17822_ (.X(_09472_),
    .B(_09471_),
    .A(_09470_));
 sg13g2_inv_2 _17823_ (.Y(_09473_),
    .A(_09472_));
 sg13g2_a21oi_1 _17824_ (.A1(net7601),
    .A2(_09473_),
    .Y(_09474_),
    .B1(net6531));
 sg13g2_nand2_1 _17825_ (.Y(_09475_),
    .A(net2969),
    .B(net5738));
 sg13g2_xor2_1 _17826_ (.B(net6502),
    .A(\atari2600.tia.diag[58] ),
    .X(_09476_));
 sg13g2_nand2_1 _17827_ (.Y(_09477_),
    .A(_08536_),
    .B(net6504));
 sg13g2_xor2_1 _17828_ (.B(net6504),
    .A(\atari2600.tia.diag[57] ),
    .X(_09478_));
 sg13g2_nor2b_2 _17829_ (.A(net6507),
    .B_N(\atari2600.tia.diag[56] ),
    .Y(_09479_));
 sg13g2_nor2_1 _17830_ (.A(_09478_),
    .B(_09479_),
    .Y(_09480_));
 sg13g2_a21oi_1 _17831_ (.A1(_08536_),
    .A2(net6504),
    .Y(_09481_),
    .B1(_09480_));
 sg13g2_nor2_1 _17832_ (.A(_09476_),
    .B(_09481_),
    .Y(_09482_));
 sg13g2_xor2_1 _17833_ (.B(_09481_),
    .A(_09476_),
    .X(_09483_));
 sg13g2_xor2_1 _17834_ (.B(net6500),
    .A(net6271),
    .X(_09484_));
 sg13g2_a21oi_2 _17835_ (.B1(_09482_),
    .Y(_09485_),
    .A2(net6502),
    .A1(_08535_));
 sg13g2_nor2_1 _17836_ (.A(_09484_),
    .B(_09485_),
    .Y(_09486_));
 sg13g2_xnor2_1 _17837_ (.Y(_09487_),
    .A(_09484_),
    .B(_09485_));
 sg13g2_nor2_1 _17838_ (.A(net6511),
    .B(_09483_),
    .Y(_09488_));
 sg13g2_a21oi_1 _17839_ (.A1(net6511),
    .A2(_09487_),
    .Y(_09489_),
    .B1(_09488_));
 sg13g2_nor2b_1 _17840_ (.A(net6510),
    .B_N(_09489_),
    .Y(_09490_));
 sg13g2_xor2_1 _17841_ (.B(net6496),
    .A(net6270),
    .X(_09491_));
 sg13g2_a21oi_2 _17842_ (.B1(_09486_),
    .Y(_09492_),
    .A2(net6499),
    .A1(_08534_));
 sg13g2_nor2_1 _17843_ (.A(_09491_),
    .B(_09492_),
    .Y(_09493_));
 sg13g2_xor2_1 _17844_ (.B(_09492_),
    .A(_09491_),
    .X(_09494_));
 sg13g2_nor2_1 _17845_ (.A(net6269),
    .B(net6119),
    .Y(_09495_));
 sg13g2_xnor2_1 _17846_ (.Y(_09496_),
    .A(net6269),
    .B(net6492));
 sg13g2_a21oi_2 _17847_ (.B1(_09493_),
    .Y(_09497_),
    .A2(net6496),
    .A1(_08533_));
 sg13g2_inv_1 _17848_ (.Y(_09498_),
    .A(_09497_));
 sg13g2_xnor2_1 _17849_ (.Y(_09499_),
    .A(_09496_),
    .B(_09497_));
 sg13g2_mux2_1 _17850_ (.A0(_09494_),
    .A1(_09499_),
    .S(net6512),
    .X(_09500_));
 sg13g2_a21oi_1 _17851_ (.A1(net6510),
    .A2(_09500_),
    .Y(_09501_),
    .B1(_09490_));
 sg13g2_xnor2_1 _17852_ (.Y(_09502_),
    .A(_00148_),
    .B(_09501_));
 sg13g2_xnor2_1 _17853_ (.Y(_09503_),
    .A(_09478_),
    .B(_09479_));
 sg13g2_nor2_1 _17854_ (.A(net6512),
    .B(_09487_),
    .Y(_09504_));
 sg13g2_a21oi_1 _17855_ (.A1(net6512),
    .A2(_09494_),
    .Y(_09505_),
    .B1(_09504_));
 sg13g2_or2_1 _17856_ (.X(_09506_),
    .B(_09503_),
    .A(net6511));
 sg13g2_a21oi_1 _17857_ (.A1(net6511),
    .A2(_09483_),
    .Y(_09507_),
    .B1(net6510));
 sg13g2_a22oi_1 _17858_ (.Y(_09508_),
    .B1(_09506_),
    .B2(_09507_),
    .A2(_09505_),
    .A1(net6510));
 sg13g2_xnor2_1 _17859_ (.Y(_09509_),
    .A(_00148_),
    .B(_09508_));
 sg13g2_nor2_1 _17860_ (.A(\atari2600.tia.diag[56] ),
    .B(_08629_),
    .Y(_09510_));
 sg13g2_or2_1 _17861_ (.X(_09511_),
    .B(_09510_),
    .A(_09479_));
 sg13g2_or2_1 _17862_ (.X(_09512_),
    .B(_09511_),
    .A(net6511));
 sg13g2_a21oi_1 _17863_ (.A1(net6511),
    .A2(_09503_),
    .Y(_09513_),
    .B1(net6510));
 sg13g2_a22oi_1 _17864_ (.Y(_09514_),
    .B1(_09512_),
    .B2(_09513_),
    .A2(_09489_),
    .A1(net6510));
 sg13g2_xnor2_1 _17865_ (.Y(_09515_),
    .A(_00148_),
    .B(_09514_));
 sg13g2_mux4_1 _17866_ (.S0(_09509_),
    .A0(\atari2600.tia.diag[98] ),
    .A1(\atari2600.tia.diag[96] ),
    .A2(\atari2600.tia.old_grp1[2] ),
    .A3(\atari2600.tia.old_grp1[0] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09516_));
 sg13g2_mux4_1 _17867_ (.S0(_09509_),
    .A0(\atari2600.tia.diag[99] ),
    .A1(\atari2600.tia.diag[97] ),
    .A2(\atari2600.tia.old_grp1[3] ),
    .A3(\atari2600.tia.old_grp1[1] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09517_));
 sg13g2_mux2_1 _17868_ (.A0(_09516_),
    .A1(_09517_),
    .S(_09515_),
    .X(_09518_));
 sg13g2_nor2_1 _17869_ (.A(_09502_),
    .B(_09518_),
    .Y(_09519_));
 sg13g2_mux4_1 _17870_ (.S0(_09509_),
    .A0(\atari2600.tia.diag[102] ),
    .A1(\atari2600.tia.diag[100] ),
    .A2(\atari2600.tia.old_grp1[6] ),
    .A3(\atari2600.tia.old_grp1[4] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09520_));
 sg13g2_nor2_1 _17871_ (.A(_09515_),
    .B(_09520_),
    .Y(_09521_));
 sg13g2_nand2b_1 _17872_ (.Y(_09522_),
    .B(\atari2600.tia.vdelp1 ),
    .A_N(\atari2600.tia.old_grp1[7] ));
 sg13g2_o21ai_1 _17873_ (.B1(_09522_),
    .Y(_09523_),
    .A1(\atari2600.tia.diag[103] ),
    .A2(\atari2600.tia.vdelp1 ));
 sg13g2_mux2_1 _17874_ (.A0(\atari2600.tia.diag[101] ),
    .A1(\atari2600.tia.old_grp1[5] ),
    .S(\atari2600.tia.vdelp1 ),
    .X(_09524_));
 sg13g2_o21ai_1 _17875_ (.B1(_09515_),
    .Y(_09525_),
    .A1(_09509_),
    .A2(_09523_));
 sg13g2_a21oi_1 _17876_ (.A1(_09509_),
    .A2(_09524_),
    .Y(_09526_),
    .B1(_09525_));
 sg13g2_o21ai_1 _17877_ (.B1(_09502_),
    .Y(_09527_),
    .A1(_09521_),
    .A2(_09526_));
 sg13g2_nand2b_1 _17878_ (.Y(_09528_),
    .B(net6487),
    .A_N(\atari2600.tia.p1_spacing[5] ));
 sg13g2_xor2_1 _17879_ (.B(net6487),
    .A(\atari2600.tia.p1_spacing[5] ),
    .X(_09529_));
 sg13g2_nor2b_1 _17880_ (.A(net6492),
    .B_N(\atari2600.tia.p1_spacing[4] ),
    .Y(_09530_));
 sg13g2_o21ai_1 _17881_ (.B1(_09528_),
    .Y(_09531_),
    .A1(_09529_),
    .A2(_09530_));
 sg13g2_xor2_1 _17882_ (.B(net6483),
    .A(\atari2600.tia.p1_spacing[6] ),
    .X(_09532_));
 sg13g2_xnor2_1 _17883_ (.Y(_09533_),
    .A(_09531_),
    .B(_09532_));
 sg13g2_xnor2_1 _17884_ (.Y(_09534_),
    .A(_09529_),
    .B(_09530_));
 sg13g2_xnor2_1 _17885_ (.Y(_09535_),
    .A(\atari2600.tia.p1_spacing[4] ),
    .B(net6492));
 sg13g2_nand2b_1 _17886_ (.Y(_09536_),
    .B(_00146_),
    .A_N(_09535_));
 sg13g2_xnor2_1 _17887_ (.Y(_09537_),
    .A(net6269),
    .B(_09535_));
 sg13g2_o21ai_1 _17888_ (.B1(_09536_),
    .Y(_09538_),
    .A1(_09497_),
    .A2(_09537_));
 sg13g2_xnor2_1 _17889_ (.Y(_09539_),
    .A(_00144_),
    .B(_09534_));
 sg13g2_nand2_1 _17890_ (.Y(_09540_),
    .A(_09538_),
    .B(_09539_));
 sg13g2_o21ai_1 _17891_ (.B1(_09540_),
    .Y(_09541_),
    .A1(\atari2600.tia.diag[62] ),
    .A2(_09534_));
 sg13g2_xnor2_1 _17892_ (.Y(_09542_),
    .A(\atari2600.tia.diag[63] ),
    .B(_09533_));
 sg13g2_a22oi_1 _17893_ (.Y(_09543_),
    .B1(_09541_),
    .B2(_09542_),
    .A2(_09533_),
    .A1(_00147_));
 sg13g2_inv_1 _17894_ (.Y(_09544_),
    .A(_09543_));
 sg13g2_nand2_1 _17895_ (.Y(_09545_),
    .A(net6269),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_xnor2_1 _17896_ (.Y(_09546_),
    .A(net6269),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_nand2_1 _17897_ (.Y(_09547_),
    .A(net6271),
    .B(\atari2600.tia.p1_w[3] ));
 sg13g2_xor2_1 _17898_ (.B(\atari2600.tia.p1_w[4] ),
    .A(net6270),
    .X(_09548_));
 sg13g2_nand2b_1 _17899_ (.Y(_09549_),
    .B(_09548_),
    .A_N(_09547_));
 sg13g2_o21ai_1 _17900_ (.B1(_09549_),
    .Y(_09550_),
    .A1(_08533_),
    .A2(_08562_));
 sg13g2_inv_1 _17901_ (.Y(_09551_),
    .A(_09550_));
 sg13g2_o21ai_1 _17902_ (.B1(_09545_),
    .Y(_09552_),
    .A1(_09546_),
    .A2(_09551_));
 sg13g2_xnor2_1 _17903_ (.Y(_09553_),
    .A(_08531_),
    .B(_09552_));
 sg13g2_nor2_1 _17904_ (.A(_09534_),
    .B(_09553_),
    .Y(_09554_));
 sg13g2_xnor2_1 _17905_ (.Y(_09555_),
    .A(_09546_),
    .B(_09550_));
 sg13g2_xnor2_1 _17906_ (.Y(_09556_),
    .A(_09547_),
    .B(_09548_));
 sg13g2_nor2_1 _17907_ (.A(net6494),
    .B(_09556_),
    .Y(_09557_));
 sg13g2_xor2_1 _17908_ (.B(\atari2600.tia.p1_w[3] ),
    .A(net6271),
    .X(_09558_));
 sg13g2_nor2_1 _17909_ (.A(_00141_),
    .B(_09558_),
    .Y(_09559_));
 sg13g2_xnor2_1 _17910_ (.Y(_09560_),
    .A(net6497),
    .B(_09558_));
 sg13g2_nor2_1 _17911_ (.A(_09476_),
    .B(_09560_),
    .Y(_09561_));
 sg13g2_o21ai_1 _17912_ (.B1(_09510_),
    .Y(_09562_),
    .A1(_08536_),
    .A2(net6504));
 sg13g2_nand3_1 _17913_ (.B(_09561_),
    .C(_09562_),
    .A(_09477_),
    .Y(_09563_));
 sg13g2_nor3_1 _17914_ (.A(_08535_),
    .B(net6502),
    .C(_09559_),
    .Y(_09564_));
 sg13g2_nand2_1 _17915_ (.Y(_09565_),
    .A(net6494),
    .B(_09556_));
 sg13g2_a221oi_1 _17916_ (.B2(net6497),
    .C1(_09564_),
    .B1(_09558_),
    .A1(net6494),
    .Y(_09566_),
    .A2(_09556_));
 sg13g2_a21oi_1 _17917_ (.A1(_09563_),
    .A2(_09566_),
    .Y(_09567_),
    .B1(_09557_));
 sg13g2_nor2_1 _17918_ (.A(_09478_),
    .B(_09511_),
    .Y(_09568_));
 sg13g2_nand3_1 _17919_ (.B(_09565_),
    .C(_09568_),
    .A(_09561_),
    .Y(_09569_));
 sg13g2_nor2_1 _17920_ (.A(_09535_),
    .B(_09555_),
    .Y(_09570_));
 sg13g2_a22oi_1 _17921_ (.Y(_09571_),
    .B1(_09567_),
    .B2(_09569_),
    .A2(_09555_),
    .A1(_09535_));
 sg13g2_nor3_1 _17922_ (.A(_09554_),
    .B(_09570_),
    .C(_09571_),
    .Y(_09572_));
 sg13g2_or3_1 _17923_ (.A(_08531_),
    .B(_09546_),
    .C(_09551_),
    .X(_09573_));
 sg13g2_o21ai_1 _17924_ (.B1(_09573_),
    .Y(_09574_),
    .A1(_00144_),
    .A2(_09545_));
 sg13g2_xnor2_1 _17925_ (.Y(_09575_),
    .A(\atari2600.tia.diag[63] ),
    .B(_09574_));
 sg13g2_nand2_1 _17926_ (.Y(_09576_),
    .A(_09534_),
    .B(_09553_));
 sg13g2_o21ai_1 _17927_ (.B1(_09576_),
    .Y(_09577_),
    .A1(_09533_),
    .A2(_09575_));
 sg13g2_o21ai_1 _17928_ (.B1(\atari2600.tia.p1_copies[1] ),
    .Y(_09578_),
    .A1(_09572_),
    .A2(_09577_));
 sg13g2_a21oi_1 _17929_ (.A1(_09533_),
    .A2(_09575_),
    .Y(_09579_),
    .B1(_09578_));
 sg13g2_xor2_1 _17930_ (.B(net6487),
    .A(\atari2600.tia.diag[62] ),
    .X(_09580_));
 sg13g2_a21oi_1 _17931_ (.A1(_09496_),
    .A2(_09498_),
    .Y(_09581_),
    .B1(_09495_));
 sg13g2_nor2_1 _17932_ (.A(_09580_),
    .B(_09581_),
    .Y(_09582_));
 sg13g2_a21oi_2 _17933_ (.B1(_09582_),
    .Y(_09583_),
    .A2(net6486),
    .A1(_08531_));
 sg13g2_o21ai_1 _17934_ (.B1(_09583_),
    .Y(_09584_),
    .A1(\atari2600.tia.diag[63] ),
    .A2(_08633_));
 sg13g2_xnor2_1 _17935_ (.Y(_09585_),
    .A(_08661_),
    .B(_09555_));
 sg13g2_a22oi_1 _17936_ (.Y(_09586_),
    .B1(_09567_),
    .B2(_09585_),
    .A2(_09555_),
    .A1(net6119));
 sg13g2_xnor2_1 _17937_ (.Y(_09587_),
    .A(net6485),
    .B(_09553_));
 sg13g2_nand2_1 _17938_ (.Y(_09588_),
    .A(net6118),
    .B(_09553_));
 sg13g2_o21ai_1 _17939_ (.B1(_09588_),
    .Y(_09589_),
    .A1(_09586_),
    .A2(_09587_));
 sg13g2_nor2_1 _17940_ (.A(_09557_),
    .B(_09569_),
    .Y(_09590_));
 sg13g2_nand2_1 _17941_ (.Y(_09591_),
    .A(_09585_),
    .B(_09590_));
 sg13g2_o21ai_1 _17942_ (.B1(_09589_),
    .Y(_09592_),
    .A1(_09587_),
    .A2(_09591_));
 sg13g2_o21ai_1 _17943_ (.B1(_09592_),
    .Y(_09593_),
    .A1(net6483),
    .A2(_09575_));
 sg13g2_nor2b_1 _17944_ (.A(net6483),
    .B_N(\atari2600.tia.diag[63] ),
    .Y(_09594_));
 sg13g2_a21oi_1 _17945_ (.A1(net6483),
    .A2(_09575_),
    .Y(_09595_),
    .B1(_09594_));
 sg13g2_nand3_1 _17946_ (.B(_09593_),
    .C(_09595_),
    .A(_09584_),
    .Y(_09596_));
 sg13g2_nand2b_1 _17947_ (.Y(_09597_),
    .B(net6487),
    .A_N(\atari2600.tia.p1_spacing[6] ));
 sg13g2_nor2_1 _17948_ (.A(\atari2600.tia.p1_spacing[5] ),
    .B(net6119),
    .Y(_09598_));
 sg13g2_nand2_1 _17949_ (.Y(_09599_),
    .A(\atari2600.tia.p1_spacing[4] ),
    .B(_08630_));
 sg13g2_xnor2_1 _17950_ (.Y(_09600_),
    .A(\atari2600.tia.p1_spacing[5] ),
    .B(net6492));
 sg13g2_a21oi_1 _17951_ (.A1(_09599_),
    .A2(_09600_),
    .Y(_09601_),
    .B1(_09598_));
 sg13g2_xor2_1 _17952_ (.B(net6487),
    .A(\atari2600.tia.p1_spacing[6] ),
    .X(_09602_));
 sg13g2_o21ai_1 _17953_ (.B1(_09597_),
    .Y(_09603_),
    .A1(_09601_),
    .A2(_09602_));
 sg13g2_xor2_1 _17954_ (.B(_09603_),
    .A(net6480),
    .X(_09604_));
 sg13g2_xnor2_1 _17955_ (.Y(_09605_),
    .A(_09601_),
    .B(_09602_));
 sg13g2_xnor2_1 _17956_ (.Y(_09606_),
    .A(_09599_),
    .B(_09600_));
 sg13g2_xnor2_1 _17957_ (.Y(_09607_),
    .A(\atari2600.tia.p1_spacing[4] ),
    .B(net6495));
 sg13g2_nor2_1 _17958_ (.A(\atari2600.tia.diag[60] ),
    .B(_09607_),
    .Y(_09608_));
 sg13g2_a21oi_1 _17959_ (.A1(\atari2600.tia.diag[60] ),
    .A2(_09607_),
    .Y(_09609_),
    .B1(_09492_));
 sg13g2_xnor2_1 _17960_ (.Y(_09610_),
    .A(_00146_),
    .B(_09606_));
 sg13g2_o21ai_1 _17961_ (.B1(_09610_),
    .Y(_09611_),
    .A1(_09608_),
    .A2(_09609_));
 sg13g2_o21ai_1 _17962_ (.B1(_09611_),
    .Y(_09612_),
    .A1(net6269),
    .A2(_09606_));
 sg13g2_xnor2_1 _17963_ (.Y(_09613_),
    .A(_00144_),
    .B(_09605_));
 sg13g2_nand2_1 _17964_ (.Y(_09614_),
    .A(_09612_),
    .B(_09613_));
 sg13g2_o21ai_1 _17965_ (.B1(_09614_),
    .Y(_09615_),
    .A1(\atari2600.tia.diag[62] ),
    .A2(_09605_));
 sg13g2_xnor2_1 _17966_ (.Y(_09616_),
    .A(\atari2600.tia.diag[63] ),
    .B(_09604_));
 sg13g2_a22oi_1 _17967_ (.Y(_09617_),
    .B1(_09615_),
    .B2(_09616_),
    .A2(_09604_),
    .A1(_00147_));
 sg13g2_nor2_1 _17968_ (.A(_09553_),
    .B(_09605_),
    .Y(_09618_));
 sg13g2_nand2b_1 _17969_ (.Y(_09619_),
    .B(net6499),
    .A_N(_09558_));
 sg13g2_o21ai_1 _17970_ (.B1(_09619_),
    .Y(_09620_),
    .A1(_09485_),
    .A2(_09560_));
 sg13g2_nor2_1 _17971_ (.A(_09556_),
    .B(_09607_),
    .Y(_09621_));
 sg13g2_nor2_1 _17972_ (.A(_09555_),
    .B(_09606_),
    .Y(_09622_));
 sg13g2_a22oi_1 _17973_ (.Y(_09623_),
    .B1(_09607_),
    .B2(_09556_),
    .A2(_09606_),
    .A1(_09555_));
 sg13g2_o21ai_1 _17974_ (.B1(_09623_),
    .Y(_09624_),
    .A1(_09620_),
    .A2(_09621_));
 sg13g2_nor2_1 _17975_ (.A(_09618_),
    .B(_09622_),
    .Y(_09625_));
 sg13g2_nor2_1 _17976_ (.A(_09575_),
    .B(_09604_),
    .Y(_09626_));
 sg13g2_a221oi_1 _17977_ (.B2(_09625_),
    .C1(_09626_),
    .B1(_09624_),
    .A1(_09553_),
    .Y(_09627_),
    .A2(_09605_));
 sg13g2_nand2_1 _17978_ (.Y(_09628_),
    .A(_09575_),
    .B(_09604_));
 sg13g2_o21ai_1 _17979_ (.B1(_09628_),
    .Y(_09629_),
    .A1(\atari2600.tia.p1_copies[2] ),
    .A2(\atari2600.tia.p1_copies[1] ));
 sg13g2_nor3_1 _17980_ (.A(_09617_),
    .B(_09627_),
    .C(_09629_),
    .Y(_09630_));
 sg13g2_a21oi_1 _17981_ (.A1(_09544_),
    .A2(_09579_),
    .Y(_09631_),
    .B1(_09630_));
 sg13g2_xor2_1 _17982_ (.B(net6483),
    .A(\atari2600.tia.diag[63] ),
    .X(_09632_));
 sg13g2_o21ai_1 _17983_ (.B1(net6511),
    .Y(_09633_),
    .A1(_09583_),
    .A2(_09632_));
 sg13g2_a21o_1 _17984_ (.A2(_09632_),
    .A1(_09583_),
    .B1(_09633_),
    .X(_09634_));
 sg13g2_xnor2_1 _17985_ (.Y(_09635_),
    .A(_09580_),
    .B(_09581_));
 sg13g2_nand2b_1 _17986_ (.Y(_09636_),
    .B(_09499_),
    .A_N(net6512));
 sg13g2_nand4_1 _17987_ (.B(_09634_),
    .C(_09635_),
    .A(\atari2600.tia.p1_scale[1] ),
    .Y(_09637_),
    .D(_09636_));
 sg13g2_nor2b_1 _17988_ (.A(net6510),
    .B_N(_09505_),
    .Y(_09638_));
 sg13g2_nand2b_1 _17989_ (.Y(_09639_),
    .B(_09638_),
    .A_N(_09500_));
 sg13g2_a221oi_1 _17990_ (.B2(_09639_),
    .C1(_09519_),
    .B1(_09637_),
    .A1(_09596_),
    .Y(_09640_),
    .A2(_09631_));
 sg13g2_nand2_1 _17991_ (.Y(_09641_),
    .A(_09527_),
    .B(_09640_));
 sg13g2_nor2_1 _17992_ (.A(\atari2600.tia.vid_ypos[3] ),
    .B(_08703_),
    .Y(_09642_));
 sg13g2_nor2_1 _17993_ (.A(\atari2600.tia.vid_ypos[5] ),
    .B(\atari2600.tia.vid_ypos[4] ),
    .Y(_09643_));
 sg13g2_nand3_1 _17994_ (.B(_08701_),
    .C(_09643_),
    .A(_00131_),
    .Y(_09644_));
 sg13g2_o21ai_1 _17995_ (.B1(\atari2600.tia.vid_ypos[8] ),
    .Y(_09645_),
    .A1(_09642_),
    .A2(_09644_));
 sg13g2_nor2b_1 _17996_ (.A(_09472_),
    .B_N(_09645_),
    .Y(_09646_));
 sg13g2_nand2_2 _17997_ (.Y(_09647_),
    .A(_09473_),
    .B(_09645_));
 sg13g2_nor2_1 _17998_ (.A(\atari2600.tia.diag[66] ),
    .B(net6123),
    .Y(_09648_));
 sg13g2_nand2_1 _17999_ (.Y(_09649_),
    .A(\atari2600.tia.diag[66] ),
    .B(net6123));
 sg13g2_nand2b_1 _18000_ (.Y(_09650_),
    .B(_09649_),
    .A_N(_09648_));
 sg13g2_nor2_1 _18001_ (.A(\atari2600.tia.diag[65] ),
    .B(net6122),
    .Y(_09651_));
 sg13g2_xor2_1 _18002_ (.B(net6505),
    .A(\atari2600.tia.diag[65] ),
    .X(_09652_));
 sg13g2_nor2_1 _18003_ (.A(_08540_),
    .B(net6506),
    .Y(_09653_));
 sg13g2_nor2_1 _18004_ (.A(_09652_),
    .B(_09653_),
    .Y(_09654_));
 sg13g2_nor2_1 _18005_ (.A(_09651_),
    .B(_09654_),
    .Y(_09655_));
 sg13g2_inv_1 _18006_ (.Y(_09656_),
    .A(_09655_));
 sg13g2_xor2_1 _18007_ (.B(_09655_),
    .A(_09650_),
    .X(_09657_));
 sg13g2_xnor2_1 _18008_ (.Y(_09658_),
    .A(_09652_),
    .B(_09653_));
 sg13g2_nand2b_1 _18009_ (.Y(_09659_),
    .B(net6498),
    .A_N(net6276));
 sg13g2_nor2b_1 _18010_ (.A(net6498),
    .B_N(net6276),
    .Y(_09660_));
 sg13g2_xnor2_1 _18011_ (.Y(_09661_),
    .A(net6276),
    .B(net6498));
 sg13g2_a21oi_1 _18012_ (.A1(_09649_),
    .A2(_09656_),
    .Y(_09662_),
    .B1(_09648_));
 sg13g2_xnor2_1 _18013_ (.Y(_09663_),
    .A(_09661_),
    .B(_09662_));
 sg13g2_xnor2_1 _18014_ (.Y(_09664_),
    .A(net6275),
    .B(net6495));
 sg13g2_a21oi_1 _18015_ (.A1(_08540_),
    .A2(net6506),
    .Y(_09665_),
    .B1(_09651_));
 sg13g2_a21oi_1 _18016_ (.A1(\atari2600.tia.diag[65] ),
    .A2(net6122),
    .Y(_09666_),
    .B1(_09665_));
 sg13g2_a21oi_1 _18017_ (.A1(_09649_),
    .A2(_09666_),
    .Y(_09667_),
    .B1(_09648_));
 sg13g2_o21ai_1 _18018_ (.B1(_09659_),
    .Y(_09668_),
    .A1(_09660_),
    .A2(_09667_));
 sg13g2_xor2_1 _18019_ (.B(net6506),
    .A(\atari2600.tia.diag[64] ),
    .X(_09669_));
 sg13g2_nor3_1 _18020_ (.A(_09650_),
    .B(_09652_),
    .C(_09669_),
    .Y(_09670_));
 sg13g2_and2_1 _18021_ (.A(_09661_),
    .B(_09670_),
    .X(_09671_));
 sg13g2_nor2_1 _18022_ (.A(_09668_),
    .B(_09671_),
    .Y(_09672_));
 sg13g2_o21ai_1 _18023_ (.B1(_09664_),
    .Y(_09673_),
    .A1(_09668_),
    .A2(_09671_));
 sg13g2_xor2_1 _18024_ (.B(_09672_),
    .A(_09664_),
    .X(_09674_));
 sg13g2_nor2_1 _18025_ (.A(_08561_),
    .B(_09674_),
    .Y(_09675_));
 sg13g2_a21oi_1 _18026_ (.A1(_08561_),
    .A2(_09663_),
    .Y(_09676_),
    .B1(_09675_));
 sg13g2_o21ai_1 _18027_ (.B1(_08560_),
    .Y(_09677_),
    .A1(\atari2600.tia.p0_scale[0] ),
    .A2(_09658_));
 sg13g2_a21oi_1 _18028_ (.A1(\atari2600.tia.p0_scale[0] ),
    .A2(_09657_),
    .Y(_09678_),
    .B1(_09677_));
 sg13g2_a21oi_2 _18029_ (.B1(_09678_),
    .Y(_09679_),
    .A2(_09676_),
    .A1(\atari2600.tia.p0_scale[1] ));
 sg13g2_xor2_1 _18030_ (.B(_09679_),
    .A(_00151_),
    .X(_09680_));
 sg13g2_a21oi_1 _18031_ (.A1(_08561_),
    .A2(_09669_),
    .Y(_09681_),
    .B1(\atari2600.tia.p0_scale[1] ));
 sg13g2_o21ai_1 _18032_ (.B1(_09681_),
    .Y(_09682_),
    .A1(_08561_),
    .A2(_09658_));
 sg13g2_mux2_1 _18033_ (.A0(_09657_),
    .A1(_09663_),
    .S(\atari2600.tia.p0_scale[0] ),
    .X(_09683_));
 sg13g2_o21ai_1 _18034_ (.B1(_09682_),
    .Y(_09684_),
    .A1(_08560_),
    .A2(_09683_));
 sg13g2_xor2_1 _18035_ (.B(_09684_),
    .A(_00151_),
    .X(_09685_));
 sg13g2_mux4_1 _18036_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[104] ),
    .A1(\atari2600.tia.old_grp0[0] ),
    .A2(\atari2600.tia.diag[106] ),
    .A3(\atari2600.tia.old_grp0[2] ),
    .S1(_09680_),
    .X(_09686_));
 sg13g2_nand2_1 _18037_ (.Y(_09687_),
    .A(_09685_),
    .B(_09686_));
 sg13g2_nor2_1 _18038_ (.A(\atari2600.tia.p0_scale[0] ),
    .B(_09674_),
    .Y(_09688_));
 sg13g2_nor2_1 _18039_ (.A(\atari2600.tia.diag[69] ),
    .B(net6119),
    .Y(_09689_));
 sg13g2_xnor2_1 _18040_ (.Y(_09690_),
    .A(\atari2600.tia.diag[69] ),
    .B(net6492));
 sg13g2_o21ai_1 _18041_ (.B1(_09673_),
    .Y(_09691_),
    .A1(net6275),
    .A2(net6121));
 sg13g2_xnor2_1 _18042_ (.Y(_09692_),
    .A(_09690_),
    .B(_09691_));
 sg13g2_inv_1 _18043_ (.Y(_09693_),
    .A(_09692_));
 sg13g2_a21oi_1 _18044_ (.A1(\atari2600.tia.p0_scale[0] ),
    .A2(_09693_),
    .Y(_09694_),
    .B1(_09688_));
 sg13g2_nor2_1 _18045_ (.A(\atari2600.tia.p0_scale[1] ),
    .B(_09683_),
    .Y(_09695_));
 sg13g2_a21oi_2 _18046_ (.B1(_09695_),
    .Y(_09696_),
    .A2(_09694_),
    .A1(\atari2600.tia.p0_scale[1] ));
 sg13g2_xnor2_1 _18047_ (.Y(_09697_),
    .A(_00151_),
    .B(_09696_));
 sg13g2_mux4_1 _18048_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[105] ),
    .A1(\atari2600.tia.old_grp0[1] ),
    .A2(\atari2600.tia.diag[107] ),
    .A3(\atari2600.tia.old_grp0[3] ),
    .S1(_09680_),
    .X(_09698_));
 sg13g2_nand2b_1 _18049_ (.Y(_09699_),
    .B(_09698_),
    .A_N(_09685_));
 sg13g2_and2_1 _18050_ (.A(_09697_),
    .B(_09699_),
    .X(_09700_));
 sg13g2_mux4_1 _18051_ (.S0(_09685_),
    .A0(\atari2600.tia.diag[111] ),
    .A1(\atari2600.tia.diag[110] ),
    .A2(\atari2600.tia.old_grp0[7] ),
    .A3(\atari2600.tia.old_grp0[6] ),
    .S1(\atari2600.tia.vdelp0 ),
    .X(_09701_));
 sg13g2_mux4_1 _18052_ (.S0(_09685_),
    .A0(\atari2600.tia.diag[109] ),
    .A1(\atari2600.tia.diag[108] ),
    .A2(\atari2600.tia.old_grp0[5] ),
    .A3(\atari2600.tia.old_grp0[4] ),
    .S1(\atari2600.tia.vdelp0 ),
    .X(_09702_));
 sg13g2_mux2_1 _18053_ (.A0(_09702_),
    .A1(_09701_),
    .S(_09680_),
    .X(_09703_));
 sg13g2_xor2_1 _18054_ (.B(net6483),
    .A(net6272),
    .X(_09704_));
 sg13g2_nand2_1 _18055_ (.Y(_09705_),
    .A(_08537_),
    .B(net6486));
 sg13g2_xnor2_1 _18056_ (.Y(_09706_),
    .A(\atari2600.tia.diag[70] ),
    .B(net6486));
 sg13g2_a21oi_1 _18057_ (.A1(_09690_),
    .A2(_09691_),
    .Y(_09707_),
    .B1(_09689_));
 sg13g2_nand2b_1 _18058_ (.Y(_09708_),
    .B(_09706_),
    .A_N(_09707_));
 sg13g2_a21o_1 _18059_ (.A2(_09708_),
    .A1(_09705_),
    .B1(_09704_),
    .X(_09709_));
 sg13g2_o21ai_1 _18060_ (.B1(_09709_),
    .Y(_09710_),
    .A1(net6272),
    .A2(_08633_));
 sg13g2_nand2_1 _18061_ (.Y(_09711_),
    .A(\atari2600.tia.diag[69] ),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_xor2_1 _18062_ (.B(\atari2600.tia.p0_w[5] ),
    .A(net6273),
    .X(_09712_));
 sg13g2_xor2_1 _18063_ (.B(\atari2600.tia.p0_w[4] ),
    .A(net6275),
    .X(_09713_));
 sg13g2_nand3_1 _18064_ (.B(\atari2600.tia.p0_w[3] ),
    .C(_09713_),
    .A(\atari2600.tia.diag[67] ),
    .Y(_09714_));
 sg13g2_o21ai_1 _18065_ (.B1(_09714_),
    .Y(_09715_),
    .A1(_08539_),
    .A2(_08559_));
 sg13g2_nand2_1 _18066_ (.Y(_09716_),
    .A(_09712_),
    .B(_09715_));
 sg13g2_nand3_1 _18067_ (.B(_09712_),
    .C(_09715_),
    .A(\atari2600.tia.diag[70] ),
    .Y(_09717_));
 sg13g2_o21ai_1 _18068_ (.B1(_09717_),
    .Y(_09718_),
    .A1(_00149_),
    .A2(_09711_));
 sg13g2_xor2_1 _18069_ (.B(_09718_),
    .A(net6272),
    .X(_09719_));
 sg13g2_nor2_1 _18070_ (.A(net6480),
    .B(_09719_),
    .Y(_09720_));
 sg13g2_nand2_1 _18071_ (.Y(_09721_),
    .A(_09711_),
    .B(_09716_));
 sg13g2_xnor2_1 _18072_ (.Y(_09722_),
    .A(_08537_),
    .B(_09721_));
 sg13g2_xor2_1 _18073_ (.B(_09715_),
    .A(_09712_),
    .X(_09723_));
 sg13g2_nor2_1 _18074_ (.A(net6119),
    .B(_09723_),
    .Y(_09724_));
 sg13g2_a21o_1 _18075_ (.A2(\atari2600.tia.p0_w[3] ),
    .A1(\atari2600.tia.diag[67] ),
    .B1(_09713_),
    .X(_09725_));
 sg13g2_and2_2 _18076_ (.A(_09714_),
    .B(_09725_),
    .X(_09726_));
 sg13g2_nor2_1 _18077_ (.A(net6494),
    .B(_09726_),
    .Y(_09727_));
 sg13g2_xor2_1 _18078_ (.B(\atari2600.tia.p0_w[3] ),
    .A(net6276),
    .X(_09728_));
 sg13g2_nor2_1 _18079_ (.A(net6497),
    .B(_09728_),
    .Y(_09729_));
 sg13g2_a21oi_1 _18080_ (.A1(net6497),
    .A2(_09728_),
    .Y(_09730_),
    .B1(_09662_));
 sg13g2_nor2_1 _18081_ (.A(_09729_),
    .B(_09730_),
    .Y(_09731_));
 sg13g2_nor3_1 _18082_ (.A(_09727_),
    .B(_09729_),
    .C(_09730_),
    .Y(_09732_));
 sg13g2_and2_1 _18083_ (.A(net6494),
    .B(_09726_),
    .X(_09733_));
 sg13g2_xnor2_1 _18084_ (.Y(_09734_),
    .A(_00142_),
    .B(_09723_));
 sg13g2_nor3_1 _18085_ (.A(_09732_),
    .B(_09733_),
    .C(_09734_),
    .Y(_09735_));
 sg13g2_xor2_1 _18086_ (.B(_09722_),
    .A(net6485),
    .X(_09736_));
 sg13g2_o21ai_1 _18087_ (.B1(_09736_),
    .Y(_09737_),
    .A1(_09724_),
    .A2(_09735_));
 sg13g2_o21ai_1 _18088_ (.B1(_09737_),
    .Y(_09738_),
    .A1(net6118),
    .A2(_09722_));
 sg13g2_xnor2_1 _18089_ (.Y(_09739_),
    .A(_09704_),
    .B(_09718_));
 sg13g2_a21oi_1 _18090_ (.A1(_09738_),
    .A2(_09739_),
    .Y(_09740_),
    .B1(_09720_));
 sg13g2_nand2_1 _18091_ (.Y(_09741_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net6119));
 sg13g2_nor2_1 _18092_ (.A(\atari2600.tia.p0_spacing[5] ),
    .B(net6118),
    .Y(_09742_));
 sg13g2_xnor2_1 _18093_ (.Y(_09743_),
    .A(\atari2600.tia.p0_spacing[5] ),
    .B(net6486));
 sg13g2_xnor2_1 _18094_ (.Y(_09744_),
    .A(_09741_),
    .B(_09743_));
 sg13g2_xnor2_1 _18095_ (.Y(_09745_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net6492));
 sg13g2_o21ai_1 _18096_ (.B1(_09668_),
    .Y(_09746_),
    .A1(_08539_),
    .A2(net6495));
 sg13g2_xnor2_1 _18097_ (.Y(_09747_),
    .A(net6273),
    .B(_09745_));
 sg13g2_inv_1 _18098_ (.Y(_09748_),
    .A(_09747_));
 sg13g2_a21oi_1 _18099_ (.A1(_08539_),
    .A2(net6495),
    .Y(_09749_),
    .B1(_09747_));
 sg13g2_a22oi_1 _18100_ (.Y(_09750_),
    .B1(_09746_),
    .B2(_09749_),
    .A2(_09745_),
    .A1(_08662_));
 sg13g2_xnor2_1 _18101_ (.Y(_09751_),
    .A(_00149_),
    .B(_09744_));
 sg13g2_nor2b_1 _18102_ (.A(_09750_),
    .B_N(_09751_),
    .Y(_09752_));
 sg13g2_a21oi_1 _18103_ (.A1(\atari2600.tia.diag[70] ),
    .A2(_09744_),
    .Y(_09753_),
    .B1(_09752_));
 sg13g2_a21oi_1 _18104_ (.A1(_09741_),
    .A2(_09743_),
    .Y(_09754_),
    .B1(_09742_));
 sg13g2_xor2_1 _18105_ (.B(net6483),
    .A(\atari2600.tia.p0_spacing[6] ),
    .X(_09755_));
 sg13g2_xnor2_1 _18106_ (.Y(_09756_),
    .A(_09754_),
    .B(_09755_));
 sg13g2_nand4_1 _18107_ (.B(_09671_),
    .C(_09748_),
    .A(_09664_),
    .Y(_09757_),
    .D(_09751_));
 sg13g2_o21ai_1 _18108_ (.B1(_09757_),
    .Y(_09758_),
    .A1(net6272),
    .A2(_09756_));
 sg13g2_or2_1 _18109_ (.X(_09759_),
    .B(_09758_),
    .A(_09753_));
 sg13g2_o21ai_1 _18110_ (.B1(\atari2600.tia.p0_copies[1] ),
    .Y(_09760_),
    .A1(_09719_),
    .A2(_09756_));
 sg13g2_xor2_1 _18111_ (.B(_09728_),
    .A(net6497),
    .X(_09761_));
 sg13g2_a22oi_1 _18112_ (.Y(_09762_),
    .B1(_09761_),
    .B2(_09667_),
    .A2(_09728_),
    .A1(_08626_));
 sg13g2_a21oi_1 _18113_ (.A1(_09670_),
    .A2(_09761_),
    .Y(_09763_),
    .B1(_09727_));
 sg13g2_nor2b_1 _18114_ (.A(_09762_),
    .B_N(_09763_),
    .Y(_09764_));
 sg13g2_a221oi_1 _18115_ (.B2(_09723_),
    .C1(_09764_),
    .B1(_09745_),
    .A1(net6494),
    .Y(_09765_),
    .A2(_09726_));
 sg13g2_nor2_1 _18116_ (.A(_09723_),
    .B(_09745_),
    .Y(_09766_));
 sg13g2_nor2_1 _18117_ (.A(_09765_),
    .B(_09766_),
    .Y(_09767_));
 sg13g2_o21ai_1 _18118_ (.B1(_09767_),
    .Y(_09768_),
    .A1(_09722_),
    .A2(_09744_));
 sg13g2_a22oi_1 _18119_ (.Y(_09769_),
    .B1(_09756_),
    .B2(_09719_),
    .A2(_09744_),
    .A1(_09722_));
 sg13g2_a221oi_1 _18120_ (.B2(_09769_),
    .C1(_09760_),
    .B1(_09768_),
    .A1(net6272),
    .Y(_09770_),
    .A2(_09756_));
 sg13g2_nand2_2 _18121_ (.Y(_09771_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net6121));
 sg13g2_nor2_1 _18122_ (.A(\atari2600.tia.p0_spacing[5] ),
    .B(net6119),
    .Y(_09772_));
 sg13g2_xnor2_1 _18123_ (.Y(_09773_),
    .A(\atari2600.tia.p0_spacing[5] ),
    .B(net6492));
 sg13g2_xor2_1 _18124_ (.B(_09773_),
    .A(_09771_),
    .X(_09774_));
 sg13g2_xnor2_1 _18125_ (.Y(_09775_),
    .A(_09771_),
    .B(_09773_));
 sg13g2_xnor2_1 _18126_ (.Y(_09776_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net6495));
 sg13g2_o21ai_1 _18127_ (.B1(_09731_),
    .Y(_09777_),
    .A1(_09726_),
    .A2(_09776_));
 sg13g2_a22oi_1 _18128_ (.Y(_09778_),
    .B1(_09776_),
    .B2(_09726_),
    .A2(_09775_),
    .A1(_09723_));
 sg13g2_nand2b_1 _18129_ (.Y(_09779_),
    .B(net6486),
    .A_N(\atari2600.tia.p0_spacing[6] ));
 sg13g2_xor2_1 _18130_ (.B(net6486),
    .A(\atari2600.tia.p0_spacing[6] ),
    .X(_09780_));
 sg13g2_a21oi_1 _18131_ (.A1(_09771_),
    .A2(_09773_),
    .Y(_09781_),
    .B1(_09772_));
 sg13g2_xnor2_1 _18132_ (.Y(_09782_),
    .A(_09780_),
    .B(_09781_));
 sg13g2_nand2b_1 _18133_ (.Y(_09783_),
    .B(_09774_),
    .A_N(_09723_));
 sg13g2_o21ai_1 _18134_ (.B1(_09783_),
    .Y(_09784_),
    .A1(_09722_),
    .A2(_09782_));
 sg13g2_a21oi_1 _18135_ (.A1(_09777_),
    .A2(_09778_),
    .Y(_09785_),
    .B1(_09784_));
 sg13g2_o21ai_1 _18136_ (.B1(_09779_),
    .Y(_09786_),
    .A1(_09780_),
    .A2(_09781_));
 sg13g2_xnor2_1 _18137_ (.Y(_09787_),
    .A(net6480),
    .B(_09786_));
 sg13g2_a221oi_1 _18138_ (.B2(_09719_),
    .C1(_09785_),
    .B1(_09787_),
    .A1(_09722_),
    .Y(_09788_),
    .A2(_09782_));
 sg13g2_xnor2_1 _18139_ (.Y(_09789_),
    .A(_00149_),
    .B(_09782_));
 sg13g2_nor2_1 _18140_ (.A(net6274),
    .B(_09776_),
    .Y(_09790_));
 sg13g2_xnor2_1 _18141_ (.Y(_09791_),
    .A(_00150_),
    .B(_09774_));
 sg13g2_nor2_1 _18142_ (.A(_09790_),
    .B(_09791_),
    .Y(_09792_));
 sg13g2_nand2_1 _18143_ (.Y(_09793_),
    .A(net6274),
    .B(_09776_));
 sg13g2_nand2_1 _18144_ (.Y(_09794_),
    .A(_09668_),
    .B(_09793_));
 sg13g2_a22oi_1 _18145_ (.Y(_09795_),
    .B1(_09792_),
    .B2(_09794_),
    .A2(_09775_),
    .A1(net6273));
 sg13g2_inv_1 _18146_ (.Y(_09796_),
    .A(_09795_));
 sg13g2_a22oi_1 _18147_ (.Y(_09797_),
    .B1(_09789_),
    .B2(_09796_),
    .A2(_09782_),
    .A1(\atari2600.tia.diag[70] ));
 sg13g2_nand4_1 _18148_ (.B(_09789_),
    .C(_09792_),
    .A(_09671_),
    .Y(_09798_),
    .D(_09793_));
 sg13g2_o21ai_1 _18149_ (.B1(_09798_),
    .Y(_09799_),
    .A1(net6272),
    .A2(_09787_));
 sg13g2_nor2_1 _18150_ (.A(_09797_),
    .B(_09799_),
    .Y(_09800_));
 sg13g2_nor2_1 _18151_ (.A(\atari2600.tia.p0_copies[2] ),
    .B(\atari2600.tia.p0_copies[1] ),
    .Y(_09801_));
 sg13g2_a21oi_1 _18152_ (.A1(net6272),
    .A2(_09787_),
    .Y(_09802_),
    .B1(_09801_));
 sg13g2_o21ai_1 _18153_ (.B1(_09802_),
    .Y(_09803_),
    .A1(_09719_),
    .A2(_09787_));
 sg13g2_or3_1 _18154_ (.A(_09788_),
    .B(_09800_),
    .C(_09803_),
    .X(_09804_));
 sg13g2_a22oi_1 _18155_ (.Y(_09805_),
    .B1(_09759_),
    .B2(_09770_),
    .A2(_09740_),
    .A1(_09710_));
 sg13g2_nand3_1 _18156_ (.B(_09705_),
    .C(_09708_),
    .A(_09704_),
    .Y(_09806_));
 sg13g2_nand3_1 _18157_ (.B(_09709_),
    .C(_09806_),
    .A(\atari2600.tia.p0_scale[0] ),
    .Y(_09807_));
 sg13g2_nand2b_1 _18158_ (.Y(_09808_),
    .B(_09707_),
    .A_N(_09706_));
 sg13g2_a22oi_1 _18159_ (.Y(_09809_),
    .B1(_09708_),
    .B2(_09808_),
    .A2(_09693_),
    .A1(_08561_));
 sg13g2_nand2_1 _18160_ (.Y(_09810_),
    .A(_09807_),
    .B(_09809_));
 sg13g2_a21oi_1 _18161_ (.A1(_09676_),
    .A2(_09694_),
    .Y(_09811_),
    .B1(\atari2600.tia.p0_scale[1] ));
 sg13g2_a221oi_1 _18162_ (.B2(\atari2600.tia.p0_scale[1] ),
    .C1(_09811_),
    .B1(_09810_),
    .A1(_09804_),
    .Y(_09812_),
    .A2(_09805_));
 sg13g2_o21ai_1 _18163_ (.B1(_09812_),
    .Y(_09813_),
    .A1(_09697_),
    .A2(_09703_));
 sg13g2_a21oi_1 _18164_ (.A1(_09687_),
    .A2(_09700_),
    .Y(_09814_),
    .B1(_09813_));
 sg13g2_nand2_2 _18165_ (.Y(_09815_),
    .A(net5758),
    .B(net5292));
 sg13g2_inv_1 _18166_ (.Y(_09816_),
    .A(_09815_));
 sg13g2_o21ai_1 _18167_ (.B1(net2970),
    .Y(_00029_),
    .A1(net5262),
    .A2(_09815_));
 sg13g2_nand2_1 _18168_ (.Y(_09817_),
    .A(net2998),
    .B(net5737));
 sg13g2_and2_1 _18169_ (.A(\atari2600.tia.diag[51] ),
    .B(\atari2600.tia.m0_w[3] ),
    .X(_09818_));
 sg13g2_nand2_1 _18170_ (.Y(_09819_),
    .A(\atari2600.tia.diag[50] ),
    .B(\atari2600.tia.m0_w[2] ));
 sg13g2_xnor2_1 _18171_ (.Y(_09820_),
    .A(\atari2600.tia.diag[50] ),
    .B(\atari2600.tia.m0_w[2] ));
 sg13g2_nand2_1 _18172_ (.Y(_09821_),
    .A(\atari2600.tia.diag[49] ),
    .B(\atari2600.tia.m0_w[1] ));
 sg13g2_nor2_1 _18173_ (.A(\atari2600.tia.diag[49] ),
    .B(\atari2600.tia.m0_w[1] ),
    .Y(_09822_));
 sg13g2_xor2_1 _18174_ (.B(\atari2600.tia.m0_w[1] ),
    .A(\atari2600.tia.diag[49] ),
    .X(_09823_));
 sg13g2_nand2_1 _18175_ (.Y(_09824_),
    .A(\atari2600.tia.diag[48] ),
    .B(\atari2600.tia.m0_w[0] ));
 sg13g2_o21ai_1 _18176_ (.B1(_09821_),
    .Y(_09825_),
    .A1(_09822_),
    .A2(_09824_));
 sg13g2_inv_1 _18177_ (.Y(_09826_),
    .A(_09825_));
 sg13g2_o21ai_1 _18178_ (.B1(_09819_),
    .Y(_09827_),
    .A1(_09820_),
    .A2(_09826_));
 sg13g2_xor2_1 _18179_ (.B(\atari2600.tia.m0_w[3] ),
    .A(\atari2600.tia.diag[51] ),
    .X(_09828_));
 sg13g2_a21o_1 _18180_ (.A2(_09828_),
    .A1(_09827_),
    .B1(_09818_),
    .X(_09829_));
 sg13g2_and2_1 _18181_ (.A(\atari2600.tia.diag[52] ),
    .B(_09829_),
    .X(_09830_));
 sg13g2_nand3_1 _18182_ (.B(\atari2600.tia.diag[53] ),
    .C(_09830_),
    .A(\atari2600.tia.diag[54] ),
    .Y(_09831_));
 sg13g2_xnor2_1 _18183_ (.Y(_09832_),
    .A(_08528_),
    .B(_09831_));
 sg13g2_a21o_1 _18184_ (.A2(_09830_),
    .A1(net6268),
    .B1(\atari2600.tia.diag[54] ),
    .X(_09833_));
 sg13g2_nand2_1 _18185_ (.Y(_09834_),
    .A(_09831_),
    .B(_09833_));
 sg13g2_xnor2_1 _18186_ (.Y(_09835_),
    .A(net6268),
    .B(_09830_));
 sg13g2_xnor2_1 _18187_ (.Y(_09836_),
    .A(_09823_),
    .B(_09824_));
 sg13g2_xnor2_1 _18188_ (.Y(_09837_),
    .A(\atari2600.tia.diag[48] ),
    .B(\atari2600.tia.m0_w[0] ));
 sg13g2_xnor2_1 _18189_ (.Y(_09838_),
    .A(_00152_),
    .B(_09836_));
 sg13g2_a21oi_1 _18190_ (.A1(net6506),
    .A2(_09837_),
    .Y(_09839_),
    .B1(_09838_));
 sg13g2_a21o_1 _18191_ (.A2(_09836_),
    .A1(net6122),
    .B1(_09839_),
    .X(_09840_));
 sg13g2_xor2_1 _18192_ (.B(_09829_),
    .A(\atari2600.tia.diag[52] ),
    .X(_09841_));
 sg13g2_nor2_1 _18193_ (.A(net6493),
    .B(_09841_),
    .Y(_09842_));
 sg13g2_xnor2_1 _18194_ (.Y(_09843_),
    .A(_09827_),
    .B(_09828_));
 sg13g2_and2_1 _18195_ (.A(net6499),
    .B(_09843_),
    .X(_09844_));
 sg13g2_nor2_1 _18196_ (.A(net6499),
    .B(_09843_),
    .Y(_09845_));
 sg13g2_xnor2_1 _18197_ (.Y(_09846_),
    .A(_09820_),
    .B(_09825_));
 sg13g2_xnor2_1 _18198_ (.Y(_09847_),
    .A(_00140_),
    .B(_09846_));
 sg13g2_nor4_1 _18199_ (.A(_09842_),
    .B(_09844_),
    .C(_09845_),
    .D(_09847_),
    .Y(_09848_));
 sg13g2_a21oi_1 _18200_ (.A1(net6123),
    .A2(_09846_),
    .Y(_09849_),
    .B1(_09845_));
 sg13g2_nor3_1 _18201_ (.A(_09842_),
    .B(_09844_),
    .C(_09849_),
    .Y(_09850_));
 sg13g2_a221oi_1 _18202_ (.B2(_09840_),
    .C1(_09850_),
    .B1(_09848_),
    .A1(net6493),
    .Y(_09851_),
    .A2(_09841_));
 sg13g2_xnor2_1 _18203_ (.Y(_09852_),
    .A(_00142_),
    .B(_09835_));
 sg13g2_nand2b_1 _18204_ (.Y(_09853_),
    .B(_09852_),
    .A_N(_09851_));
 sg13g2_o21ai_1 _18205_ (.B1(_09853_),
    .Y(_09854_),
    .A1(net6490),
    .A2(_09835_));
 sg13g2_xnor2_1 _18206_ (.Y(_09855_),
    .A(net6484),
    .B(_09834_));
 sg13g2_nand2_1 _18207_ (.Y(_09856_),
    .A(_09854_),
    .B(_09855_));
 sg13g2_o21ai_1 _18208_ (.B1(_09856_),
    .Y(_09857_),
    .A1(net6488),
    .A2(_09834_));
 sg13g2_xor2_1 _18209_ (.B(_09837_),
    .A(_00153_),
    .X(_09858_));
 sg13g2_a21oi_1 _18210_ (.A1(net6493),
    .A2(_09841_),
    .Y(_09859_),
    .B1(_09838_));
 sg13g2_nand4_1 _18211_ (.B(_09852_),
    .C(_09855_),
    .A(_09848_),
    .Y(_09860_),
    .D(_09859_));
 sg13g2_o21ai_1 _18212_ (.B1(_09857_),
    .Y(_09861_),
    .A1(_09858_),
    .A2(_09860_));
 sg13g2_o21ai_1 _18213_ (.B1(_09861_),
    .Y(_09862_),
    .A1(net6482),
    .A2(_09832_));
 sg13g2_nand2_1 _18214_ (.Y(_09863_),
    .A(net6268),
    .B(net6120));
 sg13g2_nor2_1 _18215_ (.A(\atari2600.tia.diag[52] ),
    .B(net6121),
    .Y(_09864_));
 sg13g2_nand2b_1 _18216_ (.Y(_09865_),
    .B(net6505),
    .A_N(\atari2600.tia.diag[49] ));
 sg13g2_and3_1 _18217_ (.X(_09866_),
    .A(\atari2600.tia.diag[48] ),
    .B(_08629_),
    .C(_09865_));
 sg13g2_a221oi_1 _18218_ (.B2(\atari2600.tia.diag[49] ),
    .C1(_09866_),
    .B1(net6122),
    .A1(\atari2600.tia.diag[50] ),
    .Y(_09867_),
    .A2(net6123));
 sg13g2_a221oi_1 _18219_ (.B2(_08530_),
    .C1(_09867_),
    .B1(net6502),
    .A1(_08529_),
    .Y(_09868_),
    .A2(net6499));
 sg13g2_a221oi_1 _18220_ (.B2(\atari2600.tia.diag[52] ),
    .C1(_09868_),
    .B1(net6121),
    .A1(\atari2600.tia.diag[51] ),
    .Y(_09869_),
    .A2(_08626_));
 sg13g2_o21ai_1 _18221_ (.B1(_09863_),
    .Y(_09870_),
    .A1(_09864_),
    .A2(_09869_));
 sg13g2_nand2b_1 _18222_ (.Y(_09871_),
    .B(net6488),
    .A_N(\atari2600.tia.diag[54] ));
 sg13g2_o21ai_1 _18223_ (.B1(_09871_),
    .Y(_09872_),
    .A1(net6268),
    .A2(net6120));
 sg13g2_nand2b_1 _18224_ (.Y(_09873_),
    .B(_09870_),
    .A_N(_09872_));
 sg13g2_a22oi_1 _18225_ (.Y(_09874_),
    .B1(_08633_),
    .B2(\atari2600.tia.diag[55] ),
    .A2(_08632_),
    .A1(\atari2600.tia.diag[54] ));
 sg13g2_a22oi_1 _18226_ (.Y(_09875_),
    .B1(_09873_),
    .B2(_09874_),
    .A2(net6482),
    .A1(_08528_));
 sg13g2_a21oi_1 _18227_ (.A1(net6482),
    .A2(_09832_),
    .Y(_09876_),
    .B1(_09875_));
 sg13g2_nand3_1 _18228_ (.B(_09862_),
    .C(_09876_),
    .A(net7588),
    .Y(_09877_));
 sg13g2_nand2_1 _18229_ (.Y(_09878_),
    .A(\atari2600.tia.diag[43] ),
    .B(\atari2600.tia.m1_w[3] ));
 sg13g2_and2_1 _18230_ (.A(\atari2600.tia.diag[42] ),
    .B(\atari2600.tia.m1_w[2] ),
    .X(_09879_));
 sg13g2_xor2_1 _18231_ (.B(\atari2600.tia.m1_w[2] ),
    .A(\atari2600.tia.diag[42] ),
    .X(_09880_));
 sg13g2_nand2_1 _18232_ (.Y(_09881_),
    .A(\atari2600.tia.diag[41] ),
    .B(\atari2600.tia.m1_w[1] ));
 sg13g2_nor2_1 _18233_ (.A(\atari2600.tia.diag[41] ),
    .B(\atari2600.tia.m1_w[1] ),
    .Y(_09882_));
 sg13g2_xor2_1 _18234_ (.B(\atari2600.tia.m1_w[1] ),
    .A(\atari2600.tia.diag[41] ),
    .X(_09883_));
 sg13g2_nand2_1 _18235_ (.Y(_09884_),
    .A(\atari2600.tia.diag[40] ),
    .B(\atari2600.tia.m1_w[0] ));
 sg13g2_o21ai_1 _18236_ (.B1(_09881_),
    .Y(_09885_),
    .A1(_09882_),
    .A2(_09884_));
 sg13g2_a21o_1 _18237_ (.A2(_09885_),
    .A1(_09880_),
    .B1(_09879_),
    .X(_09886_));
 sg13g2_xor2_1 _18238_ (.B(\atari2600.tia.m1_w[3] ),
    .A(\atari2600.tia.diag[43] ),
    .X(_09887_));
 sg13g2_nand2_1 _18239_ (.Y(_09888_),
    .A(_09886_),
    .B(_09887_));
 sg13g2_a21oi_2 _18240_ (.B1(_08525_),
    .Y(_09889_),
    .A2(_09888_),
    .A1(_09878_));
 sg13g2_nand3_1 _18241_ (.B(\atari2600.tia.diag[45] ),
    .C(_09889_),
    .A(\atari2600.tia.diag[46] ),
    .Y(_09890_));
 sg13g2_xnor2_1 _18242_ (.Y(_09891_),
    .A(_08522_),
    .B(_09890_));
 sg13g2_a21o_1 _18243_ (.A2(_09889_),
    .A1(\atari2600.tia.diag[45] ),
    .B1(\atari2600.tia.diag[46] ),
    .X(_09892_));
 sg13g2_nand2_1 _18244_ (.Y(_09893_),
    .A(_09890_),
    .B(_09892_));
 sg13g2_nand3_1 _18245_ (.B(_09890_),
    .C(_09892_),
    .A(net6118),
    .Y(_09894_));
 sg13g2_xnor2_1 _18246_ (.Y(_09895_),
    .A(\atari2600.tia.diag[45] ),
    .B(_09889_));
 sg13g2_nor2_1 _18247_ (.A(net6491),
    .B(_09895_),
    .Y(_09896_));
 sg13g2_nand3_1 _18248_ (.B(_09878_),
    .C(_09888_),
    .A(_08525_),
    .Y(_09897_));
 sg13g2_nor2b_1 _18249_ (.A(_09889_),
    .B_N(_09897_),
    .Y(_09898_));
 sg13g2_and2_1 _18250_ (.A(_00145_),
    .B(_09898_),
    .X(_09899_));
 sg13g2_xnor2_1 _18251_ (.Y(_09900_),
    .A(_09886_),
    .B(_09887_));
 sg13g2_nand2_1 _18252_ (.Y(_09901_),
    .A(net6499),
    .B(_09900_));
 sg13g2_o21ai_1 _18253_ (.B1(_09901_),
    .Y(_09902_),
    .A1(_00145_),
    .A2(_09898_));
 sg13g2_inv_1 _18254_ (.Y(_09903_),
    .A(_09902_));
 sg13g2_nor2_1 _18255_ (.A(net6499),
    .B(_09900_),
    .Y(_09904_));
 sg13g2_xnor2_1 _18256_ (.Y(_09905_),
    .A(_09880_),
    .B(_09885_));
 sg13g2_xnor2_1 _18257_ (.Y(_09906_),
    .A(_09883_),
    .B(_09884_));
 sg13g2_and2_1 _18258_ (.A(net6122),
    .B(_09906_),
    .X(_09907_));
 sg13g2_xnor2_1 _18259_ (.Y(_09908_),
    .A(\atari2600.tia.diag[40] ),
    .B(\atari2600.tia.m1_w[0] ));
 sg13g2_xnor2_1 _18260_ (.Y(_09909_),
    .A(_00152_),
    .B(_09906_));
 sg13g2_a21oi_1 _18261_ (.A1(net6506),
    .A2(_09908_),
    .Y(_09910_),
    .B1(_09909_));
 sg13g2_xnor2_1 _18262_ (.Y(_09911_),
    .A(_00140_),
    .B(_09905_));
 sg13g2_o21ai_1 _18263_ (.B1(_09911_),
    .Y(_09912_),
    .A1(_09907_),
    .A2(_09910_));
 sg13g2_o21ai_1 _18264_ (.B1(_09912_),
    .Y(_09913_),
    .A1(net6502),
    .A2(_09905_));
 sg13g2_o21ai_1 _18265_ (.B1(_09903_),
    .Y(_09914_),
    .A1(_09904_),
    .A2(_09913_));
 sg13g2_nand2b_1 _18266_ (.Y(_09915_),
    .B(_09914_),
    .A_N(_09899_));
 sg13g2_xnor2_1 _18267_ (.Y(_09916_),
    .A(_00142_),
    .B(_09895_));
 sg13g2_a21oi_1 _18268_ (.A1(_09915_),
    .A2(_09916_),
    .Y(_09917_),
    .B1(_09896_));
 sg13g2_xor2_1 _18269_ (.B(_09893_),
    .A(net6484),
    .X(_09918_));
 sg13g2_o21ai_1 _18270_ (.B1(_09894_),
    .Y(_09919_),
    .A1(_09917_),
    .A2(_09918_));
 sg13g2_xor2_1 _18271_ (.B(_09908_),
    .A(_00153_),
    .X(_09920_));
 sg13g2_nor4_1 _18272_ (.A(_09899_),
    .B(_09904_),
    .C(_09909_),
    .D(_09920_),
    .Y(_09921_));
 sg13g2_nand4_1 _18273_ (.B(_09911_),
    .C(_09916_),
    .A(_09903_),
    .Y(_09922_),
    .D(_09921_));
 sg13g2_o21ai_1 _18274_ (.B1(_09919_),
    .Y(_09923_),
    .A1(_09918_),
    .A2(_09922_));
 sg13g2_o21ai_1 _18275_ (.B1(_09923_),
    .Y(_09924_),
    .A1(net6481),
    .A2(_09891_));
 sg13g2_nand2b_1 _18276_ (.Y(_09925_),
    .B(net6505),
    .A_N(\atari2600.tia.diag[41] ));
 sg13g2_and3_1 _18277_ (.X(_09926_),
    .A(\atari2600.tia.diag[40] ),
    .B(_08629_),
    .C(_09925_));
 sg13g2_a221oi_1 _18278_ (.B2(\atari2600.tia.diag[41] ),
    .C1(_09926_),
    .B1(net6122),
    .A1(\atari2600.tia.diag[42] ),
    .Y(_09927_),
    .A2(net6123));
 sg13g2_a221oi_1 _18279_ (.B2(_08527_),
    .C1(_09927_),
    .B1(net6502),
    .A1(_08526_),
    .Y(_09928_),
    .A2(net6498));
 sg13g2_a221oi_1 _18280_ (.B2(\atari2600.tia.diag[44] ),
    .C1(_09928_),
    .B1(_08630_),
    .A1(\atari2600.tia.diag[43] ),
    .Y(_09929_),
    .A2(_08626_));
 sg13g2_a221oi_1 _18281_ (.B2(_08524_),
    .C1(_09929_),
    .B1(net6492),
    .A1(_08525_),
    .Y(_09930_),
    .A2(net6496));
 sg13g2_a221oi_1 _18282_ (.B2(\atari2600.tia.diag[46] ),
    .C1(_09930_),
    .B1(net6118),
    .A1(\atari2600.tia.diag[45] ),
    .Y(_09931_),
    .A2(net6120));
 sg13g2_a221oi_1 _18283_ (.B2(_08522_),
    .C1(_09931_),
    .B1(net6481),
    .A1(_08523_),
    .Y(_09932_),
    .A2(net6489));
 sg13g2_o21ai_1 _18284_ (.B1(\atari2600.tia.enam1 ),
    .Y(_09933_),
    .A1(_08522_),
    .A2(net6481));
 sg13g2_nor2_1 _18285_ (.A(_09932_),
    .B(_09933_),
    .Y(_09934_));
 sg13g2_nand2_1 _18286_ (.Y(_09935_),
    .A(_09924_),
    .B(_09934_));
 sg13g2_a21oi_2 _18287_ (.B1(_09935_),
    .Y(_09936_),
    .A2(_09891_),
    .A1(\atari2600.tia.vid_xpos[7] ));
 sg13g2_nand2_1 _18288_ (.Y(_09937_),
    .A(net5758),
    .B(net5286));
 sg13g2_o21ai_1 _18289_ (.B1(_09817_),
    .Y(_00023_),
    .A1(net5289),
    .A2(_09937_));
 sg13g2_nand2_1 _18290_ (.Y(_09938_),
    .A(net2981),
    .B(net5737));
 sg13g2_nand2_1 _18291_ (.Y(_09939_),
    .A(\atari2600.tia.diag[35] ),
    .B(\atari2600.tia.ball_w[3] ));
 sg13g2_and2_1 _18292_ (.A(\atari2600.tia.diag[34] ),
    .B(\atari2600.tia.ball_w[2] ),
    .X(_09940_));
 sg13g2_or2_1 _18293_ (.X(_09941_),
    .B(\atari2600.tia.ball_w[2] ),
    .A(\atari2600.tia.diag[34] ));
 sg13g2_nand2b_1 _18294_ (.Y(_09942_),
    .B(_09941_),
    .A_N(_09940_));
 sg13g2_nand2_1 _18295_ (.Y(_09943_),
    .A(\atari2600.tia.diag[33] ),
    .B(\atari2600.tia.ball_w[1] ));
 sg13g2_nor2_1 _18296_ (.A(\atari2600.tia.diag[33] ),
    .B(\atari2600.tia.ball_w[1] ),
    .Y(_09944_));
 sg13g2_xor2_1 _18297_ (.B(\atari2600.tia.ball_w[1] ),
    .A(\atari2600.tia.diag[33] ),
    .X(_09945_));
 sg13g2_nand2_1 _18298_ (.Y(_09946_),
    .A(\atari2600.tia.diag[32] ),
    .B(\atari2600.tia.ball_w[0] ));
 sg13g2_o21ai_1 _18299_ (.B1(_09943_),
    .Y(_09947_),
    .A1(_09944_),
    .A2(_09946_));
 sg13g2_a21oi_1 _18300_ (.A1(_09941_),
    .A2(_09947_),
    .Y(_09948_),
    .B1(_09940_));
 sg13g2_xnor2_1 _18301_ (.Y(_09949_),
    .A(\atari2600.tia.diag[35] ),
    .B(\atari2600.tia.ball_w[3] ));
 sg13g2_o21ai_1 _18302_ (.B1(_09939_),
    .Y(_09950_),
    .A1(_09948_),
    .A2(_09949_));
 sg13g2_and2_1 _18303_ (.A(\atari2600.tia.diag[36] ),
    .B(_09950_),
    .X(_09951_));
 sg13g2_nand3_1 _18304_ (.B(\atari2600.tia.diag[37] ),
    .C(_09951_),
    .A(\atari2600.tia.diag[38] ),
    .Y(_09952_));
 sg13g2_xor2_1 _18305_ (.B(_09952_),
    .A(\atari2600.tia.diag[39] ),
    .X(_09953_));
 sg13g2_a21o_1 _18306_ (.A2(_09951_),
    .A1(\atari2600.tia.diag[37] ),
    .B1(\atari2600.tia.diag[38] ),
    .X(_09954_));
 sg13g2_nand2_1 _18307_ (.Y(_09955_),
    .A(_09952_),
    .B(_09954_));
 sg13g2_nor2_1 _18308_ (.A(net6488),
    .B(_09955_),
    .Y(_09956_));
 sg13g2_xnor2_1 _18309_ (.Y(_09957_),
    .A(\atari2600.tia.diag[37] ),
    .B(_09951_));
 sg13g2_xnor2_1 _18310_ (.Y(_09958_),
    .A(_08521_),
    .B(_09950_));
 sg13g2_xnor2_1 _18311_ (.Y(_09959_),
    .A(_09948_),
    .B(_09949_));
 sg13g2_nor2_1 _18312_ (.A(net6493),
    .B(_09958_),
    .Y(_09960_));
 sg13g2_a21oi_1 _18313_ (.A1(net6498),
    .A2(_09959_),
    .Y(_09961_),
    .B1(_09960_));
 sg13g2_nor2_1 _18314_ (.A(net6498),
    .B(_09959_),
    .Y(_09962_));
 sg13g2_xnor2_1 _18315_ (.Y(_09963_),
    .A(_09942_),
    .B(_09947_));
 sg13g2_nand2_1 _18316_ (.Y(_09964_),
    .A(net6123),
    .B(_09963_));
 sg13g2_xnor2_1 _18317_ (.Y(_09965_),
    .A(_09945_),
    .B(_09946_));
 sg13g2_xnor2_1 _18318_ (.Y(_09966_),
    .A(\atari2600.tia.diag[32] ),
    .B(\atari2600.tia.ball_w[0] ));
 sg13g2_nand2_1 _18319_ (.Y(_09967_),
    .A(net6506),
    .B(_09966_));
 sg13g2_xor2_1 _18320_ (.B(_09965_),
    .A(_00152_),
    .X(_09968_));
 sg13g2_a22oi_1 _18321_ (.Y(_09969_),
    .B1(_09967_),
    .B2(_09968_),
    .A2(_09965_),
    .A1(net6122));
 sg13g2_xnor2_1 _18322_ (.Y(_09970_),
    .A(_00140_),
    .B(_09963_));
 sg13g2_o21ai_1 _18323_ (.B1(_09964_),
    .Y(_09971_),
    .A1(_09969_),
    .A2(_09970_));
 sg13g2_nor2_1 _18324_ (.A(_09962_),
    .B(_09970_),
    .Y(_09972_));
 sg13g2_or2_1 _18325_ (.X(_09973_),
    .B(_09971_),
    .A(_09962_));
 sg13g2_a22oi_1 _18326_ (.Y(_09974_),
    .B1(_09961_),
    .B2(_09973_),
    .A2(_09958_),
    .A1(net6494));
 sg13g2_xnor2_1 _18327_ (.Y(_09975_),
    .A(_00142_),
    .B(_09957_));
 sg13g2_nand2b_1 _18328_ (.Y(_09976_),
    .B(_09975_),
    .A_N(_09974_));
 sg13g2_o21ai_1 _18329_ (.B1(_09976_),
    .Y(_09977_),
    .A1(net6491),
    .A2(_09957_));
 sg13g2_xnor2_1 _18330_ (.Y(_09978_),
    .A(net6484),
    .B(_09955_));
 sg13g2_a21oi_1 _18331_ (.A1(_09977_),
    .A2(_09978_),
    .Y(_09979_),
    .B1(_09956_));
 sg13g2_xnor2_1 _18332_ (.Y(_09980_),
    .A(_00153_),
    .B(_09966_));
 sg13g2_nand3_1 _18333_ (.B(_09972_),
    .C(_09980_),
    .A(_09968_),
    .Y(_09981_));
 sg13g2_a21oi_1 _18334_ (.A1(net6493),
    .A2(_09958_),
    .Y(_09982_),
    .B1(_09981_));
 sg13g2_nand4_1 _18335_ (.B(_09975_),
    .C(_09978_),
    .A(_09961_),
    .Y(_09983_),
    .D(_09982_));
 sg13g2_nand2b_1 _18336_ (.Y(_09984_),
    .B(_09983_),
    .A_N(_09979_));
 sg13g2_o21ai_1 _18337_ (.B1(_09984_),
    .Y(_09985_),
    .A1(net6481),
    .A2(_09953_));
 sg13g2_nand2_1 _18338_ (.Y(_09986_),
    .A(net6481),
    .B(_09953_));
 sg13g2_nor2_1 _18339_ (.A(\atari2600.tia.diag[38] ),
    .B(_08632_),
    .Y(_09987_));
 sg13g2_nand2b_1 _18340_ (.Y(_09988_),
    .B(net6505),
    .A_N(\atari2600.tia.diag[33] ));
 sg13g2_nand3_1 _18341_ (.B(_08629_),
    .C(_09988_),
    .A(\atari2600.tia.diag[32] ),
    .Y(_09989_));
 sg13g2_a22oi_1 _18342_ (.Y(_09990_),
    .B1(net6122),
    .B2(\atari2600.tia.diag[33] ),
    .A2(net6123),
    .A1(\atari2600.tia.diag[34] ));
 sg13g2_nand2b_1 _18343_ (.Y(_09991_),
    .B(net6498),
    .A_N(\atari2600.tia.diag[35] ));
 sg13g2_o21ai_1 _18344_ (.B1(_09991_),
    .Y(_09992_),
    .A1(\atari2600.tia.diag[34] ),
    .A2(net6123));
 sg13g2_a21oi_1 _18345_ (.A1(_09989_),
    .A2(_09990_),
    .Y(_09993_),
    .B1(_09992_));
 sg13g2_a221oi_1 _18346_ (.B2(\atari2600.tia.diag[36] ),
    .C1(_09993_),
    .B1(net6121),
    .A1(\atari2600.tia.diag[35] ),
    .Y(_09994_),
    .A2(_08626_));
 sg13g2_a221oi_1 _18347_ (.B2(_08520_),
    .C1(_09994_),
    .B1(net6490),
    .A1(_08521_),
    .Y(_09995_),
    .A2(net6496));
 sg13g2_a21oi_1 _18348_ (.A1(\atari2600.tia.diag[37] ),
    .A2(net6120),
    .Y(_09996_),
    .B1(_09995_));
 sg13g2_a22oi_1 _18349_ (.Y(_09997_),
    .B1(_08633_),
    .B2(\atari2600.tia.diag[39] ),
    .A2(net6118),
    .A1(\atari2600.tia.diag[38] ));
 sg13g2_o21ai_1 _18350_ (.B1(_09997_),
    .Y(_09998_),
    .A1(_09987_),
    .A2(_09996_));
 sg13g2_o21ai_1 _18351_ (.B1(_09998_),
    .Y(_09999_),
    .A1(\atari2600.tia.diag[39] ),
    .A2(_08633_));
 sg13g2_nand4_1 _18352_ (.B(_09985_),
    .C(_09986_),
    .A(\atari2600.tia.enabl ),
    .Y(_10000_),
    .D(_09999_));
 sg13g2_nor2_2 _18353_ (.A(net6496),
    .B(net6490),
    .Y(_10001_));
 sg13g2_nand2_2 _18354_ (.Y(_10002_),
    .A(net6121),
    .B(net6120));
 sg13g2_a21oi_2 _18355_ (.B1(net6482),
    .Y(_10003_),
    .A2(_10002_),
    .A1(net6488));
 sg13g2_xor2_1 _18356_ (.B(net6498),
    .A(\atari2600.tia.refpf ),
    .X(_10004_));
 sg13g2_nand2_1 _18357_ (.Y(_10005_),
    .A(net6497),
    .B(_10003_));
 sg13g2_o21ai_1 _18358_ (.B1(_10005_),
    .Y(_10006_),
    .A1(_10003_),
    .A2(_10004_));
 sg13g2_nand2_1 _18359_ (.Y(_10007_),
    .A(_00140_),
    .B(_10003_));
 sg13g2_xor2_1 _18360_ (.B(net6502),
    .A(\atari2600.tia.refpf ),
    .X(_10008_));
 sg13g2_o21ai_1 _18361_ (.B1(_10007_),
    .Y(_10009_),
    .A1(_10003_),
    .A2(_10008_));
 sg13g2_mux2_1 _18362_ (.A0(\atari2600.tia.diag[91] ),
    .A1(\atari2600.tia.diag[90] ),
    .S(net5935),
    .X(_10010_));
 sg13g2_nor2_1 _18363_ (.A(\atari2600.tia.refpf ),
    .B(_10003_),
    .Y(_10011_));
 sg13g2_nor2_2 _18364_ (.A(net6496),
    .B(net6120),
    .Y(_10012_));
 sg13g2_nor2_2 _18365_ (.A(_08630_),
    .B(net6490),
    .Y(_10013_));
 sg13g2_nand2_2 _18366_ (.Y(_10014_),
    .A(net6496),
    .B(net6490));
 sg13g2_nand3_1 _18367_ (.B(_10011_),
    .C(_10014_),
    .A(_10002_),
    .Y(_10015_));
 sg13g2_o21ai_1 _18368_ (.B1(_10015_),
    .Y(_10016_),
    .A1(_08661_),
    .A2(_10011_));
 sg13g2_nand2b_1 _18369_ (.Y(_10017_),
    .B(net5935),
    .A_N(\atari2600.tia.diag[88] ));
 sg13g2_o21ai_1 _18370_ (.B1(_10017_),
    .Y(_10018_),
    .A1(\atari2600.tia.diag[89] ),
    .A2(net5935));
 sg13g2_nor2_2 _18371_ (.A(net6486),
    .B(net6483),
    .Y(_10019_));
 sg13g2_nor2_1 _18372_ (.A(net6495),
    .B(_10003_),
    .Y(_10020_));
 sg13g2_a21oi_2 _18373_ (.B1(_10020_),
    .Y(_10021_),
    .A2(net6072),
    .A1(net6495));
 sg13g2_mux2_1 _18374_ (.A0(\atari2600.tia.diag[83] ),
    .A1(\atari2600.tia.diag[82] ),
    .S(net5935),
    .X(_10022_));
 sg13g2_nand2b_1 _18375_ (.Y(_10023_),
    .B(net5935),
    .A_N(\atari2600.tia.diag[80] ));
 sg13g2_o21ai_1 _18376_ (.B1(_10023_),
    .Y(_10024_),
    .A1(\atari2600.tia.diag[81] ),
    .A2(net5935));
 sg13g2_nor2_2 _18377_ (.A(net6488),
    .B(_08633_),
    .Y(_10025_));
 sg13g2_o21ai_1 _18378_ (.B1(net6119),
    .Y(_10026_),
    .A1(\atari2600.tia.refpf ),
    .A2(net6121));
 sg13g2_mux2_1 _18379_ (.A0(_10025_),
    .A1(net6486),
    .S(_10026_),
    .X(_10027_));
 sg13g2_a21oi_2 _18380_ (.B1(_10027_),
    .Y(_10028_),
    .A2(_10003_),
    .A1(net6485));
 sg13g2_mux4_1 _18381_ (.S0(net5935),
    .A0(\atari2600.tia.diag[79] ),
    .A1(\atari2600.tia.diag[78] ),
    .A2(\atari2600.tia.diag[77] ),
    .A3(\atari2600.tia.diag[76] ),
    .S1(_10006_),
    .X(_10029_));
 sg13g2_nand2_1 _18382_ (.Y(_10030_),
    .A(_10021_),
    .B(_10029_));
 sg13g2_a21oi_1 _18383_ (.A1(_10006_),
    .A2(_10024_),
    .Y(_10031_),
    .B1(_10021_));
 sg13g2_o21ai_1 _18384_ (.B1(_10031_),
    .Y(_10032_),
    .A1(_10006_),
    .A2(_10022_));
 sg13g2_nand3_1 _18385_ (.B(_10030_),
    .C(_10032_),
    .A(_10016_),
    .Y(_10033_));
 sg13g2_a21oi_1 _18386_ (.A1(_10006_),
    .A2(_10018_),
    .Y(_10034_),
    .B1(_10021_));
 sg13g2_o21ai_1 _18387_ (.B1(_10034_),
    .Y(_10035_),
    .A1(_10006_),
    .A2(_10010_));
 sg13g2_mux4_1 _18388_ (.S0(net5935),
    .A0(\atari2600.tia.diag[87] ),
    .A1(\atari2600.tia.diag[86] ),
    .A2(\atari2600.tia.diag[85] ),
    .A3(\atari2600.tia.diag[84] ),
    .S1(_10006_),
    .X(_10036_));
 sg13g2_a21oi_1 _18389_ (.A1(_10021_),
    .A2(_10036_),
    .Y(_10037_),
    .B1(_10016_));
 sg13g2_a21oi_1 _18390_ (.A1(_10035_),
    .A2(_10037_),
    .Y(_10038_),
    .B1(_10028_));
 sg13g2_mux4_1 _18391_ (.S0(_10009_),
    .A0(\atari2600.tia.diag[95] ),
    .A1(\atari2600.tia.diag[94] ),
    .A2(\atari2600.tia.diag[93] ),
    .A3(\atari2600.tia.diag[92] ),
    .S1(_10006_),
    .X(_10039_));
 sg13g2_and3_1 _18392_ (.X(_10040_),
    .A(_10016_),
    .B(_10021_),
    .C(_10039_));
 sg13g2_a22oi_1 _18393_ (.Y(_10041_),
    .B1(_10040_),
    .B2(_10028_),
    .A2(_10038_),
    .A1(_10033_));
 sg13g2_or3_1 _18394_ (.A(net6118),
    .B(net6480),
    .C(_10001_),
    .X(_10042_));
 sg13g2_a21oi_1 _18395_ (.A1(net6482),
    .A2(_00139_),
    .Y(_10043_),
    .B1(\atari2600.tia.refpf ));
 sg13g2_o21ai_1 _18396_ (.B1(net6482),
    .Y(_10044_),
    .A1(net6490),
    .A2(net6488));
 sg13g2_a22oi_1 _18397_ (.Y(_10045_),
    .B1(net6071),
    .B2(\atari2600.tia.refpf ),
    .A2(_10043_),
    .A1(_10042_));
 sg13g2_nor2_1 _18398_ (.A(_10041_),
    .B(_10045_),
    .Y(_10046_));
 sg13g2_nor3_2 _18399_ (.A(_09647_),
    .B(_10041_),
    .C(_10045_),
    .Y(_10047_));
 sg13g2_nand2_1 _18400_ (.Y(_10048_),
    .A(net5758),
    .B(net5708));
 sg13g2_o21ai_1 _18401_ (.B1(_09938_),
    .Y(_00030_),
    .A1(net5539),
    .A2(_10048_));
 sg13g2_nand2_1 _18402_ (.Y(_10049_),
    .A(net3074),
    .B(net5737));
 sg13g2_o21ai_1 _18403_ (.B1(_10049_),
    .Y(_00031_),
    .A1(_09937_),
    .A2(net5539));
 sg13g2_a22oi_1 _18404_ (.Y(_10050_),
    .B1(net5286),
    .B2(_10047_),
    .A2(net5738),
    .A1(net3653));
 sg13g2_inv_1 _18405_ (.Y(_00032_),
    .A(_10050_));
 sg13g2_nor3_1 _18406_ (.A(_09647_),
    .B(net5287),
    .C(net5539),
    .Y(_10051_));
 sg13g2_a21o_1 _18407_ (.A2(net5738),
    .A1(net4105),
    .B1(_10051_),
    .X(_00033_));
 sg13g2_nand2_1 _18408_ (.Y(_10052_),
    .A(net3252),
    .B(net5737));
 sg13g2_o21ai_1 _18409_ (.B1(_10052_),
    .Y(_00034_),
    .A1(net5289),
    .A2(_10048_));
 sg13g2_nand2_1 _18410_ (.Y(_10053_),
    .A(net2972),
    .B(net5738));
 sg13g2_nand3_1 _18411_ (.B(_09640_),
    .C(net5758),
    .A(_09527_),
    .Y(_10054_));
 sg13g2_inv_1 _18412_ (.Y(_10055_),
    .A(_10054_));
 sg13g2_o21ai_1 _18413_ (.B1(_10053_),
    .Y(_00035_),
    .A1(net5539),
    .A2(_10054_));
 sg13g2_a22oi_1 _18414_ (.Y(_10056_),
    .B1(net5708),
    .B2(_10055_),
    .A2(net5737),
    .A1(net4479));
 sg13g2_inv_1 _18415_ (.Y(_00036_),
    .A(_10056_));
 sg13g2_nand2_1 _18416_ (.Y(_10057_),
    .A(net2992),
    .B(net5737));
 sg13g2_o21ai_1 _18417_ (.B1(_10057_),
    .Y(_00037_),
    .A1(_09815_),
    .A2(net5539));
 sg13g2_a22oi_1 _18418_ (.Y(_10058_),
    .B1(net5292),
    .B2(_10047_),
    .A2(net5738),
    .A1(net3303));
 sg13g2_inv_1 _18419_ (.Y(_00024_),
    .A(_10058_));
 sg13g2_nand2_1 _18420_ (.Y(_10059_),
    .A(net4142),
    .B(net5737));
 sg13g2_o21ai_1 _18421_ (.B1(_10059_),
    .Y(_00025_),
    .A1(net5262),
    .A2(_09937_));
 sg13g2_a22oi_1 _18422_ (.Y(_10060_),
    .B1(_09816_),
    .B2(net5286),
    .A2(net5737),
    .A1(net3240));
 sg13g2_inv_1 _18423_ (.Y(_00026_),
    .A(_10060_));
 sg13g2_nand2_1 _18424_ (.Y(_10061_),
    .A(net2999),
    .B(net5738));
 sg13g2_o21ai_1 _18425_ (.B1(net3000),
    .Y(_00027_),
    .A1(_09815_),
    .A2(net5289));
 sg13g2_nand2_1 _18426_ (.Y(_10062_),
    .A(net2959),
    .B(net5738));
 sg13g2_o21ai_1 _18427_ (.B1(net2960),
    .Y(_00028_),
    .A1(net5289),
    .A2(_10054_));
 sg13g2_nor2_2 _18428_ (.A(_09210_),
    .B(net5512),
    .Y(_10063_));
 sg13g2_nand2_2 _18429_ (.Y(_10064_),
    .A(net5402),
    .B(_09291_));
 sg13g2_nand3_1 _18430_ (.B(net5748),
    .C(_10063_),
    .A(_09127_),
    .Y(_10065_));
 sg13g2_nor2_1 _18431_ (.A(\atari2600.tia.vid_vsync ),
    .B(_10065_),
    .Y(_10066_));
 sg13g2_nor2_2 _18432_ (.A(net6540),
    .B(net5078),
    .Y(_10067_));
 sg13g2_o21ai_1 _18433_ (.B1(net6575),
    .Y(_10068_),
    .A1(\atari2600.tia.vid_vsync ),
    .A2(_10065_));
 sg13g2_nand2_2 _18434_ (.Y(_10069_),
    .A(_08626_),
    .B(net6124));
 sg13g2_nor2_2 _18435_ (.A(_08628_),
    .B(_08629_),
    .Y(_10070_));
 sg13g2_nand2_2 _18436_ (.Y(_10071_),
    .A(net6505),
    .B(net6507));
 sg13g2_nand4_1 _18437_ (.B(net6124),
    .C(net6121),
    .A(_08626_),
    .Y(_10072_),
    .D(net6067));
 sg13g2_and4_2 _18438_ (.A(net6490),
    .B(net6489),
    .C(net6481),
    .D(_10072_),
    .X(_10073_));
 sg13g2_nand4_1 _18439_ (.B(net6488),
    .C(net6481),
    .A(net6491),
    .Y(_10074_),
    .D(_10072_));
 sg13g2_nor2_1 _18440_ (.A(_09647_),
    .B(_10073_),
    .Y(_10075_));
 sg13g2_nor2_1 _18441_ (.A(_09472_),
    .B(net5706),
    .Y(_10076_));
 sg13g2_or2_1 _18442_ (.X(_10077_),
    .B(_10076_),
    .A(net2939));
 sg13g2_nand3_1 _18443_ (.B(_09646_),
    .C(_10073_),
    .A(net2939),
    .Y(_10078_));
 sg13g2_o21ai_1 _18444_ (.B1(_10078_),
    .Y(_00046_),
    .A1(_10068_),
    .A2(_10077_));
 sg13g2_nand2_1 _18445_ (.Y(_10079_),
    .A(\atari2600.tia.vid_ypos[1] ),
    .B(\atari2600.tia.vid_ypos[0] ));
 sg13g2_nand3_1 _18446_ (.B(_09646_),
    .C(_10079_),
    .A(_08702_),
    .Y(_10080_));
 sg13g2_a21oi_1 _18447_ (.A1(_10076_),
    .A2(_10080_),
    .Y(_10081_),
    .B1(net2949));
 sg13g2_nand2_1 _18448_ (.Y(_10082_),
    .A(_10067_),
    .B(_10081_));
 sg13g2_o21ai_1 _18449_ (.B1(_10082_),
    .Y(_00047_),
    .A1(_10074_),
    .A2(_10080_));
 sg13g2_xnor2_1 _18450_ (.Y(_10083_),
    .A(\atari2600.tia.vid_ypos[2] ),
    .B(_10079_));
 sg13g2_nand2_1 _18451_ (.Y(_10084_),
    .A(net5758),
    .B(_10083_));
 sg13g2_a21oi_1 _18452_ (.A1(_10076_),
    .A2(_10084_),
    .Y(_10085_),
    .B1(net3114));
 sg13g2_nand2_1 _18453_ (.Y(_10086_),
    .A(_10067_),
    .B(_10085_));
 sg13g2_o21ai_1 _18454_ (.B1(_10086_),
    .Y(_00048_),
    .A1(_10074_),
    .A2(_10084_));
 sg13g2_nor2_1 _18455_ (.A(net3114),
    .B(_10079_),
    .Y(_10087_));
 sg13g2_xnor2_1 _18456_ (.Y(_10088_),
    .A(\atari2600.tia.vid_ypos[3] ),
    .B(_10087_));
 sg13g2_a21oi_1 _18457_ (.A1(_10073_),
    .A2(_10088_),
    .Y(_10089_),
    .B1(_09647_));
 sg13g2_nor2_1 _18458_ (.A(_09472_),
    .B(_10089_),
    .Y(_10090_));
 sg13g2_nor3_1 _18459_ (.A(net4709),
    .B(_10068_),
    .C(_10090_),
    .Y(_10091_));
 sg13g2_a21o_1 _18460_ (.A2(_10089_),
    .A1(_10073_),
    .B1(_10091_),
    .X(_00049_));
 sg13g2_nand4_1 _18461_ (.B(\atari2600.tia.vid_ypos[2] ),
    .C(\atari2600.tia.vid_ypos[1] ),
    .A(\atari2600.tia.vid_ypos[3] ),
    .Y(_10092_),
    .D(\atari2600.tia.vid_ypos[0] ));
 sg13g2_o21ai_1 _18462_ (.B1(net5758),
    .Y(_10093_),
    .A1(_08571_),
    .A2(_10092_));
 sg13g2_a21oi_1 _18463_ (.A1(_08571_),
    .A2(_10092_),
    .Y(_10094_),
    .B1(_10093_));
 sg13g2_nor3_1 _18464_ (.A(_09472_),
    .B(net5706),
    .C(_10094_),
    .Y(_10095_));
 sg13g2_nor3_1 _18465_ (.A(net7127),
    .B(_10068_),
    .C(_10095_),
    .Y(_10096_));
 sg13g2_a21o_1 _18466_ (.A2(_10094_),
    .A1(_10073_),
    .B1(_10096_),
    .X(_00050_));
 sg13g2_o21ai_1 _18467_ (.B1(\atari2600.tia.vid_ypos[5] ),
    .Y(_10097_),
    .A1(_00160_),
    .A2(_10092_));
 sg13g2_nor3_1 _18468_ (.A(\atari2600.tia.vid_ypos[5] ),
    .B(_00160_),
    .C(_10092_),
    .Y(_10098_));
 sg13g2_nor2_1 _18469_ (.A(_10074_),
    .B(_10098_),
    .Y(_10099_));
 sg13g2_a21oi_1 _18470_ (.A1(_10097_),
    .A2(_10099_),
    .Y(_10100_),
    .B1(_09647_));
 sg13g2_nor2_1 _18471_ (.A(_09472_),
    .B(_10100_),
    .Y(_10101_));
 sg13g2_nor3_1 _18472_ (.A(net3456),
    .B(_10068_),
    .C(_10101_),
    .Y(_10102_));
 sg13g2_a21o_1 _18473_ (.A2(_10100_),
    .A1(_10073_),
    .B1(_10102_),
    .X(_00051_));
 sg13g2_or3_2 _18474_ (.A(_08570_),
    .B(_08571_),
    .C(_10092_),
    .X(_10103_));
 sg13g2_xnor2_1 _18475_ (.Y(_10104_),
    .A(\atari2600.tia.vid_ypos[6] ),
    .B(_10103_));
 sg13g2_o21ai_1 _18476_ (.B1(net5758),
    .Y(_10105_),
    .A1(_10074_),
    .A2(_10104_));
 sg13g2_a21oi_1 _18477_ (.A1(_09473_),
    .A2(_10105_),
    .Y(_10106_),
    .B1(net4536));
 sg13g2_nand2_1 _18478_ (.Y(_10107_),
    .A(_10067_),
    .B(_10106_));
 sg13g2_o21ai_1 _18479_ (.B1(_10107_),
    .Y(_00052_),
    .A1(_10074_),
    .A2(_10105_));
 sg13g2_o21ai_1 _18480_ (.B1(\atari2600.tia.vid_ypos[7] ),
    .Y(_10108_),
    .A1(_00161_),
    .A2(_10103_));
 sg13g2_nor3_1 _18481_ (.A(\atari2600.tia.vid_ypos[7] ),
    .B(_00161_),
    .C(_10103_),
    .Y(_10109_));
 sg13g2_nor2_1 _18482_ (.A(_10074_),
    .B(_10109_),
    .Y(_10110_));
 sg13g2_a21oi_1 _18483_ (.A1(_10108_),
    .A2(_10110_),
    .Y(_10111_),
    .B1(_09647_));
 sg13g2_nor2_1 _18484_ (.A(_09472_),
    .B(_10111_),
    .Y(_10112_));
 sg13g2_nor3_1 _18485_ (.A(net2963),
    .B(_10068_),
    .C(_10112_),
    .Y(_10113_));
 sg13g2_a21o_1 _18486_ (.A2(_10111_),
    .A1(_10073_),
    .B1(_10113_),
    .X(_00053_));
 sg13g2_nand2_1 _18487_ (.Y(_10114_),
    .A(\atari2600.tia.vid_ypos[7] ),
    .B(\atari2600.tia.vid_ypos[6] ));
 sg13g2_o21ai_1 _18488_ (.B1(\atari2600.tia.vid_ypos[8] ),
    .Y(_10115_),
    .A1(_10103_),
    .A2(_10114_));
 sg13g2_nor3_1 _18489_ (.A(\atari2600.tia.vid_ypos[8] ),
    .B(_10103_),
    .C(_10114_),
    .Y(_10116_));
 sg13g2_nor2_1 _18490_ (.A(_10074_),
    .B(_10116_),
    .Y(_10117_));
 sg13g2_a21oi_1 _18491_ (.A1(_10115_),
    .A2(_10117_),
    .Y(_10118_),
    .B1(_09647_));
 sg13g2_nor2_1 _18492_ (.A(_09472_),
    .B(_10118_),
    .Y(_10119_));
 sg13g2_nor3_1 _18493_ (.A(net7384),
    .B(_10068_),
    .C(_10119_),
    .Y(_10120_));
 sg13g2_a21o_1 _18494_ (.A2(_10118_),
    .A1(_10073_),
    .B1(_10120_),
    .X(_00054_));
 sg13g2_nand2_2 _18495_ (.Y(_10121_),
    .A(net6575),
    .B(_09647_));
 sg13g2_nor3_1 _18496_ (.A(net7542),
    .B(_10066_),
    .C(_10121_),
    .Y(_10122_));
 sg13g2_a21o_1 _18497_ (.A2(net5706),
    .A1(_08629_),
    .B1(_10122_),
    .X(_00038_));
 sg13g2_nor2_2 _18498_ (.A(net6504),
    .B(_08629_),
    .Y(_10123_));
 sg13g2_nand2_2 _18499_ (.Y(_10124_),
    .A(_08628_),
    .B(net6507));
 sg13g2_nor2_2 _18500_ (.A(_08628_),
    .B(net6507),
    .Y(_10125_));
 sg13g2_nand2_2 _18501_ (.Y(_10126_),
    .A(net6504),
    .B(_08629_));
 sg13g2_o21ai_1 _18502_ (.B1(net5706),
    .Y(_10127_),
    .A1(_10123_),
    .A2(_10125_));
 sg13g2_or2_1 _18503_ (.X(_10128_),
    .B(_10121_),
    .A(net7547));
 sg13g2_o21ai_1 _18504_ (.B1(_10127_),
    .Y(_00039_),
    .A1(net5078),
    .A2(_10128_));
 sg13g2_nor2_1 _18505_ (.A(_00140_),
    .B(net6067),
    .Y(_10129_));
 sg13g2_nand2_1 _18506_ (.Y(_10130_),
    .A(_00140_),
    .B(net6067));
 sg13g2_nand2_1 _18507_ (.Y(_10131_),
    .A(net5706),
    .B(_10130_));
 sg13g2_or3_1 _18508_ (.A(_00140_),
    .B(net5078),
    .C(_10121_),
    .X(_10132_));
 sg13g2_o21ai_1 _18509_ (.B1(_10132_),
    .Y(_00040_),
    .A1(_10129_),
    .A2(_10131_));
 sg13g2_xnor2_1 _18510_ (.Y(_10133_),
    .A(net6497),
    .B(_10129_));
 sg13g2_nor3_1 _18511_ (.A(net6497),
    .B(net5078),
    .C(_10121_),
    .Y(_10134_));
 sg13g2_a21o_1 _18512_ (.A2(_10133_),
    .A1(net5706),
    .B1(_10134_),
    .X(_00041_));
 sg13g2_nand2_1 _18513_ (.Y(_10135_),
    .A(net6503),
    .B(_10070_));
 sg13g2_nand2_2 _18514_ (.Y(_10136_),
    .A(net6501),
    .B(net6503));
 sg13g2_or2_2 _18515_ (.X(_10137_),
    .B(_10136_),
    .A(_10071_));
 sg13g2_nor2_1 _18516_ (.A(net6493),
    .B(net6029),
    .Y(_10138_));
 sg13g2_xor2_1 _18517_ (.B(net6029),
    .A(net6493),
    .X(_10139_));
 sg13g2_nor3_1 _18518_ (.A(net6493),
    .B(net5078),
    .C(_10121_),
    .Y(_10140_));
 sg13g2_a21o_1 _18519_ (.A2(_10139_),
    .A1(net5706),
    .B1(_10140_),
    .X(_00042_));
 sg13g2_xnor2_1 _18520_ (.Y(_10141_),
    .A(_00142_),
    .B(_10138_));
 sg13g2_nor3_1 _18521_ (.A(_00142_),
    .B(net5078),
    .C(_10121_),
    .Y(_10142_));
 sg13g2_a21o_1 _18522_ (.A2(_10141_),
    .A1(net5706),
    .B1(_10142_),
    .X(_00043_));
 sg13g2_nor3_1 _18523_ (.A(net6485),
    .B(_10014_),
    .C(net6029),
    .Y(_10143_));
 sg13g2_o21ai_1 _18524_ (.B1(net6484),
    .Y(_10144_),
    .A1(_10014_),
    .A2(net6029));
 sg13g2_nand2_1 _18525_ (.Y(_10145_),
    .A(_10075_),
    .B(_10144_));
 sg13g2_or3_1 _18526_ (.A(net6484),
    .B(net5078),
    .C(_10121_),
    .X(_10146_));
 sg13g2_o21ai_1 _18527_ (.B1(_10146_),
    .Y(_00044_),
    .A1(_10143_),
    .A2(_10145_));
 sg13g2_xnor2_1 _18528_ (.Y(_10147_),
    .A(net6480),
    .B(_10143_));
 sg13g2_nor3_1 _18529_ (.A(net6480),
    .B(net5078),
    .C(_10121_),
    .Y(_10148_));
 sg13g2_a21o_1 _18530_ (.A2(_10147_),
    .A1(_10075_),
    .B1(_10148_),
    .X(_00045_));
 sg13g2_a22oi_1 _18531_ (.Y(_10149_),
    .B1(net5298),
    .B2(\atari2600.ram[50][0] ),
    .A2(net5438),
    .A1(\atari2600.ram[49][0] ));
 sg13g2_a221oi_1 _18532_ (.B2(\atari2600.ram[51][0] ),
    .C1(net5280),
    .B1(net5346),
    .A1(\atari2600.ram[48][0] ),
    .Y(_10150_),
    .A2(net5391));
 sg13g2_a21oi_1 _18533_ (.A1(_10149_),
    .A2(_10150_),
    .Y(_10151_),
    .B1(_09293_));
 sg13g2_a22oi_1 _18534_ (.Y(_10152_),
    .B1(net5394),
    .B2(\atari2600.ram[56][0] ),
    .A2(net5443),
    .A1(\atari2600.ram[57][0] ));
 sg13g2_a22oi_1 _18535_ (.Y(_10153_),
    .B1(net5303),
    .B2(\atari2600.ram[58][0] ),
    .A2(net5349),
    .A1(\atari2600.ram[59][0] ));
 sg13g2_a21oi_1 _18536_ (.A1(_10152_),
    .A2(_10153_),
    .Y(_10154_),
    .B1(net5480));
 sg13g2_a22oi_1 _18537_ (.Y(_10155_),
    .B1(net5347),
    .B2(\atari2600.ram[63][0] ),
    .A2(net5393),
    .A1(\atari2600.ram[60][0] ));
 sg13g2_a22oi_1 _18538_ (.Y(_10156_),
    .B1(net5301),
    .B2(\atari2600.ram[62][0] ),
    .A2(net5441),
    .A1(\atari2600.ram[61][0] ));
 sg13g2_a21oi_1 _18539_ (.A1(_10155_),
    .A2(_10156_),
    .Y(_10157_),
    .B1(net5488));
 sg13g2_a22oi_1 _18540_ (.Y(_10158_),
    .B1(net5346),
    .B2(\atari2600.ram[55][0] ),
    .A2(net5391),
    .A1(\atari2600.ram[52][0] ));
 sg13g2_a22oi_1 _18541_ (.Y(_10159_),
    .B1(net5298),
    .B2(\atari2600.ram[54][0] ),
    .A2(net5438),
    .A1(\atari2600.ram[53][0] ));
 sg13g2_a21oi_1 _18542_ (.A1(_10158_),
    .A2(_10159_),
    .Y(_10160_),
    .B1(net5518));
 sg13g2_nor4_1 _18543_ (.A(_10151_),
    .B(_10154_),
    .C(_10157_),
    .D(_10160_),
    .Y(_10161_));
 sg13g2_a22oi_1 _18544_ (.Y(_10162_),
    .B1(net5385),
    .B2(\atari2600.ram[36][0] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][0] ));
 sg13g2_a22oi_1 _18545_ (.Y(_10163_),
    .B1(net5293),
    .B2(\atari2600.ram[38][0] ),
    .A2(net5340),
    .A1(\atari2600.ram[39][0] ));
 sg13g2_a21oi_2 _18546_ (.B1(net5515),
    .Y(_10164_),
    .A2(_10163_),
    .A1(_10162_));
 sg13g2_a22oi_1 _18547_ (.Y(_10165_),
    .B1(net5344),
    .B2(\atari2600.ram[43][0] ),
    .A2(net5389),
    .A1(\atari2600.ram[40][0] ));
 sg13g2_a22oi_1 _18548_ (.Y(_10166_),
    .B1(net5297),
    .B2(\atari2600.ram[42][0] ),
    .A2(net5437),
    .A1(\atari2600.ram[41][0] ));
 sg13g2_a21oi_1 _18549_ (.A1(_10165_),
    .A2(_10166_),
    .Y(_10167_),
    .B1(net5477));
 sg13g2_a22oi_1 _18550_ (.Y(_10168_),
    .B1(net5342),
    .B2(\atari2600.ram[47][0] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][0] ));
 sg13g2_a22oi_1 _18551_ (.Y(_10169_),
    .B1(net5305),
    .B2(\atari2600.ram[46][0] ),
    .A2(net5445),
    .A1(\atari2600.ram[45][0] ));
 sg13g2_a21oi_1 _18552_ (.A1(_10168_),
    .A2(_10169_),
    .Y(_10170_),
    .B1(net5490));
 sg13g2_a22oi_1 _18553_ (.Y(_10171_),
    .B1(net5341),
    .B2(\atari2600.ram[35][0] ),
    .A2(net5386),
    .A1(\atari2600.ram[32][0] ));
 sg13g2_a22oi_1 _18554_ (.Y(_10172_),
    .B1(net5294),
    .B2(\atari2600.ram[34][0] ),
    .A2(net5434),
    .A1(\atari2600.ram[33][0] ));
 sg13g2_a21oi_1 _18555_ (.A1(_10171_),
    .A2(_10172_),
    .Y(_10173_),
    .B1(net5501));
 sg13g2_or2_1 _18556_ (.X(_10174_),
    .B(_10173_),
    .A(_10170_));
 sg13g2_nor4_2 _18557_ (.A(net5275),
    .B(_10164_),
    .C(_10167_),
    .Y(_10175_),
    .D(_10174_));
 sg13g2_nor3_2 _18558_ (.A(net5568),
    .B(_10161_),
    .C(_10175_),
    .Y(_10176_));
 sg13g2_a22oi_1 _18559_ (.Y(_10177_),
    .B1(net5344),
    .B2(\atari2600.ram[11][0] ),
    .A2(net5390),
    .A1(\atari2600.ram[8][0] ));
 sg13g2_a22oi_1 _18560_ (.Y(_10178_),
    .B1(net5296),
    .B2(\atari2600.ram[10][0] ),
    .A2(net5436),
    .A1(\atari2600.ram[9][0] ));
 sg13g2_a21oi_2 _18561_ (.B1(net5479),
    .Y(_10179_),
    .A2(_10178_),
    .A1(_10177_));
 sg13g2_a22oi_1 _18562_ (.Y(_10180_),
    .B1(net5354),
    .B2(\atari2600.ram[7][0] ),
    .A2(net5399),
    .A1(\atari2600.ram[4][0] ));
 sg13g2_a22oi_1 _18563_ (.Y(_10181_),
    .B1(net5308),
    .B2(\atari2600.ram[6][0] ),
    .A2(net5448),
    .A1(\atari2600.ram[5][0] ));
 sg13g2_a21oi_1 _18564_ (.A1(_10180_),
    .A2(_10181_),
    .Y(_10182_),
    .B1(net5516));
 sg13g2_a22oi_1 _18565_ (.Y(_10183_),
    .B1(net5354),
    .B2(\atari2600.ram[15][0] ),
    .A2(net5399),
    .A1(\atari2600.ram[12][0] ));
 sg13g2_a22oi_1 _18566_ (.Y(_10184_),
    .B1(net5306),
    .B2(\atari2600.ram[14][0] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][0] ));
 sg13g2_a21oi_1 _18567_ (.A1(_10183_),
    .A2(_10184_),
    .Y(_10185_),
    .B1(net5491));
 sg13g2_a22oi_1 _18568_ (.Y(_10186_),
    .B1(net5353),
    .B2(\atari2600.ram[3][0] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][0] ));
 sg13g2_a22oi_1 _18569_ (.Y(_10187_),
    .B1(net5308),
    .B2(\atari2600.ram[2][0] ),
    .A2(net5448),
    .A1(\atari2600.ram[1][0] ));
 sg13g2_a21oi_2 _18570_ (.B1(net5507),
    .Y(_10188_),
    .A2(_10187_),
    .A1(_10186_));
 sg13g2_nor4_1 _18571_ (.A(_10179_),
    .B(_10182_),
    .C(_10185_),
    .D(_10188_),
    .Y(_10189_));
 sg13g2_a22oi_1 _18572_ (.Y(_10190_),
    .B1(net5373),
    .B2(\atari2600.ram[31][0] ),
    .A2(net5421),
    .A1(\atari2600.ram[28][0] ));
 sg13g2_a22oi_1 _18573_ (.Y(_10191_),
    .B1(net5328),
    .B2(\atari2600.ram[30][0] ),
    .A2(net5467),
    .A1(\atari2600.ram[29][0] ));
 sg13g2_a21oi_1 _18574_ (.A1(_10190_),
    .A2(_10191_),
    .Y(_10192_),
    .B1(net5498));
 sg13g2_a22oi_1 _18575_ (.Y(_10193_),
    .B1(net5373),
    .B2(\atari2600.ram[19][0] ),
    .A2(net5421),
    .A1(\atari2600.ram[16][0] ));
 sg13g2_a22oi_1 _18576_ (.Y(_10194_),
    .B1(net5328),
    .B2(\atari2600.ram[18][0] ),
    .A2(net5467),
    .A1(\atari2600.ram[17][0] ));
 sg13g2_a21oi_1 _18577_ (.A1(_10193_),
    .A2(_10194_),
    .Y(_10195_),
    .B1(net5505));
 sg13g2_a22oi_1 _18578_ (.Y(_10196_),
    .B1(net5356),
    .B2(\atari2600.ram[23][0] ),
    .A2(net5403),
    .A1(\atari2600.ram[20][0] ));
 sg13g2_a22oi_1 _18579_ (.Y(_10197_),
    .B1(net5309),
    .B2(\atari2600.ram[22][0] ),
    .A2(net5449),
    .A1(\atari2600.ram[21][0] ));
 sg13g2_a21oi_1 _18580_ (.A1(_10196_),
    .A2(_10197_),
    .Y(_10198_),
    .B1(net5517));
 sg13g2_a22oi_1 _18581_ (.Y(_10199_),
    .B1(net5372),
    .B2(\atari2600.ram[27][0] ),
    .A2(net5420),
    .A1(\atari2600.ram[24][0] ));
 sg13g2_a22oi_1 _18582_ (.Y(_10200_),
    .B1(net5327),
    .B2(\atari2600.ram[26][0] ),
    .A2(net5466),
    .A1(\atari2600.ram[25][0] ));
 sg13g2_a21oi_2 _18583_ (.B1(net5484),
    .Y(_10201_),
    .A2(_10200_),
    .A1(_10199_));
 sg13g2_nor4_2 _18584_ (.A(_10192_),
    .B(_10195_),
    .C(_10198_),
    .Y(_10202_),
    .D(_10201_));
 sg13g2_nor2_1 _18585_ (.A(net5265),
    .B(_10202_),
    .Y(_10203_));
 sg13g2_o21ai_1 _18586_ (.B1(net5543),
    .Y(_10204_),
    .A1(net5270),
    .A2(_10189_));
 sg13g2_nor3_1 _18587_ (.A(_10176_),
    .B(_10203_),
    .C(_10204_),
    .Y(_10205_));
 sg13g2_a22oi_1 _18588_ (.Y(_10206_),
    .B1(net5413),
    .B2(\atari2600.ram[100][0] ),
    .A2(net5460),
    .A1(\atari2600.ram[101][0] ));
 sg13g2_a22oi_1 _18589_ (.Y(_10207_),
    .B1(net5321),
    .B2(\atari2600.ram[102][0] ),
    .A2(net5366),
    .A1(\atari2600.ram[103][0] ));
 sg13g2_a21oi_1 _18590_ (.A1(_10206_),
    .A2(_10207_),
    .Y(_10208_),
    .B1(net5526));
 sg13g2_a22oi_1 _18591_ (.Y(_10209_),
    .B1(net5365),
    .B2(\atari2600.ram[111][0] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][0] ));
 sg13g2_a22oi_1 _18592_ (.Y(_10210_),
    .B1(net5319),
    .B2(\atari2600.ram[110][0] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][0] ));
 sg13g2_a21oi_1 _18593_ (.A1(_10209_),
    .A2(_10210_),
    .Y(_10211_),
    .B1(net5495));
 sg13g2_a22oi_1 _18594_ (.Y(_10212_),
    .B1(net5369),
    .B2(\atari2600.ram[99][0] ),
    .A2(net5416),
    .A1(\atari2600.ram[96][0] ));
 sg13g2_a22oi_1 _18595_ (.Y(_10213_),
    .B1(net5322),
    .B2(\atari2600.ram[98][0] ),
    .A2(net5464),
    .A1(\atari2600.ram[97][0] ));
 sg13g2_a21oi_1 _18596_ (.A1(_10212_),
    .A2(_10213_),
    .Y(_10214_),
    .B1(net5510));
 sg13g2_a22oi_1 _18597_ (.Y(_10215_),
    .B1(net5361),
    .B2(\atari2600.ram[107][0] ),
    .A2(net5406),
    .A1(\atari2600.ram[104][0] ));
 sg13g2_a22oi_1 _18598_ (.Y(_10216_),
    .B1(net5314),
    .B2(\atari2600.ram[106][0] ),
    .A2(net5453),
    .A1(\atari2600.ram[105][0] ));
 sg13g2_a21oi_1 _18599_ (.A1(_10215_),
    .A2(_10216_),
    .Y(_10217_),
    .B1(net5483));
 sg13g2_nor2_1 _18600_ (.A(net5276),
    .B(_10214_),
    .Y(_10218_));
 sg13g2_nor3_2 _18601_ (.A(_10208_),
    .B(_10211_),
    .C(_10217_),
    .Y(_10219_));
 sg13g2_a22oi_1 _18602_ (.Y(_10220_),
    .B1(net5364),
    .B2(\atari2600.ram[123][0] ),
    .A2(net5409),
    .A1(\atari2600.ram[120][0] ));
 sg13g2_a22oi_1 _18603_ (.Y(_10221_),
    .B1(net5316),
    .B2(\atari2600.ram[122][0] ),
    .A2(net5455),
    .A1(\atari2600.ram[121][0] ));
 sg13g2_a21oi_1 _18604_ (.A1(_10220_),
    .A2(_10221_),
    .Y(_10222_),
    .B1(net5482));
 sg13g2_a22oi_1 _18605_ (.Y(_10223_),
    .B1(net5362),
    .B2(\atari2600.ram[115][0] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][0] ));
 sg13g2_a22oi_1 _18606_ (.Y(_10224_),
    .B1(net5317),
    .B2(\atari2600.ram[114][0] ),
    .A2(net5456),
    .A1(\atari2600.ram[113][0] ));
 sg13g2_a21oi_1 _18607_ (.A1(_10223_),
    .A2(_10224_),
    .Y(_10225_),
    .B1(net5510));
 sg13g2_a22oi_1 _18608_ (.Y(_10226_),
    .B1(net5359),
    .B2(\atari2600.ram[127][0] ),
    .A2(net5406),
    .A1(\atari2600.ram[124][0] ));
 sg13g2_a22oi_1 _18609_ (.Y(_10227_),
    .B1(net5314),
    .B2(\atari2600.ram[126][0] ),
    .A2(net5453),
    .A1(\atari2600.ram[125][0] ));
 sg13g2_a21o_2 _18610_ (.A2(_10227_),
    .A1(_10226_),
    .B1(net5494),
    .X(_10228_));
 sg13g2_a22oi_1 _18611_ (.Y(_10229_),
    .B1(net5409),
    .B2(\atari2600.ram[116][0] ),
    .A2(net5455),
    .A1(\atari2600.ram[117][0] ));
 sg13g2_a22oi_1 _18612_ (.Y(_10230_),
    .B1(net5316),
    .B2(\atari2600.ram[118][0] ),
    .A2(net5364),
    .A1(\atari2600.ram[119][0] ));
 sg13g2_a21oi_1 _18613_ (.A1(_10229_),
    .A2(_10230_),
    .Y(_10231_),
    .B1(net5520));
 sg13g2_nor4_1 _18614_ (.A(net5283),
    .B(_10222_),
    .C(_10225_),
    .D(_10231_),
    .Y(_10232_));
 sg13g2_a221oi_1 _18615_ (.B2(_10232_),
    .C1(net5572),
    .B1(_10228_),
    .A1(_10218_),
    .Y(_10233_),
    .A2(_10219_));
 sg13g2_a22oi_1 _18616_ (.Y(_10234_),
    .B1(net5368),
    .B2(\atari2600.ram[75][0] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][0] ));
 sg13g2_a22oi_1 _18617_ (.Y(_10235_),
    .B1(net5323),
    .B2(\atari2600.ram[74][0] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][0] ));
 sg13g2_a21oi_2 _18618_ (.B1(net5485),
    .Y(_10236_),
    .A2(_10235_),
    .A1(_10234_));
 sg13g2_a22oi_1 _18619_ (.Y(_10237_),
    .B1(net5367),
    .B2(\atari2600.ram[79][0] ),
    .A2(net5418),
    .A1(\atari2600.ram[76][0] ));
 sg13g2_a22oi_1 _18620_ (.Y(_10238_),
    .B1(net5320),
    .B2(\atari2600.ram[78][0] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][0] ));
 sg13g2_a21oi_2 _18621_ (.B1(net5496),
    .Y(_10239_),
    .A2(_10238_),
    .A1(_10237_));
 sg13g2_a22oi_1 _18622_ (.Y(_10240_),
    .B1(net5378),
    .B2(\atari2600.ram[67][0] ),
    .A2(net5426),
    .A1(\atari2600.ram[64][0] ));
 sg13g2_a22oi_1 _18623_ (.Y(_10241_),
    .B1(net5331),
    .B2(\atari2600.ram[66][0] ),
    .A2(net5470),
    .A1(\atari2600.ram[65][0] ));
 sg13g2_a21oi_1 _18624_ (.A1(_10240_),
    .A2(_10241_),
    .Y(_10242_),
    .B1(net5512));
 sg13g2_a22oi_1 _18625_ (.Y(_10243_),
    .B1(net5378),
    .B2(\atari2600.ram[71][0] ),
    .A2(net5427),
    .A1(\atari2600.ram[68][0] ));
 sg13g2_a22oi_1 _18626_ (.Y(_10244_),
    .B1(net5336),
    .B2(\atari2600.ram[70][0] ),
    .A2(net5475),
    .A1(\atari2600.ram[69][0] ));
 sg13g2_a21oi_2 _18627_ (.B1(net5524),
    .Y(_10245_),
    .A2(_10244_),
    .A1(_10243_));
 sg13g2_nor4_2 _18628_ (.A(_10236_),
    .B(_10239_),
    .C(_10242_),
    .Y(_10246_),
    .D(_10245_));
 sg13g2_nor2_1 _18629_ (.A(net5271),
    .B(_10246_),
    .Y(_10247_));
 sg13g2_a22oi_1 _18630_ (.Y(_10248_),
    .B1(net5380),
    .B2(\atari2600.ram[87][0] ),
    .A2(net5428),
    .A1(\atari2600.ram[84][0] ));
 sg13g2_a22oi_1 _18631_ (.Y(_10249_),
    .B1(net5333),
    .B2(\atari2600.ram[86][0] ),
    .A2(net5472),
    .A1(\atari2600.ram[85][0] ));
 sg13g2_a21oi_1 _18632_ (.A1(_10248_),
    .A2(_10249_),
    .Y(_10250_),
    .B1(net5523));
 sg13g2_a22oi_1 _18633_ (.Y(_10251_),
    .B1(net5381),
    .B2(\atari2600.ram[91][0] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][0] ));
 sg13g2_a22oi_1 _18634_ (.Y(_10252_),
    .B1(net5334),
    .B2(\atari2600.ram[90][0] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][0] ));
 sg13g2_a21oi_1 _18635_ (.A1(_10251_),
    .A2(_10252_),
    .Y(_10253_),
    .B1(net5484));
 sg13g2_a22oi_1 _18636_ (.Y(_10254_),
    .B1(net5374),
    .B2(\atari2600.ram[83][0] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][0] ));
 sg13g2_a22oi_1 _18637_ (.Y(_10255_),
    .B1(net5329),
    .B2(\atari2600.ram[82][0] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][0] ));
 sg13g2_a21oi_1 _18638_ (.A1(_10254_),
    .A2(_10255_),
    .Y(_10256_),
    .B1(net5508));
 sg13g2_a22oi_1 _18639_ (.Y(_10257_),
    .B1(net5379),
    .B2(\atari2600.ram[95][0] ),
    .A2(net5427),
    .A1(\atari2600.ram[92][0] ));
 sg13g2_a22oi_1 _18640_ (.Y(_10258_),
    .B1(net5333),
    .B2(\atari2600.ram[94][0] ),
    .A2(net5472),
    .A1(\atari2600.ram[93][0] ));
 sg13g2_a21oi_1 _18641_ (.A1(_10257_),
    .A2(_10258_),
    .Y(_10259_),
    .B1(net5498));
 sg13g2_nor4_2 _18642_ (.A(_10250_),
    .B(_10253_),
    .C(_10256_),
    .Y(_10260_),
    .D(_10259_));
 sg13g2_o21ai_1 _18643_ (.B1(net5546),
    .Y(_10261_),
    .A1(net5266),
    .A2(_10260_));
 sg13g2_nor3_2 _18644_ (.A(_10233_),
    .B(_10247_),
    .C(_10261_),
    .Y(_10262_));
 sg13g2_nor2_1 _18645_ (.A(_10205_),
    .B(_10262_),
    .Y(_00001_));
 sg13g2_a22oi_1 _18646_ (.Y(_10263_),
    .B1(net5350),
    .B2(\atari2600.ram[115][1] ),
    .A2(net5395),
    .A1(\atari2600.ram[112][1] ));
 sg13g2_a22oi_1 _18647_ (.Y(_10264_),
    .B1(net5313),
    .B2(\atari2600.ram[114][1] ),
    .A2(net5441),
    .A1(\atari2600.ram[113][1] ));
 sg13g2_a21oi_1 _18648_ (.A1(_10263_),
    .A2(_10264_),
    .Y(_10265_),
    .B1(net5506));
 sg13g2_a22oi_1 _18649_ (.Y(_10266_),
    .B1(net5360),
    .B2(\atari2600.ram[127][1] ),
    .A2(net5407),
    .A1(\atari2600.ram[124][1] ));
 sg13g2_a22oi_1 _18650_ (.Y(_10267_),
    .B1(net5312),
    .B2(\atari2600.ram[126][1] ),
    .A2(net5452),
    .A1(\atari2600.ram[125][1] ));
 sg13g2_a21oi_2 _18651_ (.B1(net5489),
    .Y(_10268_),
    .A2(_10267_),
    .A1(_10266_));
 sg13g2_a22oi_1 _18652_ (.Y(_10269_),
    .B1(net5411),
    .B2(\atari2600.ram[116][1] ),
    .A2(net5453),
    .A1(\atari2600.ram[117][1] ));
 sg13g2_a22oi_1 _18653_ (.Y(_10270_),
    .B1(net5314),
    .B2(\atari2600.ram[118][1] ),
    .A2(net5361),
    .A1(\atari2600.ram[119][1] ));
 sg13g2_a21o_1 _18654_ (.A2(_10270_),
    .A1(_10269_),
    .B1(net5521),
    .X(_10271_));
 sg13g2_a22oi_1 _18655_ (.Y(_10272_),
    .B1(net5350),
    .B2(\atari2600.ram[123][1] ),
    .A2(net5395),
    .A1(\atari2600.ram[120][1] ));
 sg13g2_a22oi_1 _18656_ (.Y(_10273_),
    .B1(net5303),
    .B2(\atari2600.ram[122][1] ),
    .A2(net5443),
    .A1(\atari2600.ram[121][1] ));
 sg13g2_a21oi_2 _18657_ (.B1(net5480),
    .Y(_10274_),
    .A2(_10273_),
    .A1(_10272_));
 sg13g2_nor4_2 _18658_ (.A(net5281),
    .B(_10265_),
    .C(_10268_),
    .Y(_10275_),
    .D(_10274_));
 sg13g2_a22oi_1 _18659_ (.Y(_10276_),
    .B1(net5363),
    .B2(\atari2600.ram[107][1] ),
    .A2(net5409),
    .A1(\atari2600.ram[104][1] ));
 sg13g2_a22oi_1 _18660_ (.Y(_10277_),
    .B1(net5316),
    .B2(\atari2600.ram[106][1] ),
    .A2(net5455),
    .A1(\atari2600.ram[105][1] ));
 sg13g2_a21oi_1 _18661_ (.A1(_10276_),
    .A2(_10277_),
    .Y(_10278_),
    .B1(net5483));
 sg13g2_nor2_1 _18662_ (.A(net5276),
    .B(_10278_),
    .Y(_10279_));
 sg13g2_a22oi_1 _18663_ (.Y(_10280_),
    .B1(net5365),
    .B2(\atari2600.ram[111][1] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][1] ));
 sg13g2_a22oi_1 _18664_ (.Y(_10281_),
    .B1(net5319),
    .B2(\atari2600.ram[110][1] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][1] ));
 sg13g2_a21oi_2 _18665_ (.B1(net5495),
    .Y(_10282_),
    .A2(_10281_),
    .A1(_10280_));
 sg13g2_a22oi_1 _18666_ (.Y(_10283_),
    .B1(net5413),
    .B2(\atari2600.ram[100][1] ),
    .A2(net5458),
    .A1(\atari2600.ram[101][1] ));
 sg13g2_a22oi_1 _18667_ (.Y(_10284_),
    .B1(net5319),
    .B2(\atari2600.ram[102][1] ),
    .A2(net5366),
    .A1(\atari2600.ram[103][1] ));
 sg13g2_a21oi_1 _18668_ (.A1(_10283_),
    .A2(_10284_),
    .Y(_10285_),
    .B1(net5526));
 sg13g2_a22oi_1 _18669_ (.Y(_10286_),
    .B1(net5369),
    .B2(\atari2600.ram[99][1] ),
    .A2(net5416),
    .A1(\atari2600.ram[96][1] ));
 sg13g2_a22oi_1 _18670_ (.Y(_10287_),
    .B1(net5325),
    .B2(\atari2600.ram[98][1] ),
    .A2(net5461),
    .A1(\atari2600.ram[97][1] ));
 sg13g2_a21oi_2 _18671_ (.B1(net5511),
    .Y(_10288_),
    .A2(_10287_),
    .A1(_10286_));
 sg13g2_nor3_2 _18672_ (.A(_10282_),
    .B(_10285_),
    .C(_10288_),
    .Y(_10289_));
 sg13g2_a221oi_1 _18673_ (.B2(_10289_),
    .C1(net5571),
    .B1(_10279_),
    .A1(_10271_),
    .Y(_10290_),
    .A2(_10275_));
 sg13g2_a22oi_1 _18674_ (.Y(_10291_),
    .B1(net5372),
    .B2(\atari2600.ram[95][1] ),
    .A2(net5420),
    .A1(\atari2600.ram[92][1] ));
 sg13g2_a22oi_1 _18675_ (.Y(_10292_),
    .B1(net5327),
    .B2(\atari2600.ram[94][1] ),
    .A2(net5466),
    .A1(\atari2600.ram[93][1] ));
 sg13g2_a21oi_2 _18676_ (.B1(net5498),
    .Y(_10293_),
    .A2(_10292_),
    .A1(_10291_));
 sg13g2_a22oi_1 _18677_ (.Y(_10294_),
    .B1(net5381),
    .B2(\atari2600.ram[91][1] ),
    .A2(net5429),
    .A1(\atari2600.ram[88][1] ));
 sg13g2_a22oi_1 _18678_ (.Y(_10295_),
    .B1(net5334),
    .B2(\atari2600.ram[90][1] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][1] ));
 sg13g2_a21oi_1 _18679_ (.A1(_10294_),
    .A2(_10295_),
    .Y(_10296_),
    .B1(net5484));
 sg13g2_a22oi_1 _18680_ (.Y(_10297_),
    .B1(net5381),
    .B2(\atari2600.ram[87][1] ),
    .A2(net5429),
    .A1(\atari2600.ram[84][1] ));
 sg13g2_a22oi_1 _18681_ (.Y(_10298_),
    .B1(net5335),
    .B2(\atari2600.ram[86][1] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][1] ));
 sg13g2_a21oi_2 _18682_ (.B1(net5525),
    .Y(_10299_),
    .A2(_10298_),
    .A1(_10297_));
 sg13g2_a22oi_1 _18683_ (.Y(_10300_),
    .B1(net5375),
    .B2(\atari2600.ram[83][1] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][1] ));
 sg13g2_a22oi_1 _18684_ (.Y(_10301_),
    .B1(net5330),
    .B2(\atari2600.ram[82][1] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][1] ));
 sg13g2_a21oi_1 _18685_ (.A1(_10300_),
    .A2(_10301_),
    .Y(_10302_),
    .B1(net5509));
 sg13g2_nor4_2 _18686_ (.A(_10293_),
    .B(_10296_),
    .C(_10299_),
    .Y(_10303_),
    .D(_10302_));
 sg13g2_a22oi_1 _18687_ (.Y(_10304_),
    .B1(net5367),
    .B2(\atari2600.ram[79][1] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][1] ));
 sg13g2_a22oi_1 _18688_ (.Y(_10305_),
    .B1(net5320),
    .B2(\atari2600.ram[78][1] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][1] ));
 sg13g2_a21oi_2 _18689_ (.B1(net5496),
    .Y(_10306_),
    .A2(_10305_),
    .A1(_10304_));
 sg13g2_a22oi_1 _18690_ (.Y(_10307_),
    .B1(net5369),
    .B2(\atari2600.ram[67][1] ),
    .A2(net5416),
    .A1(\atari2600.ram[64][1] ));
 sg13g2_a22oi_1 _18691_ (.Y(_10308_),
    .B1(net5324),
    .B2(\atari2600.ram[66][1] ),
    .A2(net5463),
    .A1(\atari2600.ram[65][1] ));
 sg13g2_a21oi_1 _18692_ (.A1(_10307_),
    .A2(_10308_),
    .Y(_10309_),
    .B1(net5511));
 sg13g2_a22oi_1 _18693_ (.Y(_10310_),
    .B1(net5379),
    .B2(\atari2600.ram[71][1] ),
    .A2(net5426),
    .A1(\atari2600.ram[68][1] ));
 sg13g2_a22oi_1 _18694_ (.Y(_10311_),
    .B1(net5331),
    .B2(\atari2600.ram[70][1] ),
    .A2(net5470),
    .A1(\atari2600.ram[69][1] ));
 sg13g2_a21oi_1 _18695_ (.A1(_10310_),
    .A2(_10311_),
    .Y(_10312_),
    .B1(net5523));
 sg13g2_a22oi_1 _18696_ (.Y(_10313_),
    .B1(net5370),
    .B2(\atari2600.ram[75][1] ),
    .A2(net5417),
    .A1(\atari2600.ram[72][1] ));
 sg13g2_a22oi_1 _18697_ (.Y(_10314_),
    .B1(net5323),
    .B2(\atari2600.ram[74][1] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][1] ));
 sg13g2_a21oi_1 _18698_ (.A1(_10313_),
    .A2(_10314_),
    .Y(_10315_),
    .B1(net5485));
 sg13g2_nor4_1 _18699_ (.A(_10306_),
    .B(_10309_),
    .C(_10312_),
    .D(_10315_),
    .Y(_10316_));
 sg13g2_nor2_1 _18700_ (.A(net5271),
    .B(_10316_),
    .Y(_10317_));
 sg13g2_o21ai_1 _18701_ (.B1(net5545),
    .Y(_10318_),
    .A1(net5266),
    .A2(_10303_));
 sg13g2_nor3_2 _18702_ (.A(_10290_),
    .B(_10317_),
    .C(_10318_),
    .Y(_10319_));
 sg13g2_a22oi_1 _18703_ (.Y(_10320_),
    .B1(net5301),
    .B2(\atari2600.ram[50][1] ),
    .A2(net5441),
    .A1(\atari2600.ram[49][1] ));
 sg13g2_a221oi_1 _18704_ (.B2(\atari2600.ram[51][1] ),
    .C1(net5281),
    .B1(net5346),
    .A1(\atari2600.ram[48][1] ),
    .Y(_10321_),
    .A2(net5392));
 sg13g2_a21oi_1 _18705_ (.A1(_10320_),
    .A2(_10321_),
    .Y(_10322_),
    .B1(_09293_));
 sg13g2_a22oi_1 _18706_ (.Y(_10323_),
    .B1(net5395),
    .B2(\atari2600.ram[56][1] ),
    .A2(net5444),
    .A1(\atari2600.ram[57][1] ));
 sg13g2_a22oi_1 _18707_ (.Y(_10324_),
    .B1(net5304),
    .B2(\atari2600.ram[58][1] ),
    .A2(net5350),
    .A1(\atari2600.ram[59][1] ));
 sg13g2_a21oi_2 _18708_ (.B1(net5480),
    .Y(_10325_),
    .A2(_10324_),
    .A1(_10323_));
 sg13g2_a22oi_1 _18709_ (.Y(_10326_),
    .B1(net5350),
    .B2(\atari2600.ram[63][1] ),
    .A2(net5395),
    .A1(\atari2600.ram[60][1] ));
 sg13g2_a22oi_1 _18710_ (.Y(_10327_),
    .B1(net5300),
    .B2(\atari2600.ram[62][1] ),
    .A2(net5440),
    .A1(\atari2600.ram[61][1] ));
 sg13g2_a21oi_1 _18711_ (.A1(_10326_),
    .A2(_10327_),
    .Y(_10328_),
    .B1(net5489));
 sg13g2_a22oi_1 _18712_ (.Y(_10329_),
    .B1(net5347),
    .B2(\atari2600.ram[55][1] ),
    .A2(net5392),
    .A1(\atari2600.ram[52][1] ));
 sg13g2_a22oi_1 _18713_ (.Y(_10330_),
    .B1(net5300),
    .B2(\atari2600.ram[54][1] ),
    .A2(net5440),
    .A1(\atari2600.ram[53][1] ));
 sg13g2_a21oi_1 _18714_ (.A1(_10329_),
    .A2(_10330_),
    .Y(_10331_),
    .B1(net5518));
 sg13g2_nor4_2 _18715_ (.A(_10322_),
    .B(_10325_),
    .C(_10328_),
    .Y(_10332_),
    .D(_10331_));
 sg13g2_a22oi_1 _18716_ (.Y(_10333_),
    .B1(net5340),
    .B2(\atari2600.ram[47][1] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][1] ));
 sg13g2_a22oi_1 _18717_ (.Y(_10334_),
    .B1(net5293),
    .B2(\atari2600.ram[46][1] ),
    .A2(net5433),
    .A1(\atari2600.ram[45][1] ));
 sg13g2_a21oi_1 _18718_ (.A1(_10333_),
    .A2(_10334_),
    .Y(_10335_),
    .B1(net5490));
 sg13g2_nand2b_1 _18719_ (.Y(_10336_),
    .B(net5279),
    .A_N(_10335_));
 sg13g2_a22oi_1 _18720_ (.Y(_10337_),
    .B1(net5341),
    .B2(\atari2600.ram[35][1] ),
    .A2(net5386),
    .A1(\atari2600.ram[32][1] ));
 sg13g2_a22oi_1 _18721_ (.Y(_10338_),
    .B1(net5294),
    .B2(\atari2600.ram[34][1] ),
    .A2(net5434),
    .A1(\atari2600.ram[33][1] ));
 sg13g2_a21oi_1 _18722_ (.A1(_10337_),
    .A2(_10338_),
    .Y(_10339_),
    .B1(net5501));
 sg13g2_a22oi_1 _18723_ (.Y(_10340_),
    .B1(net5389),
    .B2(\atari2600.ram[40][1] ),
    .A2(net5437),
    .A1(\atari2600.ram[41][1] ));
 sg13g2_a22oi_1 _18724_ (.Y(_10341_),
    .B1(net5297),
    .B2(\atari2600.ram[42][1] ),
    .A2(net5344),
    .A1(\atari2600.ram[43][1] ));
 sg13g2_a21oi_1 _18725_ (.A1(_10340_),
    .A2(_10341_),
    .Y(_10342_),
    .B1(net5477));
 sg13g2_a22oi_1 _18726_ (.Y(_10343_),
    .B1(net5341),
    .B2(\atari2600.ram[39][1] ),
    .A2(net5386),
    .A1(\atari2600.ram[36][1] ));
 sg13g2_a22oi_1 _18727_ (.Y(_10344_),
    .B1(net5293),
    .B2(\atari2600.ram[38][1] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][1] ));
 sg13g2_a21oi_2 _18728_ (.B1(net5515),
    .Y(_10345_),
    .A2(_10344_),
    .A1(_10343_));
 sg13g2_nor4_2 _18729_ (.A(_10336_),
    .B(_10339_),
    .C(_10342_),
    .Y(_10346_),
    .D(_10345_));
 sg13g2_nor3_2 _18730_ (.A(net5568),
    .B(_10332_),
    .C(_10346_),
    .Y(_10347_));
 sg13g2_a22oi_1 _18731_ (.Y(_10348_),
    .B1(net5355),
    .B2(\atari2600.ram[7][1] ),
    .A2(net5399),
    .A1(\atari2600.ram[4][1] ));
 sg13g2_a22oi_1 _18732_ (.Y(_10349_),
    .B1(net5311),
    .B2(\atari2600.ram[6][1] ),
    .A2(net5451),
    .A1(\atari2600.ram[5][1] ));
 sg13g2_a21oi_1 _18733_ (.A1(_10348_),
    .A2(_10349_),
    .Y(_10350_),
    .B1(net5516));
 sg13g2_a22oi_1 _18734_ (.Y(_10351_),
    .B1(net5354),
    .B2(\atari2600.ram[15][1] ),
    .A2(net5399),
    .A1(\atari2600.ram[12][1] ));
 sg13g2_a22oi_1 _18735_ (.Y(_10352_),
    .B1(net5306),
    .B2(\atari2600.ram[14][1] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][1] ));
 sg13g2_a21oi_1 _18736_ (.A1(_10351_),
    .A2(_10352_),
    .Y(_10353_),
    .B1(net5491));
 sg13g2_a22oi_1 _18737_ (.Y(_10354_),
    .B1(net5353),
    .B2(\atari2600.ram[3][1] ),
    .A2(net5400),
    .A1(\atari2600.ram[0][1] ));
 sg13g2_a22oi_1 _18738_ (.Y(_10355_),
    .B1(net5307),
    .B2(\atari2600.ram[2][1] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][1] ));
 sg13g2_a21oi_1 _18739_ (.A1(_10354_),
    .A2(_10355_),
    .Y(_10356_),
    .B1(net5507));
 sg13g2_a22oi_1 _18740_ (.Y(_10357_),
    .B1(net5345),
    .B2(\atari2600.ram[11][1] ),
    .A2(net5390),
    .A1(\atari2600.ram[8][1] ));
 sg13g2_a22oi_1 _18741_ (.Y(_10358_),
    .B1(net5297),
    .B2(\atari2600.ram[10][1] ),
    .A2(net5436),
    .A1(\atari2600.ram[9][1] ));
 sg13g2_a21oi_2 _18742_ (.B1(net5478),
    .Y(_10359_),
    .A2(_10358_),
    .A1(_10357_));
 sg13g2_nor4_1 _18743_ (.A(_10350_),
    .B(_10353_),
    .C(_10356_),
    .D(_10359_),
    .Y(_10360_));
 sg13g2_nor2_1 _18744_ (.A(net5270),
    .B(_10360_),
    .Y(_10361_));
 sg13g2_a22oi_1 _18745_ (.Y(_10362_),
    .B1(net5356),
    .B2(\atari2600.ram[23][1] ),
    .A2(net5402),
    .A1(\atari2600.ram[20][1] ));
 sg13g2_a22oi_1 _18746_ (.Y(_10363_),
    .B1(net5309),
    .B2(\atari2600.ram[22][1] ),
    .A2(net5449),
    .A1(\atari2600.ram[21][1] ));
 sg13g2_a21oi_1 _18747_ (.A1(_10362_),
    .A2(_10363_),
    .Y(_10364_),
    .B1(net5517));
 sg13g2_a22oi_1 _18748_ (.Y(_10365_),
    .B1(net5371),
    .B2(\atari2600.ram[27][1] ),
    .A2(net5419),
    .A1(\atari2600.ram[24][1] ));
 sg13g2_a22oi_1 _18749_ (.Y(_10366_),
    .B1(net5326),
    .B2(\atari2600.ram[26][1] ),
    .A2(net5465),
    .A1(\atari2600.ram[25][1] ));
 sg13g2_a21oi_1 _18750_ (.A1(_10365_),
    .A2(_10366_),
    .Y(_10367_),
    .B1(net5487));
 sg13g2_a22oi_1 _18751_ (.Y(_10368_),
    .B1(net5356),
    .B2(\atari2600.ram[19][1] ),
    .A2(net5403),
    .A1(\atari2600.ram[16][1] ));
 sg13g2_a22oi_1 _18752_ (.Y(_10369_),
    .B1(net5310),
    .B2(\atari2600.ram[18][1] ),
    .A2(net5450),
    .A1(\atari2600.ram[17][1] ));
 sg13g2_a21oi_1 _18753_ (.A1(_10368_),
    .A2(_10369_),
    .Y(_10370_),
    .B1(net5505));
 sg13g2_a22oi_1 _18754_ (.Y(_10371_),
    .B1(net5374),
    .B2(\atari2600.ram[31][1] ),
    .A2(net5421),
    .A1(\atari2600.ram[28][1] ));
 sg13g2_a22oi_1 _18755_ (.Y(_10372_),
    .B1(net5330),
    .B2(\atari2600.ram[30][1] ),
    .A2(net5469),
    .A1(\atari2600.ram[29][1] ));
 sg13g2_a21oi_2 _18756_ (.B1(net5492),
    .Y(_10373_),
    .A2(_10372_),
    .A1(_10371_));
 sg13g2_nor4_2 _18757_ (.A(_10364_),
    .B(_10367_),
    .C(_10370_),
    .Y(_10374_),
    .D(_10373_));
 sg13g2_o21ai_1 _18758_ (.B1(net5542),
    .Y(_10375_),
    .A1(net5265),
    .A2(_10374_));
 sg13g2_nor3_1 _18759_ (.A(_10347_),
    .B(_10361_),
    .C(_10375_),
    .Y(_10376_));
 sg13g2_nor2_1 _18760_ (.A(_10319_),
    .B(_10376_),
    .Y(_00002_));
 sg13g2_a22oi_1 _18761_ (.Y(_10377_),
    .B1(net5298),
    .B2(\atari2600.ram[50][2] ),
    .A2(net5438),
    .A1(\atari2600.ram[49][2] ));
 sg13g2_a221oi_1 _18762_ (.B2(\atari2600.ram[51][2] ),
    .C1(net5279),
    .B1(net5349),
    .A1(\atari2600.ram[48][2] ),
    .Y(_10378_),
    .A2(net5394));
 sg13g2_a21oi_1 _18763_ (.A1(_10377_),
    .A2(_10378_),
    .Y(_10379_),
    .B1(_09293_));
 sg13g2_a22oi_1 _18764_ (.Y(_10380_),
    .B1(net5351),
    .B2(\atari2600.ram[59][2] ),
    .A2(net5396),
    .A1(\atari2600.ram[56][2] ));
 sg13g2_a22oi_1 _18765_ (.Y(_10381_),
    .B1(net5304),
    .B2(\atari2600.ram[58][2] ),
    .A2(net5444),
    .A1(\atari2600.ram[57][2] ));
 sg13g2_a21oi_2 _18766_ (.B1(net5480),
    .Y(_10382_),
    .A2(_10381_),
    .A1(_10380_));
 sg13g2_a22oi_1 _18767_ (.Y(_10383_),
    .B1(net5392),
    .B2(\atari2600.ram[52][2] ),
    .A2(net5440),
    .A1(\atari2600.ram[53][2] ));
 sg13g2_a22oi_1 _18768_ (.Y(_10384_),
    .B1(net5300),
    .B2(\atari2600.ram[54][2] ),
    .A2(net5347),
    .A1(\atari2600.ram[55][2] ));
 sg13g2_a21oi_2 _18769_ (.B1(net5518),
    .Y(_10385_),
    .A2(_10384_),
    .A1(_10383_));
 sg13g2_a22oi_1 _18770_ (.Y(_10386_),
    .B1(net5350),
    .B2(\atari2600.ram[63][2] ),
    .A2(net5395),
    .A1(\atari2600.ram[60][2] ));
 sg13g2_a22oi_1 _18771_ (.Y(_10387_),
    .B1(net5301),
    .B2(\atari2600.ram[62][2] ),
    .A2(net5441),
    .A1(\atari2600.ram[61][2] ));
 sg13g2_a21oi_1 _18772_ (.A1(_10386_),
    .A2(_10387_),
    .Y(_10388_),
    .B1(net5489));
 sg13g2_nor4_2 _18773_ (.A(_10379_),
    .B(_10382_),
    .C(_10385_),
    .Y(_10389_),
    .D(_10388_));
 sg13g2_a22oi_1 _18774_ (.Y(_10390_),
    .B1(net5342),
    .B2(\atari2600.ram[47][2] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][2] ));
 sg13g2_a22oi_1 _18775_ (.Y(_10391_),
    .B1(net5295),
    .B2(\atari2600.ram[46][2] ),
    .A2(net5435),
    .A1(\atari2600.ram[45][2] ));
 sg13g2_a21oi_2 _18776_ (.B1(net5490),
    .Y(_10392_),
    .A2(_10391_),
    .A1(_10390_));
 sg13g2_nand2b_1 _18777_ (.Y(_10393_),
    .B(net5279),
    .A_N(_10392_));
 sg13g2_a22oi_1 _18778_ (.Y(_10394_),
    .B1(net5389),
    .B2(\atari2600.ram[40][2] ),
    .A2(net5437),
    .A1(\atari2600.ram[41][2] ));
 sg13g2_a22oi_1 _18779_ (.Y(_10395_),
    .B1(net5297),
    .B2(\atari2600.ram[42][2] ),
    .A2(net5344),
    .A1(\atari2600.ram[43][2] ));
 sg13g2_a21oi_1 _18780_ (.A1(_10394_),
    .A2(_10395_),
    .Y(_10396_),
    .B1(net5477));
 sg13g2_a22oi_1 _18781_ (.Y(_10397_),
    .B1(net5340),
    .B2(\atari2600.ram[39][2] ),
    .A2(net5385),
    .A1(\atari2600.ram[36][2] ));
 sg13g2_a22oi_1 _18782_ (.Y(_10398_),
    .B1(net5293),
    .B2(\atari2600.ram[38][2] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][2] ));
 sg13g2_a21oi_2 _18783_ (.B1(net5515),
    .Y(_10399_),
    .A2(_10398_),
    .A1(_10397_));
 sg13g2_a22oi_1 _18784_ (.Y(_10400_),
    .B1(net5341),
    .B2(\atari2600.ram[35][2] ),
    .A2(net5386),
    .A1(\atari2600.ram[32][2] ));
 sg13g2_a22oi_1 _18785_ (.Y(_10401_),
    .B1(net5294),
    .B2(\atari2600.ram[34][2] ),
    .A2(net5434),
    .A1(\atari2600.ram[33][2] ));
 sg13g2_a21oi_1 _18786_ (.A1(_10400_),
    .A2(_10401_),
    .Y(_10402_),
    .B1(net5501));
 sg13g2_nor4_2 _18787_ (.A(_10393_),
    .B(_10396_),
    .C(_10399_),
    .Y(_10403_),
    .D(_10402_));
 sg13g2_nor3_2 _18788_ (.A(net5568),
    .B(_10389_),
    .C(_10403_),
    .Y(_10404_));
 sg13g2_a22oi_1 _18789_ (.Y(_10405_),
    .B1(net5373),
    .B2(\atari2600.ram[31][2] ),
    .A2(net5422),
    .A1(\atari2600.ram[28][2] ));
 sg13g2_a22oi_1 _18790_ (.Y(_10406_),
    .B1(net5328),
    .B2(\atari2600.ram[30][2] ),
    .A2(net5467),
    .A1(\atari2600.ram[29][2] ));
 sg13g2_a21oi_2 _18791_ (.B1(net5498),
    .Y(_10407_),
    .A2(_10406_),
    .A1(_10405_));
 sg13g2_a22oi_1 _18792_ (.Y(_10408_),
    .B1(net5372),
    .B2(\atari2600.ram[27][2] ),
    .A2(net5420),
    .A1(\atari2600.ram[24][2] ));
 sg13g2_a22oi_1 _18793_ (.Y(_10409_),
    .B1(net5327),
    .B2(\atari2600.ram[26][2] ),
    .A2(net5466),
    .A1(\atari2600.ram[25][2] ));
 sg13g2_a21oi_1 _18794_ (.A1(_10408_),
    .A2(_10409_),
    .Y(_10410_),
    .B1(net5484));
 sg13g2_a22oi_1 _18795_ (.Y(_10411_),
    .B1(net5356),
    .B2(\atari2600.ram[19][2] ),
    .A2(net5402),
    .A1(\atari2600.ram[16][2] ));
 sg13g2_a22oi_1 _18796_ (.Y(_10412_),
    .B1(net5310),
    .B2(\atari2600.ram[18][2] ),
    .A2(net5449),
    .A1(\atari2600.ram[17][2] ));
 sg13g2_a21oi_1 _18797_ (.A1(_10411_),
    .A2(_10412_),
    .Y(_10413_),
    .B1(net5504));
 sg13g2_a22oi_1 _18798_ (.Y(_10414_),
    .B1(net5372),
    .B2(\atari2600.ram[23][2] ),
    .A2(net5420),
    .A1(\atari2600.ram[20][2] ));
 sg13g2_a22oi_1 _18799_ (.Y(_10415_),
    .B1(net5327),
    .B2(\atari2600.ram[22][2] ),
    .A2(net5465),
    .A1(\atari2600.ram[21][2] ));
 sg13g2_a21oi_1 _18800_ (.A1(_10414_),
    .A2(_10415_),
    .Y(_10416_),
    .B1(net5517));
 sg13g2_nor4_2 _18801_ (.A(_10407_),
    .B(_10410_),
    .C(_10413_),
    .Y(_10417_),
    .D(_10416_));
 sg13g2_a22oi_1 _18802_ (.Y(_10418_),
    .B1(net5358),
    .B2(\atari2600.ram[7][2] ),
    .A2(net5401),
    .A1(\atari2600.ram[4][2] ));
 sg13g2_a22oi_1 _18803_ (.Y(_10419_),
    .B1(net5308),
    .B2(\atari2600.ram[6][2] ),
    .A2(net5448),
    .A1(\atari2600.ram[5][2] ));
 sg13g2_a21oi_1 _18804_ (.A1(_10418_),
    .A2(_10419_),
    .Y(_10420_),
    .B1(net5516));
 sg13g2_a22oi_1 _18805_ (.Y(_10421_),
    .B1(net5353),
    .B2(\atari2600.ram[3][2] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][2] ));
 sg13g2_a22oi_1 _18806_ (.Y(_10422_),
    .B1(net5307),
    .B2(\atari2600.ram[2][2] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][2] ));
 sg13g2_a21oi_1 _18807_ (.A1(_10421_),
    .A2(_10422_),
    .Y(_10423_),
    .B1(net5503));
 sg13g2_a22oi_1 _18808_ (.Y(_10424_),
    .B1(net5357),
    .B2(\atari2600.ram[15][2] ),
    .A2(net5404),
    .A1(\atari2600.ram[12][2] ));
 sg13g2_a22oi_1 _18809_ (.Y(_10425_),
    .B1(net5306),
    .B2(\atari2600.ram[14][2] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][2] ));
 sg13g2_a21oi_1 _18810_ (.A1(_10424_),
    .A2(_10425_),
    .Y(_10426_),
    .B1(net5492));
 sg13g2_a22oi_1 _18811_ (.Y(_10427_),
    .B1(net5349),
    .B2(\atari2600.ram[11][2] ),
    .A2(net5394),
    .A1(\atari2600.ram[8][2] ));
 sg13g2_a22oi_1 _18812_ (.Y(_10428_),
    .B1(net5296),
    .B2(\atari2600.ram[10][2] ),
    .A2(net5436),
    .A1(\atari2600.ram[9][2] ));
 sg13g2_a21oi_2 _18813_ (.B1(net5478),
    .Y(_10429_),
    .A2(_10428_),
    .A1(_10427_));
 sg13g2_nor4_1 _18814_ (.A(_10420_),
    .B(_10423_),
    .C(_10426_),
    .D(_10429_),
    .Y(_10430_));
 sg13g2_nor2_1 _18815_ (.A(net5270),
    .B(_10430_),
    .Y(_10431_));
 sg13g2_o21ai_1 _18816_ (.B1(net5542),
    .Y(_10432_),
    .A1(net5264),
    .A2(_10417_));
 sg13g2_nor3_1 _18817_ (.A(_10404_),
    .B(_10431_),
    .C(_10432_),
    .Y(_10433_));
 sg13g2_a22oi_1 _18818_ (.Y(_10434_),
    .B1(net5366),
    .B2(\atari2600.ram[103][2] ),
    .A2(net5413),
    .A1(\atari2600.ram[100][2] ));
 sg13g2_a22oi_1 _18819_ (.Y(_10435_),
    .B1(net5322),
    .B2(\atari2600.ram[102][2] ),
    .A2(net5461),
    .A1(\atari2600.ram[101][2] ));
 sg13g2_a21oi_1 _18820_ (.A1(_10434_),
    .A2(_10435_),
    .Y(_10436_),
    .B1(net5521));
 sg13g2_a22oi_1 _18821_ (.Y(_10437_),
    .B1(net5369),
    .B2(\atari2600.ram[99][2] ),
    .A2(net5416),
    .A1(\atari2600.ram[96][2] ));
 sg13g2_a22oi_1 _18822_ (.Y(_10438_),
    .B1(net5322),
    .B2(\atari2600.ram[98][2] ),
    .A2(net5461),
    .A1(\atari2600.ram[97][2] ));
 sg13g2_a21oi_1 _18823_ (.A1(_10437_),
    .A2(_10438_),
    .Y(_10439_),
    .B1(net5511));
 sg13g2_a22oi_1 _18824_ (.Y(_10440_),
    .B1(net5363),
    .B2(\atari2600.ram[107][2] ),
    .A2(net5409),
    .A1(\atari2600.ram[104][2] ));
 sg13g2_a22oi_1 _18825_ (.Y(_10441_),
    .B1(net5316),
    .B2(\atari2600.ram[106][2] ),
    .A2(net5455),
    .A1(\atari2600.ram[105][2] ));
 sg13g2_a21oi_1 _18826_ (.A1(_10440_),
    .A2(_10441_),
    .Y(_10442_),
    .B1(net5483));
 sg13g2_a22oi_1 _18827_ (.Y(_10443_),
    .B1(net5365),
    .B2(\atari2600.ram[111][2] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][2] ));
 sg13g2_a22oi_1 _18828_ (.Y(_10444_),
    .B1(net5319),
    .B2(\atari2600.ram[110][2] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][2] ));
 sg13g2_a21oi_2 _18829_ (.B1(net5495),
    .Y(_10445_),
    .A2(_10444_),
    .A1(_10443_));
 sg13g2_nor4_1 _18830_ (.A(_10436_),
    .B(_10439_),
    .C(_10442_),
    .D(_10445_),
    .Y(_10446_));
 sg13g2_a22oi_1 _18831_ (.Y(_10447_),
    .B1(net5381),
    .B2(\atari2600.ram[91][2] ),
    .A2(net5429),
    .A1(\atari2600.ram[88][2] ));
 sg13g2_a22oi_1 _18832_ (.Y(_10448_),
    .B1(net5334),
    .B2(\atari2600.ram[90][2] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][2] ));
 sg13g2_a22oi_1 _18833_ (.Y(_10449_),
    .B1(net5372),
    .B2(\atari2600.ram[95][2] ),
    .A2(net5420),
    .A1(\atari2600.ram[92][2] ));
 sg13g2_a22oi_1 _18834_ (.Y(_10450_),
    .B1(net5329),
    .B2(\atari2600.ram[94][2] ),
    .A2(net5468),
    .A1(\atari2600.ram[93][2] ));
 sg13g2_a21oi_1 _18835_ (.A1(_10449_),
    .A2(_10450_),
    .Y(_10451_),
    .B1(net5498));
 sg13g2_a22oi_1 _18836_ (.Y(_10452_),
    .B1(net5374),
    .B2(\atari2600.ram[83][2] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][2] ));
 sg13g2_a22oi_1 _18837_ (.Y(_10453_),
    .B1(net5330),
    .B2(\atari2600.ram[82][2] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][2] ));
 sg13g2_a21oi_1 _18838_ (.A1(_10452_),
    .A2(_10453_),
    .Y(_10454_),
    .B1(net5508));
 sg13g2_a22oi_1 _18839_ (.Y(_10455_),
    .B1(net5381),
    .B2(\atari2600.ram[87][2] ),
    .A2(net5429),
    .A1(\atari2600.ram[84][2] ));
 sg13g2_a22oi_1 _18840_ (.Y(_10456_),
    .B1(net5335),
    .B2(\atari2600.ram[86][2] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][2] ));
 sg13g2_a21oi_1 _18841_ (.A1(_10455_),
    .A2(_10456_),
    .Y(_10457_),
    .B1(net5523));
 sg13g2_a22oi_1 _18842_ (.Y(_10458_),
    .B1(net5370),
    .B2(\atari2600.ram[79][2] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][2] ));
 sg13g2_a22oi_1 _18843_ (.Y(_10459_),
    .B1(net5320),
    .B2(\atari2600.ram[78][2] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][2] ));
 sg13g2_a21oi_2 _18844_ (.B1(net5496),
    .Y(_10460_),
    .A2(_10459_),
    .A1(_10458_));
 sg13g2_a22oi_1 _18845_ (.Y(_10461_),
    .B1(net5368),
    .B2(\atari2600.ram[75][2] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][2] ));
 sg13g2_a22oi_1 _18846_ (.Y(_10462_),
    .B1(net5323),
    .B2(\atari2600.ram[74][2] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][2] ));
 sg13g2_a21oi_1 _18847_ (.A1(_10461_),
    .A2(_10462_),
    .Y(_10463_),
    .B1(net5485));
 sg13g2_a22oi_1 _18848_ (.Y(_10464_),
    .B1(net5377),
    .B2(\atari2600.ram[71][2] ),
    .A2(net5427),
    .A1(\atari2600.ram[68][2] ));
 sg13g2_a22oi_1 _18849_ (.Y(_10465_),
    .B1(net5332),
    .B2(\atari2600.ram[70][2] ),
    .A2(net5471),
    .A1(\atari2600.ram[69][2] ));
 sg13g2_a21oi_2 _18850_ (.B1(net5523),
    .Y(_10466_),
    .A2(_10465_),
    .A1(_10464_));
 sg13g2_a22oi_1 _18851_ (.Y(_10467_),
    .B1(net5370),
    .B2(\atari2600.ram[67][2] ),
    .A2(net5417),
    .A1(\atari2600.ram[64][2] ));
 sg13g2_a22oi_1 _18852_ (.Y(_10468_),
    .B1(net5324),
    .B2(\atari2600.ram[66][2] ),
    .A2(net5463),
    .A1(\atari2600.ram[65][2] ));
 sg13g2_a21oi_1 _18853_ (.A1(_10467_),
    .A2(_10468_),
    .Y(_10469_),
    .B1(net5511));
 sg13g2_nor4_2 _18854_ (.A(_10460_),
    .B(_10463_),
    .C(_10466_),
    .Y(_10470_),
    .D(_10469_));
 sg13g2_a22oi_1 _18855_ (.Y(_10471_),
    .B1(net5362),
    .B2(\atari2600.ram[115][2] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][2] ));
 sg13g2_a22oi_1 _18856_ (.Y(_10472_),
    .B1(net5317),
    .B2(\atari2600.ram[114][2] ),
    .A2(net5456),
    .A1(\atari2600.ram[113][2] ));
 sg13g2_a21oi_1 _18857_ (.A1(_10471_),
    .A2(_10472_),
    .Y(_10473_),
    .B1(net5510));
 sg13g2_a22oi_1 _18858_ (.Y(_10474_),
    .B1(net5362),
    .B2(\atari2600.ram[123][2] ),
    .A2(net5410),
    .A1(\atari2600.ram[120][2] ));
 sg13g2_a22oi_1 _18859_ (.Y(_10475_),
    .B1(net5318),
    .B2(\atari2600.ram[122][2] ),
    .A2(net5457),
    .A1(\atari2600.ram[121][2] ));
 sg13g2_a21oi_1 _18860_ (.A1(_10474_),
    .A2(_10475_),
    .Y(_10476_),
    .B1(net5482));
 sg13g2_a22oi_1 _18861_ (.Y(_10477_),
    .B1(net5359),
    .B2(\atari2600.ram[127][2] ),
    .A2(net5406),
    .A1(\atari2600.ram[124][2] ));
 sg13g2_a22oi_1 _18862_ (.Y(_10478_),
    .B1(net5314),
    .B2(\atari2600.ram[126][2] ),
    .A2(net5453),
    .A1(\atari2600.ram[125][2] ));
 sg13g2_a21oi_2 _18863_ (.B1(net5494),
    .Y(_10479_),
    .A2(_10478_),
    .A1(_10477_));
 sg13g2_a22oi_1 _18864_ (.Y(_10480_),
    .B1(net5361),
    .B2(\atari2600.ram[119][2] ),
    .A2(net5409),
    .A1(\atari2600.ram[116][2] ));
 sg13g2_a22oi_1 _18865_ (.Y(_10481_),
    .B1(net5315),
    .B2(\atari2600.ram[118][2] ),
    .A2(net5454),
    .A1(\atari2600.ram[117][2] ));
 sg13g2_a21oi_1 _18866_ (.A1(_10480_),
    .A2(_10481_),
    .Y(_10482_),
    .B1(net5520));
 sg13g2_nor4_2 _18867_ (.A(_10473_),
    .B(_10476_),
    .C(_10479_),
    .Y(_10483_),
    .D(_10482_));
 sg13g2_a21oi_1 _18868_ (.A1(_10447_),
    .A2(_10448_),
    .Y(_10484_),
    .B1(net5484));
 sg13g2_nor4_2 _18869_ (.A(_10451_),
    .B(_10454_),
    .C(_10457_),
    .Y(_10485_),
    .D(_10484_));
 sg13g2_mux4_1 _18870_ (.S0(net5571),
    .A0(_10446_),
    .A1(_10470_),
    .A2(_10483_),
    .A3(_10485_),
    .S1(net5276),
    .X(_10486_));
 sg13g2_a21oi_1 _18871_ (.A1(net5544),
    .A2(_10486_),
    .Y(_00003_),
    .B1(_10433_));
 sg13g2_a22oi_1 _18872_ (.Y(_10487_),
    .B1(net5394),
    .B2(\atari2600.ram[56][3] ),
    .A2(net5443),
    .A1(\atari2600.ram[57][3] ));
 sg13g2_a22oi_1 _18873_ (.Y(_10488_),
    .B1(net5303),
    .B2(\atari2600.ram[58][3] ),
    .A2(net5349),
    .A1(\atari2600.ram[59][3] ));
 sg13g2_a21oi_1 _18874_ (.A1(_10487_),
    .A2(_10488_),
    .Y(_10489_),
    .B1(net5480));
 sg13g2_a22oi_1 _18875_ (.Y(_10490_),
    .B1(net5346),
    .B2(\atari2600.ram[55][3] ),
    .A2(net5391),
    .A1(\atari2600.ram[52][3] ));
 sg13g2_a22oi_1 _18876_ (.Y(_10491_),
    .B1(net5298),
    .B2(\atari2600.ram[54][3] ),
    .A2(net5438),
    .A1(\atari2600.ram[53][3] ));
 sg13g2_a21oi_1 _18877_ (.A1(_10490_),
    .A2(_10491_),
    .Y(_10492_),
    .B1(net5518));
 sg13g2_a22oi_1 _18878_ (.Y(_10493_),
    .B1(net5347),
    .B2(\atari2600.ram[63][3] ),
    .A2(net5392),
    .A1(\atari2600.ram[60][3] ));
 sg13g2_a22oi_1 _18879_ (.Y(_10494_),
    .B1(net5300),
    .B2(\atari2600.ram[62][3] ),
    .A2(net5440),
    .A1(\atari2600.ram[61][3] ));
 sg13g2_a21oi_1 _18880_ (.A1(_10493_),
    .A2(_10494_),
    .Y(_10495_),
    .B1(net5488));
 sg13g2_a22oi_1 _18881_ (.Y(_10496_),
    .B1(net5342),
    .B2(\atari2600.ram[51][3] ),
    .A2(net5393),
    .A1(\atari2600.ram[48][3] ));
 sg13g2_a22oi_1 _18882_ (.Y(_10497_),
    .B1(net5299),
    .B2(\atari2600.ram[50][3] ),
    .A2(net5439),
    .A1(\atari2600.ram[49][3] ));
 sg13g2_a21o_1 _18883_ (.A2(_10497_),
    .A1(_10496_),
    .B1(net5502),
    .X(_10498_));
 sg13g2_nor4_1 _18884_ (.A(net5280),
    .B(_10489_),
    .C(_10492_),
    .D(_10495_),
    .Y(_10499_));
 sg13g2_a22oi_1 _18885_ (.Y(_10500_),
    .B1(net5385),
    .B2(\atari2600.ram[36][3] ),
    .A2(net5434),
    .A1(\atari2600.ram[37][3] ));
 sg13g2_a22oi_1 _18886_ (.Y(_10501_),
    .B1(net5294),
    .B2(\atari2600.ram[38][3] ),
    .A2(net5341),
    .A1(\atari2600.ram[39][3] ));
 sg13g2_a21oi_1 _18887_ (.A1(_10500_),
    .A2(_10501_),
    .Y(_10502_),
    .B1(net5515));
 sg13g2_a22oi_1 _18888_ (.Y(_10503_),
    .B1(net5343),
    .B2(\atari2600.ram[35][3] ),
    .A2(net5388),
    .A1(\atari2600.ram[32][3] ));
 sg13g2_a22oi_1 _18889_ (.Y(_10504_),
    .B1(net5295),
    .B2(\atari2600.ram[34][3] ),
    .A2(net5435),
    .A1(\atari2600.ram[33][3] ));
 sg13g2_a21oi_1 _18890_ (.A1(_10503_),
    .A2(_10504_),
    .Y(_10505_),
    .B1(net5502));
 sg13g2_a22oi_1 _18891_ (.Y(_10506_),
    .B1(net5342),
    .B2(\atari2600.ram[47][3] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][3] ));
 sg13g2_a22oi_1 _18892_ (.Y(_10507_),
    .B1(net5295),
    .B2(\atari2600.ram[46][3] ),
    .A2(net5435),
    .A1(\atari2600.ram[45][3] ));
 sg13g2_a21oi_1 _18893_ (.A1(_10506_),
    .A2(_10507_),
    .Y(_10508_),
    .B1(net5490));
 sg13g2_a22oi_1 _18894_ (.Y(_10509_),
    .B1(net5345),
    .B2(\atari2600.ram[43][3] ),
    .A2(net5390),
    .A1(\atari2600.ram[40][3] ));
 sg13g2_a22oi_1 _18895_ (.Y(_10510_),
    .B1(net5296),
    .B2(\atari2600.ram[42][3] ),
    .A2(net5436),
    .A1(\atari2600.ram[41][3] ));
 sg13g2_a21oi_2 _18896_ (.B1(net5477),
    .Y(_10511_),
    .A2(_10510_),
    .A1(_10509_));
 sg13g2_nor2_1 _18897_ (.A(net5275),
    .B(_10505_),
    .Y(_10512_));
 sg13g2_nor3_2 _18898_ (.A(_10502_),
    .B(_10508_),
    .C(_10511_),
    .Y(_10513_));
 sg13g2_a221oi_1 _18899_ (.B2(_10513_),
    .C1(net5568),
    .B1(_10512_),
    .A1(_10498_),
    .Y(_10514_),
    .A2(_10499_));
 sg13g2_a22oi_1 _18900_ (.Y(_10515_),
    .B1(net5353),
    .B2(\atari2600.ram[11][3] ),
    .A2(net5398),
    .A1(\atari2600.ram[8][3] ));
 sg13g2_a22oi_1 _18901_ (.Y(_10516_),
    .B1(net5307),
    .B2(\atari2600.ram[10][3] ),
    .A2(net5447),
    .A1(\atari2600.ram[9][3] ));
 sg13g2_a21oi_2 _18902_ (.B1(net5478),
    .Y(_10517_),
    .A2(_10516_),
    .A1(_10515_));
 sg13g2_a22oi_1 _18903_ (.Y(_10518_),
    .B1(net5355),
    .B2(\atari2600.ram[7][3] ),
    .A2(net5401),
    .A1(\atari2600.ram[4][3] ));
 sg13g2_a22oi_1 _18904_ (.Y(_10519_),
    .B1(net5308),
    .B2(\atari2600.ram[6][3] ),
    .A2(net5448),
    .A1(\atari2600.ram[5][3] ));
 sg13g2_a21oi_1 _18905_ (.A1(_10518_),
    .A2(_10519_),
    .Y(_10520_),
    .B1(net5516));
 sg13g2_a22oi_1 _18906_ (.Y(_10521_),
    .B1(net5354),
    .B2(\atari2600.ram[3][3] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][3] ));
 sg13g2_a22oi_1 _18907_ (.Y(_10522_),
    .B1(net5307),
    .B2(\atari2600.ram[2][3] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][3] ));
 sg13g2_a21oi_1 _18908_ (.A1(_10521_),
    .A2(_10522_),
    .Y(_10523_),
    .B1(net5503));
 sg13g2_a22oi_1 _18909_ (.Y(_10524_),
    .B1(net5354),
    .B2(\atari2600.ram[15][3] ),
    .A2(net5400),
    .A1(\atari2600.ram[12][3] ));
 sg13g2_a22oi_1 _18910_ (.Y(_10525_),
    .B1(net5306),
    .B2(\atari2600.ram[14][3] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][3] ));
 sg13g2_a21oi_1 _18911_ (.A1(_10524_),
    .A2(_10525_),
    .Y(_10526_),
    .B1(net5491));
 sg13g2_nor4_2 _18912_ (.A(_10517_),
    .B(_10520_),
    .C(_10523_),
    .Y(_10527_),
    .D(_10526_));
 sg13g2_nor2_1 _18913_ (.A(net5270),
    .B(_10527_),
    .Y(_10528_));
 sg13g2_a22oi_1 _18914_ (.Y(_10529_),
    .B1(net5373),
    .B2(\atari2600.ram[19][3] ),
    .A2(net5421),
    .A1(\atari2600.ram[16][3] ));
 sg13g2_a22oi_1 _18915_ (.Y(_10530_),
    .B1(net5328),
    .B2(\atari2600.ram[18][3] ),
    .A2(net5467),
    .A1(\atari2600.ram[17][3] ));
 sg13g2_a21oi_2 _18916_ (.B1(net5505),
    .Y(_10531_),
    .A2(_10530_),
    .A1(_10529_));
 sg13g2_a22oi_1 _18917_ (.Y(_10532_),
    .B1(net5374),
    .B2(\atari2600.ram[31][3] ),
    .A2(net5421),
    .A1(\atari2600.ram[28][3] ));
 sg13g2_a22oi_1 _18918_ (.Y(_10533_),
    .B1(net5328),
    .B2(\atari2600.ram[30][3] ),
    .A2(net5467),
    .A1(\atari2600.ram[29][3] ));
 sg13g2_a21oi_2 _18919_ (.B1(net5492),
    .Y(_10534_),
    .A2(_10533_),
    .A1(_10532_));
 sg13g2_a22oi_1 _18920_ (.Y(_10535_),
    .B1(net5371),
    .B2(\atari2600.ram[23][3] ),
    .A2(net5419),
    .A1(\atari2600.ram[20][3] ));
 sg13g2_a22oi_1 _18921_ (.Y(_10536_),
    .B1(net5326),
    .B2(\atari2600.ram[22][3] ),
    .A2(net5465),
    .A1(\atari2600.ram[21][3] ));
 sg13g2_a21oi_1 _18922_ (.A1(_10535_),
    .A2(_10536_),
    .Y(_10537_),
    .B1(net5522));
 sg13g2_a22oi_1 _18923_ (.Y(_10538_),
    .B1(net5371),
    .B2(\atari2600.ram[27][3] ),
    .A2(net5419),
    .A1(\atari2600.ram[24][3] ));
 sg13g2_a22oi_1 _18924_ (.Y(_10539_),
    .B1(net5326),
    .B2(\atari2600.ram[26][3] ),
    .A2(net5465),
    .A1(\atari2600.ram[25][3] ));
 sg13g2_a21oi_1 _18925_ (.A1(_10538_),
    .A2(_10539_),
    .Y(_10540_),
    .B1(net5484));
 sg13g2_nor4_2 _18926_ (.A(_10531_),
    .B(_10534_),
    .C(_10537_),
    .Y(_10541_),
    .D(_10540_));
 sg13g2_o21ai_1 _18927_ (.B1(net5542),
    .Y(_10542_),
    .A1(net5264),
    .A2(_10541_));
 sg13g2_nor3_1 _18928_ (.A(_10514_),
    .B(_10528_),
    .C(_10542_),
    .Y(_10543_));
 sg13g2_a22oi_1 _18929_ (.Y(_10544_),
    .B1(net5377),
    .B2(\atari2600.ram[67][3] ),
    .A2(net5425),
    .A1(\atari2600.ram[64][3] ));
 sg13g2_a22oi_1 _18930_ (.Y(_10545_),
    .B1(net5331),
    .B2(\atari2600.ram[66][3] ),
    .A2(net5470),
    .A1(\atari2600.ram[65][3] ));
 sg13g2_a21oi_1 _18931_ (.A1(_10544_),
    .A2(_10545_),
    .Y(_10546_),
    .B1(net5512));
 sg13g2_a22oi_1 _18932_ (.Y(_10547_),
    .B1(net5365),
    .B2(\atari2600.ram[79][3] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][3] ));
 sg13g2_a22oi_1 _18933_ (.Y(_10548_),
    .B1(net5320),
    .B2(\atari2600.ram[78][3] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][3] ));
 sg13g2_a21oi_2 _18934_ (.B1(net5496),
    .Y(_10549_),
    .A2(_10548_),
    .A1(_10547_));
 sg13g2_a22oi_1 _18935_ (.Y(_10550_),
    .B1(net5377),
    .B2(\atari2600.ram[71][3] ),
    .A2(net5425),
    .A1(\atari2600.ram[68][3] ));
 sg13g2_a22oi_1 _18936_ (.Y(_10551_),
    .B1(net5332),
    .B2(\atari2600.ram[70][3] ),
    .A2(net5471),
    .A1(\atari2600.ram[69][3] ));
 sg13g2_a21oi_1 _18937_ (.A1(_10550_),
    .A2(_10551_),
    .Y(_10552_),
    .B1(net5523));
 sg13g2_a22oi_1 _18938_ (.Y(_10553_),
    .B1(net5369),
    .B2(\atari2600.ram[75][3] ),
    .A2(net5416),
    .A1(\atari2600.ram[72][3] ));
 sg13g2_a22oi_1 _18939_ (.Y(_10554_),
    .B1(net5323),
    .B2(\atari2600.ram[74][3] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][3] ));
 sg13g2_a21oi_1 _18940_ (.A1(_10553_),
    .A2(_10554_),
    .Y(_10555_),
    .B1(net5485));
 sg13g2_nor4_1 _18941_ (.A(_10546_),
    .B(_10549_),
    .C(_10552_),
    .D(_10555_),
    .Y(_10556_));
 sg13g2_a22oi_1 _18942_ (.Y(_10557_),
    .B1(net5380),
    .B2(\atari2600.ram[91][3] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][3] ));
 sg13g2_a22oi_1 _18943_ (.Y(_10558_),
    .B1(net5333),
    .B2(\atari2600.ram[90][3] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][3] ));
 sg13g2_a22oi_1 _18944_ (.Y(_10559_),
    .B1(net5377),
    .B2(\atari2600.ram[99][3] ),
    .A2(net5425),
    .A1(\atari2600.ram[96][3] ));
 sg13g2_a22oi_1 _18945_ (.Y(_10560_),
    .B1(net5332),
    .B2(\atari2600.ram[98][3] ),
    .A2(net5471),
    .A1(\atari2600.ram[97][3] ));
 sg13g2_a21oi_1 _18946_ (.A1(_10559_),
    .A2(_10560_),
    .Y(_10561_),
    .B1(net5508));
 sg13g2_a22oi_1 _18947_ (.Y(_10562_),
    .B1(net5365),
    .B2(\atari2600.ram[103][3] ),
    .A2(net5416),
    .A1(\atari2600.ram[100][3] ));
 sg13g2_a22oi_1 _18948_ (.Y(_10563_),
    .B1(net5322),
    .B2(\atari2600.ram[102][3] ),
    .A2(net5461),
    .A1(\atari2600.ram[101][3] ));
 sg13g2_a21oi_2 _18949_ (.B1(net5521),
    .Y(_10564_),
    .A2(_10563_),
    .A1(_10562_));
 sg13g2_a22oi_1 _18950_ (.Y(_10565_),
    .B1(net5376),
    .B2(\atari2600.ram[107][3] ),
    .A2(net5424),
    .A1(\atari2600.ram[104][3] ));
 sg13g2_a22oi_1 _18951_ (.Y(_10566_),
    .B1(net5316),
    .B2(\atari2600.ram[106][3] ),
    .A2(net5455),
    .A1(\atari2600.ram[105][3] ));
 sg13g2_a21oi_1 _18952_ (.A1(_10565_),
    .A2(_10566_),
    .Y(_10567_),
    .B1(net5482));
 sg13g2_a22oi_1 _18953_ (.Y(_10568_),
    .B1(net5365),
    .B2(\atari2600.ram[111][3] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][3] ));
 sg13g2_a22oi_1 _18954_ (.Y(_10569_),
    .B1(net5319),
    .B2(\atari2600.ram[110][3] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][3] ));
 sg13g2_a21oi_2 _18955_ (.B1(net5495),
    .Y(_10570_),
    .A2(_10569_),
    .A1(_10568_));
 sg13g2_nor4_1 _18956_ (.A(_10561_),
    .B(_10564_),
    .C(_10567_),
    .D(_10570_),
    .Y(_10571_));
 sg13g2_a22oi_1 _18957_ (.Y(_10572_),
    .B1(net5363),
    .B2(\atari2600.ram[123][3] ),
    .A2(net5410),
    .A1(\atari2600.ram[120][3] ));
 sg13g2_a22oi_1 _18958_ (.Y(_10573_),
    .B1(net5317),
    .B2(\atari2600.ram[122][3] ),
    .A2(net5456),
    .A1(\atari2600.ram[121][3] ));
 sg13g2_a21oi_1 _18959_ (.A1(_10572_),
    .A2(_10573_),
    .Y(_10574_),
    .B1(net5482));
 sg13g2_a22oi_1 _18960_ (.Y(_10575_),
    .B1(net5360),
    .B2(\atari2600.ram[127][3] ),
    .A2(net5407),
    .A1(\atari2600.ram[124][3] ));
 sg13g2_a22oi_1 _18961_ (.Y(_10576_),
    .B1(net5312),
    .B2(\atari2600.ram[126][3] ),
    .A2(net5452),
    .A1(\atari2600.ram[125][3] ));
 sg13g2_a21oi_2 _18962_ (.B1(net5494),
    .Y(_10577_),
    .A2(_10576_),
    .A1(_10575_));
 sg13g2_a22oi_1 _18963_ (.Y(_10578_),
    .B1(net5360),
    .B2(\atari2600.ram[119][3] ),
    .A2(net5407),
    .A1(\atari2600.ram[116][3] ));
 sg13g2_a22oi_1 _18964_ (.Y(_10579_),
    .B1(net5312),
    .B2(\atari2600.ram[118][3] ),
    .A2(net5452),
    .A1(\atari2600.ram[117][3] ));
 sg13g2_a21oi_2 _18965_ (.B1(net5520),
    .Y(_10580_),
    .A2(_10579_),
    .A1(_10578_));
 sg13g2_a22oi_1 _18966_ (.Y(_10581_),
    .B1(net5362),
    .B2(\atari2600.ram[115][3] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][3] ));
 sg13g2_a22oi_1 _18967_ (.Y(_10582_),
    .B1(net5312),
    .B2(\atari2600.ram[114][3] ),
    .A2(net5452),
    .A1(\atari2600.ram[113][3] ));
 sg13g2_a21oi_1 _18968_ (.A1(_10581_),
    .A2(_10582_),
    .Y(_10583_),
    .B1(net5510));
 sg13g2_nor4_2 _18969_ (.A(_10574_),
    .B(_10577_),
    .C(_10580_),
    .Y(_10584_),
    .D(_10583_));
 sg13g2_or2_1 _18970_ (.X(_10585_),
    .B(_10584_),
    .A(_09361_));
 sg13g2_a22oi_1 _18971_ (.Y(_10586_),
    .B1(net5379),
    .B2(\atari2600.ram[95][3] ),
    .A2(net5427),
    .A1(\atari2600.ram[92][3] ));
 sg13g2_a22oi_1 _18972_ (.Y(_10587_),
    .B1(net5329),
    .B2(\atari2600.ram[94][3] ),
    .A2(net5468),
    .A1(\atari2600.ram[93][3] ));
 sg13g2_a21oi_1 _18973_ (.A1(_10586_),
    .A2(_10587_),
    .Y(_10588_),
    .B1(net5498));
 sg13g2_a22oi_1 _18974_ (.Y(_10589_),
    .B1(net5374),
    .B2(\atari2600.ram[83][3] ),
    .A2(net5423),
    .A1(\atari2600.ram[80][3] ));
 sg13g2_a22oi_1 _18975_ (.Y(_10590_),
    .B1(net5329),
    .B2(\atari2600.ram[82][3] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][3] ));
 sg13g2_a21oi_1 _18976_ (.A1(_10589_),
    .A2(_10590_),
    .Y(_10591_),
    .B1(net5508));
 sg13g2_a22oi_1 _18977_ (.Y(_10592_),
    .B1(net5380),
    .B2(\atari2600.ram[87][3] ),
    .A2(net5428),
    .A1(\atari2600.ram[84][3] ));
 sg13g2_a22oi_1 _18978_ (.Y(_10593_),
    .B1(net5333),
    .B2(\atari2600.ram[86][3] ),
    .A2(net5472),
    .A1(\atari2600.ram[85][3] ));
 sg13g2_a21oi_1 _18979_ (.A1(_10592_),
    .A2(_10593_),
    .Y(_10594_),
    .B1(net5523));
 sg13g2_o21ai_1 _18980_ (.B1(net5545),
    .Y(_10595_),
    .A1(net5268),
    .A2(_10571_));
 sg13g2_a21oi_1 _18981_ (.A1(_10557_),
    .A2(_10558_),
    .Y(_10596_),
    .B1(net5486));
 sg13g2_nor4_2 _18982_ (.A(_10588_),
    .B(_10591_),
    .C(_10594_),
    .Y(_10597_),
    .D(_10596_));
 sg13g2_nor2_1 _18983_ (.A(net5266),
    .B(_10597_),
    .Y(_10598_));
 sg13g2_o21ai_1 _18984_ (.B1(_10585_),
    .Y(_10599_),
    .A1(net5271),
    .A2(_10556_));
 sg13g2_nor3_2 _18985_ (.A(_10595_),
    .B(_10598_),
    .C(_10599_),
    .Y(_10600_));
 sg13g2_nor2_1 _18986_ (.A(_10543_),
    .B(_10600_),
    .Y(_00004_));
 sg13g2_a22oi_1 _18987_ (.Y(_10601_),
    .B1(net5394),
    .B2(\atari2600.ram[56][4] ),
    .A2(net5443),
    .A1(\atari2600.ram[57][4] ));
 sg13g2_a22oi_1 _18988_ (.Y(_10602_),
    .B1(net5303),
    .B2(\atari2600.ram[58][4] ),
    .A2(net5349),
    .A1(\atari2600.ram[59][4] ));
 sg13g2_a21o_1 _18989_ (.A2(_10602_),
    .A1(_10601_),
    .B1(net5478),
    .X(_10603_));
 sg13g2_a22oi_1 _18990_ (.Y(_10604_),
    .B1(net5348),
    .B2(\atari2600.ram[63][4] ),
    .A2(net5393),
    .A1(\atari2600.ram[60][4] ));
 sg13g2_a22oi_1 _18991_ (.Y(_10605_),
    .B1(net5300),
    .B2(\atari2600.ram[62][4] ),
    .A2(net5440),
    .A1(\atari2600.ram[61][4] ));
 sg13g2_a21oi_1 _18992_ (.A1(_10604_),
    .A2(_10605_),
    .Y(_10606_),
    .B1(net5488));
 sg13g2_a22oi_1 _18993_ (.Y(_10607_),
    .B1(net5346),
    .B2(\atari2600.ram[55][4] ),
    .A2(net5391),
    .A1(\atari2600.ram[52][4] ));
 sg13g2_a22oi_1 _18994_ (.Y(_10608_),
    .B1(net5298),
    .B2(\atari2600.ram[54][4] ),
    .A2(net5438),
    .A1(\atari2600.ram[53][4] ));
 sg13g2_a21oi_1 _18995_ (.A1(_10607_),
    .A2(_10608_),
    .Y(_10609_),
    .B1(net5518));
 sg13g2_a22oi_1 _18996_ (.Y(_10610_),
    .B1(net5348),
    .B2(\atari2600.ram[51][4] ),
    .A2(net5393),
    .A1(\atari2600.ram[48][4] ));
 sg13g2_a22oi_1 _18997_ (.Y(_10611_),
    .B1(net5299),
    .B2(\atari2600.ram[50][4] ),
    .A2(net5439),
    .A1(\atari2600.ram[49][4] ));
 sg13g2_a21oi_1 _18998_ (.A1(_10610_),
    .A2(_10611_),
    .Y(_10612_),
    .B1(net5506));
 sg13g2_nor4_1 _18999_ (.A(net5279),
    .B(_10606_),
    .C(_10609_),
    .D(_10612_),
    .Y(_10613_));
 sg13g2_a22oi_1 _19000_ (.Y(_10614_),
    .B1(net5344),
    .B2(\atari2600.ram[43][4] ),
    .A2(net5389),
    .A1(\atari2600.ram[40][4] ));
 sg13g2_a22oi_1 _19001_ (.Y(_10615_),
    .B1(net5297),
    .B2(\atari2600.ram[42][4] ),
    .A2(net5437),
    .A1(\atari2600.ram[41][4] ));
 sg13g2_a21oi_1 _19002_ (.A1(_10614_),
    .A2(_10615_),
    .Y(_10616_),
    .B1(net5477));
 sg13g2_a22oi_1 _19003_ (.Y(_10617_),
    .B1(net5385),
    .B2(\atari2600.ram[36][4] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][4] ));
 sg13g2_a22oi_1 _19004_ (.Y(_10618_),
    .B1(net5294),
    .B2(\atari2600.ram[38][4] ),
    .A2(net5340),
    .A1(\atari2600.ram[39][4] ));
 sg13g2_a21oi_2 _19005_ (.B1(net5515),
    .Y(_10619_),
    .A2(_10618_),
    .A1(_10617_));
 sg13g2_a22oi_1 _19006_ (.Y(_10620_),
    .B1(net5342),
    .B2(\atari2600.ram[47][4] ),
    .A2(net5391),
    .A1(\atari2600.ram[44][4] ));
 sg13g2_a22oi_1 _19007_ (.Y(_10621_),
    .B1(net5298),
    .B2(\atari2600.ram[46][4] ),
    .A2(net5438),
    .A1(\atari2600.ram[45][4] ));
 sg13g2_a21oi_1 _19008_ (.A1(_10620_),
    .A2(_10621_),
    .Y(_10622_),
    .B1(net5490));
 sg13g2_a22oi_1 _19009_ (.Y(_10623_),
    .B1(net5341),
    .B2(\atari2600.ram[35][4] ),
    .A2(net5389),
    .A1(\atari2600.ram[32][4] ));
 sg13g2_a22oi_1 _19010_ (.Y(_10624_),
    .B1(net5294),
    .B2(\atari2600.ram[34][4] ),
    .A2(net5434),
    .A1(\atari2600.ram[33][4] ));
 sg13g2_a21oi_1 _19011_ (.A1(_10623_),
    .A2(_10624_),
    .Y(_10625_),
    .B1(net5501));
 sg13g2_nor2_1 _19012_ (.A(net5275),
    .B(_10622_),
    .Y(_10626_));
 sg13g2_nor3_2 _19013_ (.A(_10616_),
    .B(_10619_),
    .C(_10625_),
    .Y(_10627_));
 sg13g2_a221oi_1 _19014_ (.B2(_10627_),
    .C1(net5568),
    .B1(_10626_),
    .A1(_10603_),
    .Y(_10628_),
    .A2(_10613_));
 sg13g2_a22oi_1 _19015_ (.Y(_10629_),
    .B1(net5357),
    .B2(\atari2600.ram[23][4] ),
    .A2(net5403),
    .A1(\atari2600.ram[20][4] ));
 sg13g2_a22oi_1 _19016_ (.Y(_10630_),
    .B1(net5304),
    .B2(\atari2600.ram[22][4] ),
    .A2(net5444),
    .A1(\atari2600.ram[21][4] ));
 sg13g2_a21oi_1 _19017_ (.A1(_10629_),
    .A2(_10630_),
    .Y(_10631_),
    .B1(net5517));
 sg13g2_a22oi_1 _19018_ (.Y(_10632_),
    .B1(net5371),
    .B2(\atari2600.ram[27][4] ),
    .A2(net5419),
    .A1(\atari2600.ram[24][4] ));
 sg13g2_a22oi_1 _19019_ (.Y(_10633_),
    .B1(net5326),
    .B2(\atari2600.ram[26][4] ),
    .A2(net5465),
    .A1(\atari2600.ram[25][4] ));
 sg13g2_a21oi_1 _19020_ (.A1(_10632_),
    .A2(_10633_),
    .Y(_10634_),
    .B1(net5487));
 sg13g2_a22oi_1 _19021_ (.Y(_10635_),
    .B1(net5374),
    .B2(\atari2600.ram[31][4] ),
    .A2(net5423),
    .A1(\atari2600.ram[28][4] ));
 sg13g2_a22oi_1 _19022_ (.Y(_10636_),
    .B1(net5330),
    .B2(\atari2600.ram[30][4] ),
    .A2(net5469),
    .A1(\atari2600.ram[29][4] ));
 sg13g2_a21oi_2 _19023_ (.B1(net5492),
    .Y(_10637_),
    .A2(_10636_),
    .A1(_10635_));
 sg13g2_a22oi_1 _19024_ (.Y(_10638_),
    .B1(net5358),
    .B2(\atari2600.ram[19][4] ),
    .A2(net5405),
    .A1(\atari2600.ram[16][4] ));
 sg13g2_a22oi_1 _19025_ (.Y(_10639_),
    .B1(net5310),
    .B2(\atari2600.ram[18][4] ),
    .A2(net5450),
    .A1(\atari2600.ram[17][4] ));
 sg13g2_a21oi_1 _19026_ (.A1(_10638_),
    .A2(_10639_),
    .Y(_10640_),
    .B1(net5505));
 sg13g2_or4_2 _19027_ (.A(_10631_),
    .B(_10634_),
    .C(_10637_),
    .D(_10640_),
    .X(_10641_));
 sg13g2_a22oi_1 _19028_ (.Y(_10642_),
    .B1(net5353),
    .B2(\atari2600.ram[3][4] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][4] ));
 sg13g2_a22oi_1 _19029_ (.Y(_10643_),
    .B1(net5307),
    .B2(\atari2600.ram[2][4] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][4] ));
 sg13g2_a21oi_1 _19030_ (.A1(_10642_),
    .A2(_10643_),
    .Y(_10644_),
    .B1(net5503));
 sg13g2_a22oi_1 _19031_ (.Y(_10645_),
    .B1(net5349),
    .B2(\atari2600.ram[11][4] ),
    .A2(net5394),
    .A1(\atari2600.ram[8][4] ));
 sg13g2_a22oi_1 _19032_ (.Y(_10646_),
    .B1(net5296),
    .B2(\atari2600.ram[10][4] ),
    .A2(net5436),
    .A1(\atari2600.ram[9][4] ));
 sg13g2_a21oi_1 _19033_ (.A1(_10645_),
    .A2(_10646_),
    .Y(_10647_),
    .B1(net5479));
 sg13g2_a22oi_1 _19034_ (.Y(_10648_),
    .B1(net5355),
    .B2(\atari2600.ram[7][4] ),
    .A2(net5401),
    .A1(\atari2600.ram[4][4] ));
 sg13g2_a22oi_1 _19035_ (.Y(_10649_),
    .B1(net5308),
    .B2(\atari2600.ram[6][4] ),
    .A2(net5448),
    .A1(\atari2600.ram[5][4] ));
 sg13g2_a21oi_1 _19036_ (.A1(_10648_),
    .A2(_10649_),
    .Y(_10650_),
    .B1(net5516));
 sg13g2_a22oi_1 _19037_ (.Y(_10651_),
    .B1(net5357),
    .B2(\atari2600.ram[15][4] ),
    .A2(net5404),
    .A1(\atari2600.ram[12][4] ));
 sg13g2_a22oi_1 _19038_ (.Y(_10652_),
    .B1(net5306),
    .B2(\atari2600.ram[14][4] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][4] ));
 sg13g2_a21oi_1 _19039_ (.A1(_10651_),
    .A2(_10652_),
    .Y(_10653_),
    .B1(net5491));
 sg13g2_or4_1 _19040_ (.A(_10644_),
    .B(_10647_),
    .C(_10650_),
    .D(_10653_),
    .X(_10654_));
 sg13g2_a221oi_1 _19041_ (.B2(_09105_),
    .C1(_10628_),
    .B1(_10654_),
    .A1(_09319_),
    .Y(_10655_),
    .A2(_10641_));
 sg13g2_a22oi_1 _19042_ (.Y(_10656_),
    .B1(net5412),
    .B2(\atari2600.ram[100][4] ),
    .A2(net5458),
    .A1(\atari2600.ram[101][4] ));
 sg13g2_a22oi_1 _19043_ (.Y(_10657_),
    .B1(net5319),
    .B2(\atari2600.ram[102][4] ),
    .A2(net5366),
    .A1(\atari2600.ram[103][4] ));
 sg13g2_a21oi_1 _19044_ (.A1(_10656_),
    .A2(_10657_),
    .Y(_10658_),
    .B1(net5521));
 sg13g2_a22oi_1 _19045_ (.Y(_10659_),
    .B1(net5359),
    .B2(\atari2600.ram[111][4] ),
    .A2(net5406),
    .A1(\atari2600.ram[108][4] ));
 sg13g2_a22oi_1 _19046_ (.Y(_10660_),
    .B1(net5314),
    .B2(\atari2600.ram[110][4] ),
    .A2(net5453),
    .A1(\atari2600.ram[109][4] ));
 sg13g2_a21o_1 _19047_ (.A2(_10660_),
    .A1(_10659_),
    .B1(net5494),
    .X(_10661_));
 sg13g2_a22oi_1 _19048_ (.Y(_10662_),
    .B1(net5359),
    .B2(\atari2600.ram[107][4] ),
    .A2(net5406),
    .A1(\atari2600.ram[104][4] ));
 sg13g2_a22oi_1 _19049_ (.Y(_10663_),
    .B1(net5314),
    .B2(\atari2600.ram[106][4] ),
    .A2(net5453),
    .A1(\atari2600.ram[105][4] ));
 sg13g2_a21oi_1 _19050_ (.A1(_10662_),
    .A2(_10663_),
    .Y(_10664_),
    .B1(net5483));
 sg13g2_a22oi_1 _19051_ (.Y(_10665_),
    .B1(net5369),
    .B2(\atari2600.ram[99][4] ),
    .A2(net5416),
    .A1(\atari2600.ram[96][4] ));
 sg13g2_a22oi_1 _19052_ (.Y(_10666_),
    .B1(net5322),
    .B2(\atari2600.ram[98][4] ),
    .A2(net5461),
    .A1(\atari2600.ram[97][4] ));
 sg13g2_a21oi_1 _19053_ (.A1(_10665_),
    .A2(_10666_),
    .Y(_10667_),
    .B1(net5510));
 sg13g2_nor4_1 _19054_ (.A(net5276),
    .B(_10658_),
    .C(_10664_),
    .D(_10667_),
    .Y(_10668_));
 sg13g2_a22oi_1 _19055_ (.Y(_10669_),
    .B1(net5312),
    .B2(\atari2600.ram[114][4] ),
    .A2(net5452),
    .A1(\atari2600.ram[113][4] ));
 sg13g2_a22oi_1 _19056_ (.Y(_10670_),
    .B1(net5362),
    .B2(\atari2600.ram[115][4] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][4] ));
 sg13g2_a21oi_1 _19057_ (.A1(_10669_),
    .A2(_10670_),
    .Y(_10671_),
    .B1(net5510));
 sg13g2_a22oi_1 _19058_ (.Y(_10672_),
    .B1(net5359),
    .B2(\atari2600.ram[127][4] ),
    .A2(net5406),
    .A1(\atari2600.ram[124][4] ));
 sg13g2_a22oi_1 _19059_ (.Y(_10673_),
    .B1(net5314),
    .B2(\atari2600.ram[126][4] ),
    .A2(net5453),
    .A1(\atari2600.ram[125][4] ));
 sg13g2_a21o_1 _19060_ (.A2(_10673_),
    .A1(_10672_),
    .B1(net5494),
    .X(_10674_));
 sg13g2_a22oi_1 _19061_ (.Y(_10675_),
    .B1(net5409),
    .B2(\atari2600.ram[120][4] ),
    .A2(net5455),
    .A1(\atari2600.ram[121][4] ));
 sg13g2_a22oi_1 _19062_ (.Y(_10676_),
    .B1(net5316),
    .B2(\atari2600.ram[122][4] ),
    .A2(net5364),
    .A1(\atari2600.ram[123][4] ));
 sg13g2_a21oi_1 _19063_ (.A1(_10675_),
    .A2(_10676_),
    .Y(_10677_),
    .B1(net5482));
 sg13g2_a22oi_1 _19064_ (.Y(_10678_),
    .B1(net5359),
    .B2(\atari2600.ram[119][4] ),
    .A2(net5406),
    .A1(\atari2600.ram[116][4] ));
 sg13g2_a22oi_1 _19065_ (.Y(_10679_),
    .B1(net5315),
    .B2(\atari2600.ram[118][4] ),
    .A2(net5454),
    .A1(\atari2600.ram[117][4] ));
 sg13g2_a21oi_1 _19066_ (.A1(_10678_),
    .A2(_10679_),
    .Y(_10680_),
    .B1(net5520));
 sg13g2_nor4_1 _19067_ (.A(net5283),
    .B(_10671_),
    .C(_10677_),
    .D(_10680_),
    .Y(_10681_));
 sg13g2_a221oi_1 _19068_ (.B2(_10681_),
    .C1(net5571),
    .B1(_10674_),
    .A1(_10661_),
    .Y(_10682_),
    .A2(_10668_));
 sg13g2_a22oi_1 _19069_ (.Y(_10683_),
    .B1(net5381),
    .B2(\atari2600.ram[87][4] ),
    .A2(net5429),
    .A1(\atari2600.ram[84][4] ));
 sg13g2_a22oi_1 _19070_ (.Y(_10684_),
    .B1(net5335),
    .B2(\atari2600.ram[86][4] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][4] ));
 sg13g2_a21oi_1 _19071_ (.A1(_10683_),
    .A2(_10684_),
    .Y(_10685_),
    .B1(net5523));
 sg13g2_a22oi_1 _19072_ (.Y(_10686_),
    .B1(net5380),
    .B2(\atari2600.ram[95][4] ),
    .A2(net5427),
    .A1(\atari2600.ram[92][4] ));
 sg13g2_a22oi_1 _19073_ (.Y(_10687_),
    .B1(net5333),
    .B2(\atari2600.ram[94][4] ),
    .A2(net5472),
    .A1(\atari2600.ram[93][4] ));
 sg13g2_a21oi_1 _19074_ (.A1(_10686_),
    .A2(_10687_),
    .Y(_10688_),
    .B1(net5499));
 sg13g2_a22oi_1 _19075_ (.Y(_10689_),
    .B1(net5375),
    .B2(\atari2600.ram[83][4] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][4] ));
 sg13g2_a22oi_1 _19076_ (.Y(_10690_),
    .B1(net5329),
    .B2(\atari2600.ram[82][4] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][4] ));
 sg13g2_a21oi_2 _19077_ (.B1(net5509),
    .Y(_10691_),
    .A2(_10690_),
    .A1(_10689_));
 sg13g2_a22oi_1 _19078_ (.Y(_10692_),
    .B1(net5378),
    .B2(\atari2600.ram[71][4] ),
    .A2(net5426),
    .A1(\atari2600.ram[68][4] ));
 sg13g2_a22oi_1 _19079_ (.Y(_10693_),
    .B1(net5331),
    .B2(\atari2600.ram[70][4] ),
    .A2(net5470),
    .A1(\atari2600.ram[69][4] ));
 sg13g2_a21oi_1 _19080_ (.A1(_10692_),
    .A2(_10693_),
    .Y(_10694_),
    .B1(net5523));
 sg13g2_a22oi_1 _19081_ (.Y(_10695_),
    .B1(net5378),
    .B2(\atari2600.ram[67][4] ),
    .A2(net5426),
    .A1(\atari2600.ram[64][4] ));
 sg13g2_a22oi_1 _19082_ (.Y(_10696_),
    .B1(net5331),
    .B2(\atari2600.ram[66][4] ),
    .A2(net5470),
    .A1(\atari2600.ram[65][4] ));
 sg13g2_a21oi_1 _19083_ (.A1(_10695_),
    .A2(_10696_),
    .Y(_10697_),
    .B1(net5512));
 sg13g2_a22oi_1 _19084_ (.Y(_10698_),
    .B1(net5367),
    .B2(\atari2600.ram[79][4] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][4] ));
 sg13g2_a22oi_1 _19085_ (.Y(_10699_),
    .B1(net5320),
    .B2(\atari2600.ram[78][4] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][4] ));
 sg13g2_a21oi_2 _19086_ (.B1(net5496),
    .Y(_10700_),
    .A2(_10699_),
    .A1(_10698_));
 sg13g2_a22oi_1 _19087_ (.Y(_10701_),
    .B1(net5368),
    .B2(\atari2600.ram[75][4] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][4] ));
 sg13g2_a22oi_1 _19088_ (.Y(_10702_),
    .B1(net5323),
    .B2(\atari2600.ram[74][4] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][4] ));
 sg13g2_a21oi_1 _19089_ (.A1(_10701_),
    .A2(_10702_),
    .Y(_10703_),
    .B1(net5486));
 sg13g2_nor4_2 _19090_ (.A(_10694_),
    .B(_10697_),
    .C(_10700_),
    .Y(_10704_),
    .D(_10703_));
 sg13g2_a22oi_1 _19091_ (.Y(_10705_),
    .B1(net5380),
    .B2(\atari2600.ram[91][4] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][4] ));
 sg13g2_a22oi_1 _19092_ (.Y(_10706_),
    .B1(net5334),
    .B2(\atari2600.ram[90][4] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][4] ));
 sg13g2_a21oi_1 _19093_ (.A1(_10705_),
    .A2(_10706_),
    .Y(_10707_),
    .B1(net5486));
 sg13g2_nor4_2 _19094_ (.A(_10685_),
    .B(_10688_),
    .C(_10691_),
    .Y(_10708_),
    .D(_10707_));
 sg13g2_nor2_1 _19095_ (.A(net5266),
    .B(_10708_),
    .Y(_10709_));
 sg13g2_o21ai_1 _19096_ (.B1(net5545),
    .Y(_10710_),
    .A1(net5271),
    .A2(_10704_));
 sg13g2_nor3_2 _19097_ (.A(_10682_),
    .B(_10709_),
    .C(_10710_),
    .Y(_10711_));
 sg13g2_a21oi_1 _19098_ (.A1(net5543),
    .A2(_10655_),
    .Y(_00005_),
    .B1(_10711_));
 sg13g2_a22oi_1 _19099_ (.Y(_10712_),
    .B1(net5390),
    .B2(\atari2600.ram[40][5] ),
    .A2(net5436),
    .A1(\atari2600.ram[41][5] ));
 sg13g2_a22oi_1 _19100_ (.Y(_10713_),
    .B1(net5296),
    .B2(\atari2600.ram[42][5] ),
    .A2(net5345),
    .A1(\atari2600.ram[43][5] ));
 sg13g2_a21o_1 _19101_ (.A2(_10713_),
    .A1(_10712_),
    .B1(net5479),
    .X(_10714_));
 sg13g2_a22oi_1 _19102_ (.Y(_10715_),
    .B1(net5340),
    .B2(\atari2600.ram[39][5] ),
    .A2(net5385),
    .A1(\atari2600.ram[36][5] ));
 sg13g2_a22oi_1 _19103_ (.Y(_10716_),
    .B1(net5293),
    .B2(\atari2600.ram[38][5] ),
    .A2(net5434),
    .A1(\atari2600.ram[37][5] ));
 sg13g2_a21oi_2 _19104_ (.B1(net5515),
    .Y(_10717_),
    .A2(_10716_),
    .A1(_10715_));
 sg13g2_a22oi_1 _19105_ (.Y(_10718_),
    .B1(net5342),
    .B2(\atari2600.ram[47][5] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][5] ));
 sg13g2_a22oi_1 _19106_ (.Y(_10719_),
    .B1(net5295),
    .B2(\atari2600.ram[46][5] ),
    .A2(net5435),
    .A1(\atari2600.ram[45][5] ));
 sg13g2_a21oi_1 _19107_ (.A1(_10718_),
    .A2(_10719_),
    .Y(_10720_),
    .B1(net5490));
 sg13g2_a22oi_1 _19108_ (.Y(_10721_),
    .B1(net5343),
    .B2(\atari2600.ram[35][5] ),
    .A2(net5388),
    .A1(\atari2600.ram[32][5] ));
 sg13g2_a22oi_1 _19109_ (.Y(_10722_),
    .B1(net5295),
    .B2(\atari2600.ram[34][5] ),
    .A2(net5435),
    .A1(\atari2600.ram[33][5] ));
 sg13g2_a21oi_1 _19110_ (.A1(_10721_),
    .A2(_10722_),
    .Y(_10723_),
    .B1(net5501));
 sg13g2_nor4_2 _19111_ (.A(net5275),
    .B(_10717_),
    .C(_10720_),
    .Y(_10724_),
    .D(_10723_));
 sg13g2_a22oi_1 _19112_ (.Y(_10725_),
    .B1(net5351),
    .B2(\atari2600.ram[59][5] ),
    .A2(net5396),
    .A1(\atari2600.ram[56][5] ));
 sg13g2_a22oi_1 _19113_ (.Y(_10726_),
    .B1(net5303),
    .B2(\atari2600.ram[58][5] ),
    .A2(net5443),
    .A1(\atari2600.ram[57][5] ));
 sg13g2_a21oi_1 _19114_ (.A1(_10725_),
    .A2(_10726_),
    .Y(_10727_),
    .B1(net5478));
 sg13g2_nor2_1 _19115_ (.A(net5279),
    .B(_10727_),
    .Y(_10728_));
 sg13g2_a22oi_1 _19116_ (.Y(_10729_),
    .B1(net5391),
    .B2(\atari2600.ram[52][5] ),
    .A2(net5438),
    .A1(\atari2600.ram[53][5] ));
 sg13g2_a22oi_1 _19117_ (.Y(_10730_),
    .B1(net5298),
    .B2(\atari2600.ram[54][5] ),
    .A2(net5346),
    .A1(\atari2600.ram[55][5] ));
 sg13g2_a21oi_1 _19118_ (.A1(_10729_),
    .A2(_10730_),
    .Y(_10731_),
    .B1(net5518));
 sg13g2_a22oi_1 _19119_ (.Y(_10732_),
    .B1(net5299),
    .B2(\atari2600.ram[50][5] ),
    .A2(net5439),
    .A1(\atari2600.ram[49][5] ));
 sg13g2_a22oi_1 _19120_ (.Y(_10733_),
    .B1(net5346),
    .B2(\atari2600.ram[51][5] ),
    .A2(net5393),
    .A1(\atari2600.ram[48][5] ));
 sg13g2_a21oi_1 _19121_ (.A1(_10732_),
    .A2(_10733_),
    .Y(_10734_),
    .B1(net5502));
 sg13g2_a22oi_1 _19122_ (.Y(_10735_),
    .B1(net5347),
    .B2(\atari2600.ram[63][5] ),
    .A2(net5392),
    .A1(\atari2600.ram[60][5] ));
 sg13g2_a22oi_1 _19123_ (.Y(_10736_),
    .B1(net5300),
    .B2(\atari2600.ram[62][5] ),
    .A2(net5440),
    .A1(\atari2600.ram[61][5] ));
 sg13g2_a21oi_2 _19124_ (.B1(net5488),
    .Y(_10737_),
    .A2(_10736_),
    .A1(_10735_));
 sg13g2_nor3_1 _19125_ (.A(_10731_),
    .B(_10734_),
    .C(_10737_),
    .Y(_10738_));
 sg13g2_a221oi_1 _19126_ (.B2(_10738_),
    .C1(net5568),
    .B1(_10728_),
    .A1(_10714_),
    .Y(_10739_),
    .A2(_10724_));
 sg13g2_a22oi_1 _19127_ (.Y(_10740_),
    .B1(net5373),
    .B2(\atari2600.ram[31][5] ),
    .A2(net5423),
    .A1(\atari2600.ram[28][5] ));
 sg13g2_a22oi_1 _19128_ (.Y(_10741_),
    .B1(net5330),
    .B2(\atari2600.ram[30][5] ),
    .A2(net5469),
    .A1(\atari2600.ram[29][5] ));
 sg13g2_a21oi_1 _19129_ (.A1(_10740_),
    .A2(_10741_),
    .Y(_10742_),
    .B1(net5493));
 sg13g2_a22oi_1 _19130_ (.Y(_10743_),
    .B1(net5326),
    .B2(\atari2600.ram[26][5] ),
    .A2(net5419),
    .A1(\atari2600.ram[24][5] ));
 sg13g2_a22oi_1 _19131_ (.Y(_10744_),
    .B1(net5371),
    .B2(\atari2600.ram[27][5] ),
    .A2(net5466),
    .A1(\atari2600.ram[25][5] ));
 sg13g2_a21oi_1 _19132_ (.A1(_10743_),
    .A2(_10744_),
    .Y(_10745_),
    .B1(net5481));
 sg13g2_a22oi_1 _19133_ (.Y(_10746_),
    .B1(net5358),
    .B2(\atari2600.ram[19][5] ),
    .A2(net5405),
    .A1(\atari2600.ram[16][5] ));
 sg13g2_a22oi_1 _19134_ (.Y(_10747_),
    .B1(net5310),
    .B2(\atari2600.ram[18][5] ),
    .A2(net5450),
    .A1(\atari2600.ram[17][5] ));
 sg13g2_a21oi_2 _19135_ (.B1(net5504),
    .Y(_10748_),
    .A2(_10747_),
    .A1(_10746_));
 sg13g2_a22oi_1 _19136_ (.Y(_10749_),
    .B1(net5371),
    .B2(\atari2600.ram[23][5] ),
    .A2(net5419),
    .A1(\atari2600.ram[20][5] ));
 sg13g2_a22oi_1 _19137_ (.Y(_10750_),
    .B1(net5326),
    .B2(\atari2600.ram[22][5] ),
    .A2(net5465),
    .A1(\atari2600.ram[21][5] ));
 sg13g2_a21oi_1 _19138_ (.A1(_10749_),
    .A2(_10750_),
    .Y(_10751_),
    .B1(net5519));
 sg13g2_nor4_2 _19139_ (.A(_10742_),
    .B(_10745_),
    .C(_10748_),
    .Y(_10752_),
    .D(_10751_));
 sg13g2_a22oi_1 _19140_ (.Y(_10753_),
    .B1(net5355),
    .B2(\atari2600.ram[7][5] ),
    .A2(net5399),
    .A1(\atari2600.ram[4][5] ));
 sg13g2_a22oi_1 _19141_ (.Y(_10754_),
    .B1(net5311),
    .B2(\atari2600.ram[6][5] ),
    .A2(net5451),
    .A1(\atari2600.ram[5][5] ));
 sg13g2_a21oi_2 _19142_ (.B1(net5516),
    .Y(_10755_),
    .A2(_10754_),
    .A1(_10753_));
 sg13g2_a22oi_1 _19143_ (.Y(_10756_),
    .B1(net5344),
    .B2(\atari2600.ram[11][5] ),
    .A2(net5389),
    .A1(\atari2600.ram[8][5] ));
 sg13g2_a22oi_1 _19144_ (.Y(_10757_),
    .B1(net5297),
    .B2(\atari2600.ram[10][5] ),
    .A2(net5437),
    .A1(\atari2600.ram[9][5] ));
 sg13g2_a21oi_2 _19145_ (.B1(net5477),
    .Y(_10758_),
    .A2(_10757_),
    .A1(_10756_));
 sg13g2_a22oi_1 _19146_ (.Y(_10759_),
    .B1(net5353),
    .B2(\atari2600.ram[3][5] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][5] ));
 sg13g2_a22oi_1 _19147_ (.Y(_10760_),
    .B1(net5307),
    .B2(\atari2600.ram[2][5] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][5] ));
 sg13g2_a21oi_2 _19148_ (.B1(net5503),
    .Y(_10761_),
    .A2(_10760_),
    .A1(_10759_));
 sg13g2_a22oi_1 _19149_ (.Y(_10762_),
    .B1(net5354),
    .B2(\atari2600.ram[15][5] ),
    .A2(net5399),
    .A1(\atari2600.ram[12][5] ));
 sg13g2_a22oi_1 _19150_ (.Y(_10763_),
    .B1(net5306),
    .B2(\atari2600.ram[14][5] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][5] ));
 sg13g2_a21oi_1 _19151_ (.A1(_10762_),
    .A2(_10763_),
    .Y(_10764_),
    .B1(net5491));
 sg13g2_nor4_2 _19152_ (.A(_10755_),
    .B(_10758_),
    .C(_10761_),
    .Y(_10765_),
    .D(_10764_));
 sg13g2_nor2_1 _19153_ (.A(net5270),
    .B(_10765_),
    .Y(_10766_));
 sg13g2_o21ai_1 _19154_ (.B1(net5542),
    .Y(_10767_),
    .A1(net5264),
    .A2(_10752_));
 sg13g2_nor3_1 _19155_ (.A(_10739_),
    .B(_10766_),
    .C(_10767_),
    .Y(_10768_));
 sg13g2_a22oi_1 _19156_ (.Y(_10769_),
    .B1(net5304),
    .B2(\atari2600.ram[114][5] ),
    .A2(net5444),
    .A1(\atari2600.ram[113][5] ));
 sg13g2_a221oi_1 _19157_ (.B2(\atari2600.ram[115][5] ),
    .C1(net5281),
    .B1(net5350),
    .A1(\atari2600.ram[112][5] ),
    .Y(_10770_),
    .A2(net5395));
 sg13g2_a21oi_1 _19158_ (.A1(_10769_),
    .A2(_10770_),
    .Y(_10771_),
    .B1(_09293_));
 sg13g2_a22oi_1 _19159_ (.Y(_10772_),
    .B1(net5363),
    .B2(\atari2600.ram[123][5] ),
    .A2(net5410),
    .A1(\atari2600.ram[120][5] ));
 sg13g2_a22oi_1 _19160_ (.Y(_10773_),
    .B1(net5317),
    .B2(\atari2600.ram[122][5] ),
    .A2(net5456),
    .A1(\atari2600.ram[121][5] ));
 sg13g2_a21oi_1 _19161_ (.A1(_10772_),
    .A2(_10773_),
    .Y(_10774_),
    .B1(net5482));
 sg13g2_a22oi_1 _19162_ (.Y(_10775_),
    .B1(net5408),
    .B2(\atari2600.ram[116][5] ),
    .A2(net5456),
    .A1(\atari2600.ram[117][5] ));
 sg13g2_a22oi_1 _19163_ (.Y(_10776_),
    .B1(net5317),
    .B2(\atari2600.ram[118][5] ),
    .A2(net5362),
    .A1(\atari2600.ram[119][5] ));
 sg13g2_a21oi_1 _19164_ (.A1(_10775_),
    .A2(_10776_),
    .Y(_10777_),
    .B1(net5520));
 sg13g2_a22oi_1 _19165_ (.Y(_10778_),
    .B1(net5360),
    .B2(\atari2600.ram[127][5] ),
    .A2(net5407),
    .A1(\atari2600.ram[124][5] ));
 sg13g2_a22oi_1 _19166_ (.Y(_10779_),
    .B1(net5312),
    .B2(\atari2600.ram[126][5] ),
    .A2(net5452),
    .A1(\atari2600.ram[125][5] ));
 sg13g2_a21oi_2 _19167_ (.B1(net5489),
    .Y(_10780_),
    .A2(_10779_),
    .A1(_10778_));
 sg13g2_nor4_2 _19168_ (.A(_10771_),
    .B(_10774_),
    .C(_10777_),
    .Y(_10781_),
    .D(_10780_));
 sg13g2_a22oi_1 _19169_ (.Y(_10782_),
    .B1(net5359),
    .B2(\atari2600.ram[111][5] ),
    .A2(net5406),
    .A1(\atari2600.ram[108][5] ));
 sg13g2_a22oi_1 _19170_ (.Y(_10783_),
    .B1(net5314),
    .B2(\atari2600.ram[110][5] ),
    .A2(net5453),
    .A1(\atari2600.ram[109][5] ));
 sg13g2_a21oi_1 _19171_ (.A1(_10782_),
    .A2(_10783_),
    .Y(_10784_),
    .B1(net5494));
 sg13g2_nand2b_1 _19172_ (.Y(_10785_),
    .B(net5281),
    .A_N(_10784_));
 sg13g2_a22oi_1 _19173_ (.Y(_10786_),
    .B1(net5409),
    .B2(\atari2600.ram[104][5] ),
    .A2(net5455),
    .A1(\atari2600.ram[105][5] ));
 sg13g2_a22oi_1 _19174_ (.Y(_10787_),
    .B1(net5316),
    .B2(\atari2600.ram[106][5] ),
    .A2(net5363),
    .A1(\atari2600.ram[107][5] ));
 sg13g2_a21oi_1 _19175_ (.A1(_10786_),
    .A2(_10787_),
    .Y(_10788_),
    .B1(net5483));
 sg13g2_a22oi_1 _19176_ (.Y(_10789_),
    .B1(net5363),
    .B2(\atari2600.ram[99][5] ),
    .A2(net5409),
    .A1(\atari2600.ram[96][5] ));
 sg13g2_a22oi_1 _19177_ (.Y(_10790_),
    .B1(net5322),
    .B2(\atari2600.ram[98][5] ),
    .A2(net5461),
    .A1(\atari2600.ram[97][5] ));
 sg13g2_a21oi_1 _19178_ (.A1(_10789_),
    .A2(_10790_),
    .Y(_10791_),
    .B1(net5510));
 sg13g2_a22oi_1 _19179_ (.Y(_10792_),
    .B1(net5359),
    .B2(\atari2600.ram[103][5] ),
    .A2(net5412),
    .A1(\atari2600.ram[100][5] ));
 sg13g2_a22oi_1 _19180_ (.Y(_10793_),
    .B1(net5321),
    .B2(\atari2600.ram[102][5] ),
    .A2(net5460),
    .A1(\atari2600.ram[101][5] ));
 sg13g2_a21oi_1 _19181_ (.A1(_10792_),
    .A2(_10793_),
    .Y(_10794_),
    .B1(net5520));
 sg13g2_nor4_1 _19182_ (.A(_10785_),
    .B(_10788_),
    .C(_10791_),
    .D(_10794_),
    .Y(_10795_));
 sg13g2_nor3_2 _19183_ (.A(net5571),
    .B(_10781_),
    .C(_10795_),
    .Y(_10796_));
 sg13g2_a22oi_1 _19184_ (.Y(_10797_),
    .B1(net5368),
    .B2(\atari2600.ram[75][5] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][5] ));
 sg13g2_a22oi_1 _19185_ (.Y(_10798_),
    .B1(net5323),
    .B2(\atari2600.ram[74][5] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][5] ));
 sg13g2_a21oi_1 _19186_ (.A1(_10797_),
    .A2(_10798_),
    .Y(_10799_),
    .B1(net5486));
 sg13g2_a22oi_1 _19187_ (.Y(_10800_),
    .B1(net5378),
    .B2(\atari2600.ram[67][5] ),
    .A2(net5426),
    .A1(\atari2600.ram[64][5] ));
 sg13g2_a22oi_1 _19188_ (.Y(_10801_),
    .B1(net5331),
    .B2(\atari2600.ram[66][5] ),
    .A2(net5470),
    .A1(\atari2600.ram[65][5] ));
 sg13g2_a21oi_1 _19189_ (.A1(_10800_),
    .A2(_10801_),
    .Y(_10802_),
    .B1(net5511));
 sg13g2_a22oi_1 _19190_ (.Y(_10803_),
    .B1(net5378),
    .B2(\atari2600.ram[71][5] ),
    .A2(net5426),
    .A1(\atari2600.ram[68][5] ));
 sg13g2_a22oi_1 _19191_ (.Y(_10804_),
    .B1(net5332),
    .B2(\atari2600.ram[70][5] ),
    .A2(net5471),
    .A1(\atari2600.ram[69][5] ));
 sg13g2_a21oi_2 _19192_ (.B1(net5524),
    .Y(_10805_),
    .A2(_10804_),
    .A1(_10803_));
 sg13g2_a22oi_1 _19193_ (.Y(_10806_),
    .B1(net5367),
    .B2(\atari2600.ram[79][5] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][5] ));
 sg13g2_a22oi_1 _19194_ (.Y(_10807_),
    .B1(net5320),
    .B2(\atari2600.ram[78][5] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][5] ));
 sg13g2_a21oi_2 _19195_ (.B1(net5496),
    .Y(_10808_),
    .A2(_10807_),
    .A1(_10806_));
 sg13g2_nor4_2 _19196_ (.A(_10799_),
    .B(_10802_),
    .C(_10805_),
    .Y(_10809_),
    .D(_10808_));
 sg13g2_a22oi_1 _19197_ (.Y(_10810_),
    .B1(net5374),
    .B2(\atari2600.ram[83][5] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][5] ));
 sg13g2_a22oi_1 _19198_ (.Y(_10811_),
    .B1(net5329),
    .B2(\atari2600.ram[82][5] ),
    .A2(net5468),
    .A1(\atari2600.ram[81][5] ));
 sg13g2_a21oi_1 _19199_ (.A1(_10810_),
    .A2(_10811_),
    .Y(_10812_),
    .B1(net5508));
 sg13g2_a22oi_1 _19200_ (.Y(_10813_),
    .B1(net5379),
    .B2(\atari2600.ram[95][5] ),
    .A2(net5425),
    .A1(\atari2600.ram[92][5] ));
 sg13g2_a22oi_1 _19201_ (.Y(_10814_),
    .B1(net5333),
    .B2(\atari2600.ram[94][5] ),
    .A2(net5472),
    .A1(\atari2600.ram[93][5] ));
 sg13g2_a21oi_1 _19202_ (.A1(_10813_),
    .A2(_10814_),
    .Y(_10815_),
    .B1(net5499));
 sg13g2_a22oi_1 _19203_ (.Y(_10816_),
    .B1(net5380),
    .B2(\atari2600.ram[91][5] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][5] ));
 sg13g2_a22oi_1 _19204_ (.Y(_10817_),
    .B1(net5334),
    .B2(\atari2600.ram[90][5] ),
    .A2(net5473),
    .A1(\atari2600.ram[89][5] ));
 sg13g2_a21oi_1 _19205_ (.A1(_10816_),
    .A2(_10817_),
    .Y(_10818_),
    .B1(net5486));
 sg13g2_a22oi_1 _19206_ (.Y(_10819_),
    .B1(net5381),
    .B2(\atari2600.ram[87][5] ),
    .A2(net5429),
    .A1(\atari2600.ram[84][5] ));
 sg13g2_a22oi_1 _19207_ (.Y(_10820_),
    .B1(net5335),
    .B2(\atari2600.ram[86][5] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][5] ));
 sg13g2_a21oi_1 _19208_ (.A1(_10819_),
    .A2(_10820_),
    .Y(_10821_),
    .B1(net5525));
 sg13g2_nor4_2 _19209_ (.A(_10812_),
    .B(_10815_),
    .C(_10818_),
    .Y(_10822_),
    .D(_10821_));
 sg13g2_nor2_1 _19210_ (.A(net5266),
    .B(_10822_),
    .Y(_10823_));
 sg13g2_o21ai_1 _19211_ (.B1(net5545),
    .Y(_10824_),
    .A1(net5271),
    .A2(_10809_));
 sg13g2_nor3_2 _19212_ (.A(_10796_),
    .B(_10823_),
    .C(_10824_),
    .Y(_10825_));
 sg13g2_nor2_1 _19213_ (.A(_10768_),
    .B(_10825_),
    .Y(_00006_));
 sg13g2_a22oi_1 _19214_ (.Y(_10826_),
    .B1(net5360),
    .B2(\atari2600.ram[119][6] ),
    .A2(net5407),
    .A1(\atari2600.ram[116][6] ));
 sg13g2_a22oi_1 _19215_ (.Y(_10827_),
    .B1(net5313),
    .B2(\atari2600.ram[118][6] ),
    .A2(net5454),
    .A1(\atari2600.ram[117][6] ));
 sg13g2_a21oi_2 _19216_ (.B1(net5520),
    .Y(_10828_),
    .A2(_10827_),
    .A1(_10826_));
 sg13g2_a22oi_1 _19217_ (.Y(_10829_),
    .B1(net5362),
    .B2(\atari2600.ram[115][6] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][6] ));
 sg13g2_a22oi_1 _19218_ (.Y(_10830_),
    .B1(net5317),
    .B2(\atari2600.ram[114][6] ),
    .A2(net5456),
    .A1(\atari2600.ram[113][6] ));
 sg13g2_a21oi_1 _19219_ (.A1(_10829_),
    .A2(_10830_),
    .Y(_10831_),
    .B1(net5506));
 sg13g2_a22oi_1 _19220_ (.Y(_10832_),
    .B1(net5363),
    .B2(\atari2600.ram[123][6] ),
    .A2(net5408),
    .A1(\atari2600.ram[120][6] ));
 sg13g2_a22oi_1 _19221_ (.Y(_10833_),
    .B1(net5317),
    .B2(\atari2600.ram[122][6] ),
    .A2(net5456),
    .A1(\atari2600.ram[121][6] ));
 sg13g2_a21oi_1 _19222_ (.A1(_10832_),
    .A2(_10833_),
    .Y(_10834_),
    .B1(net5480));
 sg13g2_a22oi_1 _19223_ (.Y(_10835_),
    .B1(net5360),
    .B2(\atari2600.ram[127][6] ),
    .A2(net5407),
    .A1(\atari2600.ram[124][6] ));
 sg13g2_a22oi_1 _19224_ (.Y(_10836_),
    .B1(net5312),
    .B2(\atari2600.ram[126][6] ),
    .A2(net5452),
    .A1(\atari2600.ram[125][6] ));
 sg13g2_a21oi_2 _19225_ (.B1(net5488),
    .Y(_10837_),
    .A2(_10836_),
    .A1(_10835_));
 sg13g2_nor4_2 _19226_ (.A(_10828_),
    .B(_10831_),
    .C(_10834_),
    .Y(_10838_),
    .D(_10837_));
 sg13g2_nor2_2 _19227_ (.A(_09361_),
    .B(_10838_),
    .Y(_10839_));
 sg13g2_a22oi_1 _19228_ (.Y(_10840_),
    .B1(net5365),
    .B2(\atari2600.ram[111][6] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][6] ));
 sg13g2_a22oi_1 _19229_ (.Y(_10841_),
    .B1(net5319),
    .B2(\atari2600.ram[110][6] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][6] ));
 sg13g2_a21oi_2 _19230_ (.B1(net5494),
    .Y(_10842_),
    .A2(_10841_),
    .A1(_10840_));
 sg13g2_a22oi_1 _19231_ (.Y(_10843_),
    .B1(net5377),
    .B2(\atari2600.ram[99][6] ),
    .A2(net5425),
    .A1(\atari2600.ram[96][6] ));
 sg13g2_a22oi_1 _19232_ (.Y(_10844_),
    .B1(net5332),
    .B2(\atari2600.ram[98][6] ),
    .A2(net5471),
    .A1(\atari2600.ram[97][6] ));
 sg13g2_a21oi_1 _19233_ (.A1(_10843_),
    .A2(_10844_),
    .Y(_10845_),
    .B1(net5508));
 sg13g2_a22oi_1 _19234_ (.Y(_10846_),
    .B1(net5376),
    .B2(\atari2600.ram[107][6] ),
    .A2(net5424),
    .A1(\atari2600.ram[104][6] ));
 sg13g2_a22oi_1 _19235_ (.Y(_10847_),
    .B1(net5316),
    .B2(\atari2600.ram[106][6] ),
    .A2(net5455),
    .A1(\atari2600.ram[105][6] ));
 sg13g2_a21oi_1 _19236_ (.A1(_10846_),
    .A2(_10847_),
    .Y(_10848_),
    .B1(net5483));
 sg13g2_a22oi_1 _19237_ (.Y(_10849_),
    .B1(net5369),
    .B2(\atari2600.ram[103][6] ),
    .A2(net5416),
    .A1(\atari2600.ram[100][6] ));
 sg13g2_a22oi_1 _19238_ (.Y(_10850_),
    .B1(net5322),
    .B2(\atari2600.ram[102][6] ),
    .A2(net5461),
    .A1(\atari2600.ram[101][6] ));
 sg13g2_a21oi_1 _19239_ (.A1(_10849_),
    .A2(_10850_),
    .Y(_10851_),
    .B1(net5526));
 sg13g2_nor4_1 _19240_ (.A(_10842_),
    .B(_10845_),
    .C(_10848_),
    .D(_10851_),
    .Y(_10852_));
 sg13g2_a22oi_1 _19241_ (.Y(_10853_),
    .B1(net5377),
    .B2(\atari2600.ram[95][6] ),
    .A2(net5425),
    .A1(\atari2600.ram[92][6] ));
 sg13g2_a22oi_1 _19242_ (.Y(_10854_),
    .B1(net5333),
    .B2(\atari2600.ram[94][6] ),
    .A2(net5472),
    .A1(\atari2600.ram[93][6] ));
 sg13g2_a21oi_1 _19243_ (.A1(_10853_),
    .A2(_10854_),
    .Y(_10855_),
    .B1(net5498));
 sg13g2_a22oi_1 _19244_ (.Y(_10856_),
    .B1(net5382),
    .B2(\atari2600.ram[87][6] ),
    .A2(net5429),
    .A1(\atari2600.ram[84][6] ));
 sg13g2_a22oi_1 _19245_ (.Y(_10857_),
    .B1(net5335),
    .B2(\atari2600.ram[86][6] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][6] ));
 sg13g2_a21oi_1 _19246_ (.A1(_10856_),
    .A2(_10857_),
    .Y(_10858_),
    .B1(net5525));
 sg13g2_a22oi_1 _19247_ (.Y(_10859_),
    .B1(net5380),
    .B2(\atari2600.ram[91][6] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][6] ));
 sg13g2_a22oi_1 _19248_ (.Y(_10860_),
    .B1(net5334),
    .B2(\atari2600.ram[90][6] ),
    .A2(net5472),
    .A1(\atari2600.ram[89][6] ));
 sg13g2_a21oi_1 _19249_ (.A1(_10859_),
    .A2(_10860_),
    .Y(_10861_),
    .B1(net5486));
 sg13g2_a22oi_1 _19250_ (.Y(_10862_),
    .B1(net5375),
    .B2(\atari2600.ram[83][6] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][6] ));
 sg13g2_a22oi_1 _19251_ (.Y(_10863_),
    .B1(net5329),
    .B2(\atari2600.ram[82][6] ),
    .A2(net5469),
    .A1(\atari2600.ram[81][6] ));
 sg13g2_a21oi_1 _19252_ (.A1(_10862_),
    .A2(_10863_),
    .Y(_10864_),
    .B1(net5509));
 sg13g2_nor4_2 _19253_ (.A(_10855_),
    .B(_10858_),
    .C(_10861_),
    .Y(_10865_),
    .D(_10864_));
 sg13g2_nor2_1 _19254_ (.A(net5266),
    .B(_10865_),
    .Y(_10866_));
 sg13g2_a22oi_1 _19255_ (.Y(_10867_),
    .B1(net5368),
    .B2(\atari2600.ram[67][6] ),
    .A2(net5415),
    .A1(\atari2600.ram[64][6] ));
 sg13g2_a22oi_1 _19256_ (.Y(_10868_),
    .B1(net5324),
    .B2(\atari2600.ram[66][6] ),
    .A2(net5463),
    .A1(\atari2600.ram[65][6] ));
 sg13g2_a21oi_1 _19257_ (.A1(_10867_),
    .A2(_10868_),
    .Y(_10869_),
    .B1(net5511));
 sg13g2_a22oi_1 _19258_ (.Y(_10870_),
    .B1(net5378),
    .B2(\atari2600.ram[71][6] ),
    .A2(net5426),
    .A1(\atari2600.ram[68][6] ));
 sg13g2_a22oi_1 _19259_ (.Y(_10871_),
    .B1(net5331),
    .B2(\atari2600.ram[70][6] ),
    .A2(net5470),
    .A1(\atari2600.ram[69][6] ));
 sg13g2_a21oi_2 _19260_ (.B1(net5524),
    .Y(_10872_),
    .A2(_10871_),
    .A1(_10870_));
 sg13g2_a22oi_1 _19261_ (.Y(_10873_),
    .B1(net5370),
    .B2(\atari2600.ram[75][6] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][6] ));
 sg13g2_a22oi_1 _19262_ (.Y(_10874_),
    .B1(net5323),
    .B2(\atari2600.ram[74][6] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][6] ));
 sg13g2_a21oi_1 _19263_ (.A1(_10873_),
    .A2(_10874_),
    .Y(_10875_),
    .B1(net5485));
 sg13g2_a22oi_1 _19264_ (.Y(_10876_),
    .B1(net5367),
    .B2(\atari2600.ram[79][6] ),
    .A2(net5418),
    .A1(\atari2600.ram[76][6] ));
 sg13g2_a22oi_1 _19265_ (.Y(_10877_),
    .B1(net5320),
    .B2(\atari2600.ram[78][6] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][6] ));
 sg13g2_a21oi_2 _19266_ (.B1(net5496),
    .Y(_10878_),
    .A2(_10877_),
    .A1(_10876_));
 sg13g2_nor4_2 _19267_ (.A(_10869_),
    .B(_10872_),
    .C(_10875_),
    .Y(_10879_),
    .D(_10878_));
 sg13g2_nor2_1 _19268_ (.A(net5271),
    .B(_10879_),
    .Y(_10880_));
 sg13g2_o21ai_1 _19269_ (.B1(net5545),
    .Y(_10881_),
    .A1(net5269),
    .A2(_10852_));
 sg13g2_nor4_2 _19270_ (.A(_10839_),
    .B(_10866_),
    .C(_10880_),
    .Y(_10882_),
    .D(_10881_));
 sg13g2_a22oi_1 _19271_ (.Y(_10883_),
    .B1(net5392),
    .B2(\atari2600.ram[52][6] ),
    .A2(net5440),
    .A1(\atari2600.ram[53][6] ));
 sg13g2_a22oi_1 _19272_ (.Y(_10884_),
    .B1(net5300),
    .B2(\atari2600.ram[54][6] ),
    .A2(net5347),
    .A1(\atari2600.ram[55][6] ));
 sg13g2_a21oi_1 _19273_ (.A1(_10883_),
    .A2(_10884_),
    .Y(_10885_),
    .B1(net5518));
 sg13g2_a22oi_1 _19274_ (.Y(_10886_),
    .B1(net5347),
    .B2(\atari2600.ram[63][6] ),
    .A2(net5392),
    .A1(\atari2600.ram[60][6] ));
 sg13g2_a22oi_1 _19275_ (.Y(_10887_),
    .B1(net5301),
    .B2(\atari2600.ram[62][6] ),
    .A2(net5441),
    .A1(\atari2600.ram[61][6] ));
 sg13g2_a21oi_1 _19276_ (.A1(_10886_),
    .A2(_10887_),
    .Y(_10888_),
    .B1(net5488));
 sg13g2_a22oi_1 _19277_ (.Y(_10889_),
    .B1(net5350),
    .B2(\atari2600.ram[59][6] ),
    .A2(net5395),
    .A1(\atari2600.ram[56][6] ));
 sg13g2_a22oi_1 _19278_ (.Y(_10890_),
    .B1(net5304),
    .B2(\atari2600.ram[58][6] ),
    .A2(net5444),
    .A1(\atari2600.ram[57][6] ));
 sg13g2_a21oi_2 _19279_ (.B1(net5480),
    .Y(_10891_),
    .A2(_10890_),
    .A1(_10889_));
 sg13g2_a22oi_1 _19280_ (.Y(_10892_),
    .B1(net5342),
    .B2(\atari2600.ram[51][6] ),
    .A2(net5391),
    .A1(\atari2600.ram[48][6] ));
 sg13g2_a22oi_1 _19281_ (.Y(_10893_),
    .B1(net5299),
    .B2(\atari2600.ram[50][6] ),
    .A2(net5439),
    .A1(\atari2600.ram[49][6] ));
 sg13g2_a21o_1 _19282_ (.A2(_10893_),
    .A1(_10892_),
    .B1(net5501),
    .X(_10894_));
 sg13g2_nor4_2 _19283_ (.A(net5281),
    .B(_10885_),
    .C(_10888_),
    .Y(_10895_),
    .D(_10891_));
 sg13g2_a22oi_1 _19284_ (.Y(_10896_),
    .B1(net5342),
    .B2(\atari2600.ram[47][6] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][6] ));
 sg13g2_a22oi_1 _19285_ (.Y(_10897_),
    .B1(net5295),
    .B2(\atari2600.ram[46][6] ),
    .A2(net5435),
    .A1(\atari2600.ram[45][6] ));
 sg13g2_a21oi_1 _19286_ (.A1(_10896_),
    .A2(_10897_),
    .Y(_10898_),
    .B1(net5490));
 sg13g2_a22oi_1 _19287_ (.Y(_10899_),
    .B1(net5343),
    .B2(\atari2600.ram[35][6] ),
    .A2(net5387),
    .A1(\atari2600.ram[32][6] ));
 sg13g2_a22oi_1 _19288_ (.Y(_10900_),
    .B1(net5295),
    .B2(\atari2600.ram[34][6] ),
    .A2(net5435),
    .A1(\atari2600.ram[33][6] ));
 sg13g2_a21oi_1 _19289_ (.A1(_10899_),
    .A2(_10900_),
    .Y(_10901_),
    .B1(net5502));
 sg13g2_a22oi_1 _19290_ (.Y(_10902_),
    .B1(net5390),
    .B2(\atari2600.ram[40][6] ),
    .A2(net5436),
    .A1(\atari2600.ram[41][6] ));
 sg13g2_a22oi_1 _19291_ (.Y(_10903_),
    .B1(net5296),
    .B2(\atari2600.ram[42][6] ),
    .A2(net5345),
    .A1(\atari2600.ram[43][6] ));
 sg13g2_a21oi_1 _19292_ (.A1(_10902_),
    .A2(_10903_),
    .Y(_10904_),
    .B1(net5477));
 sg13g2_a22oi_1 _19293_ (.Y(_10905_),
    .B1(net5340),
    .B2(\atari2600.ram[39][6] ),
    .A2(net5385),
    .A1(\atari2600.ram[36][6] ));
 sg13g2_a22oi_1 _19294_ (.Y(_10906_),
    .B1(net5293),
    .B2(\atari2600.ram[38][6] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][6] ));
 sg13g2_a21oi_2 _19295_ (.B1(net5515),
    .Y(_10907_),
    .A2(_10906_),
    .A1(_10905_));
 sg13g2_nor2_1 _19296_ (.A(net5275),
    .B(_10901_),
    .Y(_10908_));
 sg13g2_nor3_1 _19297_ (.A(_10898_),
    .B(_10904_),
    .C(_10907_),
    .Y(_10909_));
 sg13g2_a221oi_1 _19298_ (.B2(_10909_),
    .C1(net5568),
    .B1(_10908_),
    .A1(_10894_),
    .Y(_10910_),
    .A2(_10895_));
 sg13g2_a22oi_1 _19299_ (.Y(_10911_),
    .B1(net5373),
    .B2(\atari2600.ram[31][6] ),
    .A2(net5421),
    .A1(\atari2600.ram[28][6] ));
 sg13g2_a22oi_1 _19300_ (.Y(_10912_),
    .B1(net5328),
    .B2(\atari2600.ram[30][6] ),
    .A2(net5467),
    .A1(\atari2600.ram[29][6] ));
 sg13g2_a21oi_2 _19301_ (.B1(net5492),
    .Y(_10913_),
    .A2(_10912_),
    .A1(_10911_));
 sg13g2_a22oi_1 _19302_ (.Y(_10914_),
    .B1(net5356),
    .B2(\atari2600.ram[19][6] ),
    .A2(net5403),
    .A1(\atari2600.ram[16][6] ));
 sg13g2_a22oi_1 _19303_ (.Y(_10915_),
    .B1(net5310),
    .B2(\atari2600.ram[18][6] ),
    .A2(net5449),
    .A1(\atari2600.ram[17][6] ));
 sg13g2_a21oi_2 _19304_ (.B1(net5504),
    .Y(_10916_),
    .A2(_10915_),
    .A1(_10914_));
 sg13g2_a22oi_1 _19305_ (.Y(_10917_),
    .B1(net5356),
    .B2(\atari2600.ram[23][6] ),
    .A2(net5402),
    .A1(\atari2600.ram[20][6] ));
 sg13g2_a22oi_1 _19306_ (.Y(_10918_),
    .B1(net5310),
    .B2(\atari2600.ram[22][6] ),
    .A2(net5449),
    .A1(\atari2600.ram[21][6] ));
 sg13g2_a21oi_1 _19307_ (.A1(_10917_),
    .A2(_10918_),
    .Y(_10919_),
    .B1(net5517));
 sg13g2_a22oi_1 _19308_ (.Y(_10920_),
    .B1(net5355),
    .B2(\atari2600.ram[7][6] ),
    .A2(net5401),
    .A1(\atari2600.ram[4][6] ));
 sg13g2_a22oi_1 _19309_ (.Y(_10921_),
    .B1(net5311),
    .B2(\atari2600.ram[6][6] ),
    .A2(net5451),
    .A1(\atari2600.ram[5][6] ));
 sg13g2_a21oi_2 _19310_ (.B1(net5516),
    .Y(_10922_),
    .A2(_10921_),
    .A1(_10920_));
 sg13g2_a22oi_1 _19311_ (.Y(_10923_),
    .B1(net5353),
    .B2(\atari2600.ram[3][6] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][6] ));
 sg13g2_a22oi_1 _19312_ (.Y(_10924_),
    .B1(net5307),
    .B2(\atari2600.ram[2][6] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][6] ));
 sg13g2_a21oi_1 _19313_ (.A1(_10923_),
    .A2(_10924_),
    .Y(_10925_),
    .B1(net5503));
 sg13g2_a22oi_1 _19314_ (.Y(_10926_),
    .B1(net5344),
    .B2(\atari2600.ram[11][6] ),
    .A2(net5389),
    .A1(\atari2600.ram[8][6] ));
 sg13g2_a22oi_1 _19315_ (.Y(_10927_),
    .B1(net5297),
    .B2(\atari2600.ram[10][6] ),
    .A2(net5437),
    .A1(\atari2600.ram[9][6] ));
 sg13g2_a21oi_2 _19316_ (.B1(net5477),
    .Y(_10928_),
    .A2(_10927_),
    .A1(_10926_));
 sg13g2_a22oi_1 _19317_ (.Y(_10929_),
    .B1(net5355),
    .B2(\atari2600.ram[15][6] ),
    .A2(net5399),
    .A1(\atari2600.ram[12][6] ));
 sg13g2_a22oi_1 _19318_ (.Y(_10930_),
    .B1(net5306),
    .B2(\atari2600.ram[14][6] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][6] ));
 sg13g2_a21oi_1 _19319_ (.A1(_10929_),
    .A2(_10930_),
    .Y(_10931_),
    .B1(net5491));
 sg13g2_nor4_2 _19320_ (.A(_10922_),
    .B(_10925_),
    .C(_10928_),
    .Y(_10932_),
    .D(_10931_));
 sg13g2_nor2_1 _19321_ (.A(net5270),
    .B(_10932_),
    .Y(_10933_));
 sg13g2_a22oi_1 _19322_ (.Y(_10934_),
    .B1(net5371),
    .B2(\atari2600.ram[27][6] ),
    .A2(net5419),
    .A1(\atari2600.ram[24][6] ));
 sg13g2_a22oi_1 _19323_ (.Y(_10935_),
    .B1(net5326),
    .B2(\atari2600.ram[26][6] ),
    .A2(net5465),
    .A1(\atari2600.ram[25][6] ));
 sg13g2_a21oi_2 _19324_ (.B1(net5482),
    .Y(_10936_),
    .A2(_10935_),
    .A1(_10934_));
 sg13g2_nor4_2 _19325_ (.A(_10913_),
    .B(_10916_),
    .C(_10919_),
    .Y(_10937_),
    .D(_10936_));
 sg13g2_nor2_2 _19326_ (.A(net5264),
    .B(_10937_),
    .Y(_10938_));
 sg13g2_nor4_1 _19327_ (.A(net5544),
    .B(_10910_),
    .C(_10933_),
    .D(_10938_),
    .Y(_10939_));
 sg13g2_nor2_1 _19328_ (.A(_10882_),
    .B(_10939_),
    .Y(_00007_));
 sg13g2_a22oi_1 _19329_ (.Y(_10940_),
    .B1(net5394),
    .B2(\atari2600.ram[56][7] ),
    .A2(net5443),
    .A1(\atari2600.ram[57][7] ));
 sg13g2_a22oi_1 _19330_ (.Y(_10941_),
    .B1(net5303),
    .B2(\atari2600.ram[58][7] ),
    .A2(net5349),
    .A1(\atari2600.ram[59][7] ));
 sg13g2_a21oi_1 _19331_ (.A1(_10940_),
    .A2(_10941_),
    .Y(_10942_),
    .B1(net5478));
 sg13g2_a22oi_1 _19332_ (.Y(_10943_),
    .B1(net5347),
    .B2(\atari2600.ram[63][7] ),
    .A2(net5392),
    .A1(\atari2600.ram[60][7] ));
 sg13g2_a22oi_1 _19333_ (.Y(_10944_),
    .B1(net5300),
    .B2(\atari2600.ram[62][7] ),
    .A2(net5440),
    .A1(\atari2600.ram[61][7] ));
 sg13g2_a21oi_1 _19334_ (.A1(_10943_),
    .A2(_10944_),
    .Y(_10945_),
    .B1(net5488));
 sg13g2_a22oi_1 _19335_ (.Y(_10946_),
    .B1(net5346),
    .B2(\atari2600.ram[55][7] ),
    .A2(net5391),
    .A1(\atari2600.ram[52][7] ));
 sg13g2_a22oi_1 _19336_ (.Y(_10947_),
    .B1(net5298),
    .B2(\atari2600.ram[54][7] ),
    .A2(net5438),
    .A1(\atari2600.ram[53][7] ));
 sg13g2_a21oi_1 _19337_ (.A1(_10946_),
    .A2(_10947_),
    .Y(_10948_),
    .B1(net5518));
 sg13g2_a22oi_1 _19338_ (.Y(_10949_),
    .B1(net5349),
    .B2(\atari2600.ram[51][7] ),
    .A2(net5394),
    .A1(\atari2600.ram[48][7] ));
 sg13g2_a22oi_1 _19339_ (.Y(_10950_),
    .B1(net5303),
    .B2(\atari2600.ram[50][7] ),
    .A2(net5443),
    .A1(\atari2600.ram[49][7] ));
 sg13g2_a21o_1 _19340_ (.A2(_10950_),
    .A1(_10949_),
    .B1(net5501),
    .X(_10951_));
 sg13g2_nor4_1 _19341_ (.A(net5280),
    .B(_10942_),
    .C(_10945_),
    .D(_10948_),
    .Y(_10952_));
 sg13g2_a22oi_1 _19342_ (.Y(_10953_),
    .B1(net5385),
    .B2(\atari2600.ram[36][7] ),
    .A2(net5433),
    .A1(\atari2600.ram[37][7] ));
 sg13g2_a22oi_1 _19343_ (.Y(_10954_),
    .B1(net5293),
    .B2(\atari2600.ram[38][7] ),
    .A2(net5340),
    .A1(\atari2600.ram[39][7] ));
 sg13g2_a21oi_1 _19344_ (.A1(_10953_),
    .A2(_10954_),
    .Y(_10955_),
    .B1(net5515));
 sg13g2_a22oi_1 _19345_ (.Y(_10956_),
    .B1(net5341),
    .B2(\atari2600.ram[35][7] ),
    .A2(net5385),
    .A1(\atari2600.ram[32][7] ));
 sg13g2_a22oi_1 _19346_ (.Y(_10957_),
    .B1(net5294),
    .B2(\atari2600.ram[34][7] ),
    .A2(net5434),
    .A1(\atari2600.ram[33][7] ));
 sg13g2_a21oi_1 _19347_ (.A1(_10956_),
    .A2(_10957_),
    .Y(_10958_),
    .B1(net5501));
 sg13g2_a22oi_1 _19348_ (.Y(_10959_),
    .B1(net5345),
    .B2(\atari2600.ram[43][7] ),
    .A2(net5390),
    .A1(\atari2600.ram[40][7] ));
 sg13g2_a22oi_1 _19349_ (.Y(_10960_),
    .B1(net5296),
    .B2(\atari2600.ram[42][7] ),
    .A2(net5436),
    .A1(\atari2600.ram[41][7] ));
 sg13g2_a21oi_1 _19350_ (.A1(_10959_),
    .A2(_10960_),
    .Y(_10961_),
    .B1(net5479));
 sg13g2_a22oi_1 _19351_ (.Y(_10962_),
    .B1(net5340),
    .B2(\atari2600.ram[47][7] ),
    .A2(net5387),
    .A1(\atari2600.ram[44][7] ));
 sg13g2_a22oi_1 _19352_ (.Y(_10963_),
    .B1(net5293),
    .B2(\atari2600.ram[46][7] ),
    .A2(net5433),
    .A1(\atari2600.ram[45][7] ));
 sg13g2_a21oi_1 _19353_ (.A1(_10962_),
    .A2(_10963_),
    .Y(_10964_),
    .B1(net5490));
 sg13g2_nor2_1 _19354_ (.A(net5275),
    .B(_10961_),
    .Y(_10965_));
 sg13g2_nor3_2 _19355_ (.A(_10955_),
    .B(_10958_),
    .C(_10964_),
    .Y(_10966_));
 sg13g2_a221oi_1 _19356_ (.B2(_10966_),
    .C1(net5568),
    .B1(_10965_),
    .A1(_10951_),
    .Y(_10967_),
    .A2(_10952_));
 sg13g2_a22oi_1 _19357_ (.Y(_10968_),
    .B1(net5373),
    .B2(\atari2600.ram[31][7] ),
    .A2(net5421),
    .A1(\atari2600.ram[28][7] ));
 sg13g2_a22oi_1 _19358_ (.Y(_10969_),
    .B1(net5328),
    .B2(\atari2600.ram[30][7] ),
    .A2(net5467),
    .A1(\atari2600.ram[29][7] ));
 sg13g2_a21oi_2 _19359_ (.B1(net5492),
    .Y(_10970_),
    .A2(_10969_),
    .A1(_10968_));
 sg13g2_a22oi_1 _19360_ (.Y(_10971_),
    .B1(net5371),
    .B2(\atari2600.ram[23][7] ),
    .A2(net5419),
    .A1(\atari2600.ram[20][7] ));
 sg13g2_a22oi_1 _19361_ (.Y(_10972_),
    .B1(net5326),
    .B2(\atari2600.ram[22][7] ),
    .A2(net5465),
    .A1(\atari2600.ram[21][7] ));
 sg13g2_a21oi_1 _19362_ (.A1(_10971_),
    .A2(_10972_),
    .Y(_10973_),
    .B1(net5522));
 sg13g2_a22oi_1 _19363_ (.Y(_10974_),
    .B1(net5372),
    .B2(\atari2600.ram[27][7] ),
    .A2(net5420),
    .A1(\atari2600.ram[24][7] ));
 sg13g2_a22oi_1 _19364_ (.Y(_10975_),
    .B1(net5327),
    .B2(\atari2600.ram[26][7] ),
    .A2(net5466),
    .A1(\atari2600.ram[25][7] ));
 sg13g2_a21oi_1 _19365_ (.A1(_10974_),
    .A2(_10975_),
    .Y(_10976_),
    .B1(net5482));
 sg13g2_a22oi_1 _19366_ (.Y(_10977_),
    .B1(net5373),
    .B2(\atari2600.ram[19][7] ),
    .A2(net5421),
    .A1(\atari2600.ram[16][7] ));
 sg13g2_a22oi_1 _19367_ (.Y(_10978_),
    .B1(net5328),
    .B2(\atari2600.ram[18][7] ),
    .A2(net5467),
    .A1(\atari2600.ram[17][7] ));
 sg13g2_a21oi_2 _19368_ (.B1(net5509),
    .Y(_10979_),
    .A2(_10978_),
    .A1(_10977_));
 sg13g2_nor4_2 _19369_ (.A(_10970_),
    .B(_10973_),
    .C(_10976_),
    .Y(_10980_),
    .D(_10979_));
 sg13g2_nor2_2 _19370_ (.A(net5265),
    .B(_10980_),
    .Y(_10981_));
 sg13g2_a22oi_1 _19371_ (.Y(_10982_),
    .B1(net5344),
    .B2(\atari2600.ram[11][7] ),
    .A2(net5389),
    .A1(\atari2600.ram[8][7] ));
 sg13g2_a22oi_1 _19372_ (.Y(_10983_),
    .B1(net5296),
    .B2(\atari2600.ram[10][7] ),
    .A2(net5437),
    .A1(\atari2600.ram[9][7] ));
 sg13g2_a21oi_2 _19373_ (.B1(net5478),
    .Y(_10984_),
    .A2(_10983_),
    .A1(_10982_));
 sg13g2_a22oi_1 _19374_ (.Y(_10985_),
    .B1(net5355),
    .B2(\atari2600.ram[7][7] ),
    .A2(net5401),
    .A1(\atari2600.ram[4][7] ));
 sg13g2_a22oi_1 _19375_ (.Y(_10986_),
    .B1(net5308),
    .B2(\atari2600.ram[6][7] ),
    .A2(net5448),
    .A1(\atari2600.ram[5][7] ));
 sg13g2_a21oi_2 _19376_ (.B1(net5516),
    .Y(_10987_),
    .A2(_10986_),
    .A1(_10985_));
 sg13g2_a22oi_1 _19377_ (.Y(_10988_),
    .B1(net5353),
    .B2(\atari2600.ram[3][7] ),
    .A2(net5398),
    .A1(\atari2600.ram[0][7] ));
 sg13g2_a22oi_1 _19378_ (.Y(_10989_),
    .B1(net5307),
    .B2(\atari2600.ram[2][7] ),
    .A2(net5447),
    .A1(\atari2600.ram[1][7] ));
 sg13g2_a21oi_1 _19379_ (.A1(_10988_),
    .A2(_10989_),
    .Y(_10990_),
    .B1(net5503));
 sg13g2_a22oi_1 _19380_ (.Y(_10991_),
    .B1(net5354),
    .B2(\atari2600.ram[15][7] ),
    .A2(net5399),
    .A1(\atari2600.ram[12][7] ));
 sg13g2_a22oi_1 _19381_ (.Y(_10992_),
    .B1(net5306),
    .B2(\atari2600.ram[14][7] ),
    .A2(net5446),
    .A1(\atari2600.ram[13][7] ));
 sg13g2_a21oi_1 _19382_ (.A1(_10991_),
    .A2(_10992_),
    .Y(_10993_),
    .B1(net5491));
 sg13g2_nor4_2 _19383_ (.A(_10984_),
    .B(_10987_),
    .C(_10990_),
    .Y(_10994_),
    .D(_10993_));
 sg13g2_o21ai_1 _19384_ (.B1(net5543),
    .Y(_10995_),
    .A1(net5270),
    .A2(_10994_));
 sg13g2_nor3_1 _19385_ (.A(_10967_),
    .B(_10981_),
    .C(_10995_),
    .Y(_10996_));
 sg13g2_a22oi_1 _19386_ (.Y(_10997_),
    .B1(net5372),
    .B2(\atari2600.ram[107][7] ),
    .A2(net5420),
    .A1(\atari2600.ram[104][7] ));
 sg13g2_a22oi_1 _19387_ (.Y(_10998_),
    .B1(net5325),
    .B2(\atari2600.ram[106][7] ),
    .A2(net5464),
    .A1(\atari2600.ram[105][7] ));
 sg13g2_a21oi_1 _19388_ (.A1(_10997_),
    .A2(_10998_),
    .Y(_10999_),
    .B1(net5483));
 sg13g2_a22oi_1 _19389_ (.Y(_11000_),
    .B1(net5366),
    .B2(\atari2600.ram[103][7] ),
    .A2(net5413),
    .A1(\atari2600.ram[100][7] ));
 sg13g2_a22oi_1 _19390_ (.Y(_11001_),
    .B1(net5322),
    .B2(\atari2600.ram[102][7] ),
    .A2(net5461),
    .A1(\atari2600.ram[101][7] ));
 sg13g2_a21oi_2 _19391_ (.B1(net5526),
    .Y(_11002_),
    .A2(_11001_),
    .A1(_11000_));
 sg13g2_a22oi_1 _19392_ (.Y(_11003_),
    .B1(net5377),
    .B2(\atari2600.ram[99][7] ),
    .A2(net5425),
    .A1(\atari2600.ram[96][7] ));
 sg13g2_a22oi_1 _19393_ (.Y(_11004_),
    .B1(net5332),
    .B2(\atari2600.ram[98][7] ),
    .A2(net5471),
    .A1(\atari2600.ram[97][7] ));
 sg13g2_a21oi_1 _19394_ (.A1(_11003_),
    .A2(_11004_),
    .Y(_11005_),
    .B1(net5511));
 sg13g2_a22oi_1 _19395_ (.Y(_11006_),
    .B1(net5365),
    .B2(\atari2600.ram[111][7] ),
    .A2(net5412),
    .A1(\atari2600.ram[108][7] ));
 sg13g2_a22oi_1 _19396_ (.Y(_11007_),
    .B1(net5319),
    .B2(\atari2600.ram[110][7] ),
    .A2(net5458),
    .A1(\atari2600.ram[109][7] ));
 sg13g2_a21oi_2 _19397_ (.B1(net5494),
    .Y(_11008_),
    .A2(_11007_),
    .A1(_11006_));
 sg13g2_nor4_1 _19398_ (.A(_10999_),
    .B(_11002_),
    .C(_11005_),
    .D(_11008_),
    .Y(_11009_));
 sg13g2_nor2_1 _19399_ (.A(net5269),
    .B(_11009_),
    .Y(_11010_));
 sg13g2_a22oi_1 _19400_ (.Y(_11011_),
    .B1(net5367),
    .B2(\atari2600.ram[79][7] ),
    .A2(net5414),
    .A1(\atari2600.ram[76][7] ));
 sg13g2_a22oi_1 _19401_ (.Y(_11012_),
    .B1(net5320),
    .B2(\atari2600.ram[78][7] ),
    .A2(net5459),
    .A1(\atari2600.ram[77][7] ));
 sg13g2_a21oi_2 _19402_ (.B1(net5496),
    .Y(_11013_),
    .A2(_11012_),
    .A1(_11011_));
 sg13g2_a22oi_1 _19403_ (.Y(_11014_),
    .B1(net5368),
    .B2(\atari2600.ram[67][7] ),
    .A2(net5417),
    .A1(\atari2600.ram[64][7] ));
 sg13g2_a22oi_1 _19404_ (.Y(_11015_),
    .B1(net5324),
    .B2(\atari2600.ram[66][7] ),
    .A2(net5463),
    .A1(\atari2600.ram[65][7] ));
 sg13g2_a21oi_1 _19405_ (.A1(_11014_),
    .A2(_11015_),
    .Y(_11016_),
    .B1(net5511));
 sg13g2_a22oi_1 _19406_ (.Y(_11017_),
    .B1(net5368),
    .B2(\atari2600.ram[75][7] ),
    .A2(net5415),
    .A1(\atari2600.ram[72][7] ));
 sg13g2_a22oi_1 _19407_ (.Y(_11018_),
    .B1(net5323),
    .B2(\atari2600.ram[74][7] ),
    .A2(net5462),
    .A1(\atari2600.ram[73][7] ));
 sg13g2_a21oi_1 _19408_ (.A1(_11017_),
    .A2(_11018_),
    .Y(_11019_),
    .B1(net5485));
 sg13g2_a22oi_1 _19409_ (.Y(_11020_),
    .B1(net5378),
    .B2(\atari2600.ram[71][7] ),
    .A2(net5426),
    .A1(\atari2600.ram[68][7] ));
 sg13g2_a22oi_1 _19410_ (.Y(_11021_),
    .B1(net5331),
    .B2(\atari2600.ram[70][7] ),
    .A2(net5470),
    .A1(\atari2600.ram[69][7] ));
 sg13g2_a21oi_2 _19411_ (.B1(net5524),
    .Y(_11022_),
    .A2(_11021_),
    .A1(_11020_));
 sg13g2_nor4_2 _19412_ (.A(_11013_),
    .B(_11016_),
    .C(_11019_),
    .Y(_11023_),
    .D(_11022_));
 sg13g2_nor2_1 _19413_ (.A(net5271),
    .B(_11023_),
    .Y(_11024_));
 sg13g2_a22oi_1 _19414_ (.Y(_11025_),
    .B1(net5377),
    .B2(\atari2600.ram[95][7] ),
    .A2(net5425),
    .A1(\atari2600.ram[92][7] ));
 sg13g2_a22oi_1 _19415_ (.Y(_11026_),
    .B1(net5332),
    .B2(\atari2600.ram[94][7] ),
    .A2(net5471),
    .A1(\atari2600.ram[93][7] ));
 sg13g2_a21oi_1 _19416_ (.A1(_11025_),
    .A2(_11026_),
    .Y(_11027_),
    .B1(net5498));
 sg13g2_a22oi_1 _19417_ (.Y(_11028_),
    .B1(net5375),
    .B2(\atari2600.ram[83][7] ),
    .A2(net5422),
    .A1(\atari2600.ram[80][7] ));
 sg13g2_a22oi_1 _19418_ (.Y(_11029_),
    .B1(net5329),
    .B2(\atari2600.ram[82][7] ),
    .A2(net5469),
    .A1(\atari2600.ram[81][7] ));
 sg13g2_a21oi_2 _19419_ (.B1(net5508),
    .Y(_11030_),
    .A2(_11029_),
    .A1(_11028_));
 sg13g2_a22oi_1 _19420_ (.Y(_11031_),
    .B1(net5382),
    .B2(\atari2600.ram[87][7] ),
    .A2(net5430),
    .A1(\atari2600.ram[84][7] ));
 sg13g2_a22oi_1 _19421_ (.Y(_11032_),
    .B1(net5335),
    .B2(\atari2600.ram[86][7] ),
    .A2(net5474),
    .A1(\atari2600.ram[85][7] ));
 sg13g2_a21oi_1 _19422_ (.A1(_11031_),
    .A2(_11032_),
    .Y(_11033_),
    .B1(net5524));
 sg13g2_a22oi_1 _19423_ (.Y(_11034_),
    .B1(net5380),
    .B2(\atari2600.ram[91][7] ),
    .A2(net5428),
    .A1(\atari2600.ram[88][7] ));
 sg13g2_a22oi_1 _19424_ (.Y(_11035_),
    .B1(net5333),
    .B2(\atari2600.ram[90][7] ),
    .A2(net5472),
    .A1(\atari2600.ram[89][7] ));
 sg13g2_a21oi_1 _19425_ (.A1(_11034_),
    .A2(_11035_),
    .Y(_11036_),
    .B1(net5486));
 sg13g2_nor4_2 _19426_ (.A(_11027_),
    .B(_11030_),
    .C(_11033_),
    .Y(_11037_),
    .D(_11036_));
 sg13g2_a22oi_1 _19427_ (.Y(_11038_),
    .B1(net5360),
    .B2(\atari2600.ram[127][7] ),
    .A2(net5407),
    .A1(\atari2600.ram[124][7] ));
 sg13g2_a22oi_1 _19428_ (.Y(_11039_),
    .B1(net5312),
    .B2(\atari2600.ram[126][7] ),
    .A2(net5452),
    .A1(\atari2600.ram[125][7] ));
 sg13g2_a21oi_2 _19429_ (.B1(net5488),
    .Y(_11040_),
    .A2(_11039_),
    .A1(_11038_));
 sg13g2_a22oi_1 _19430_ (.Y(_11041_),
    .B1(net5360),
    .B2(\atari2600.ram[119][7] ),
    .A2(net5407),
    .A1(\atari2600.ram[116][7] ));
 sg13g2_a22oi_1 _19431_ (.Y(_11042_),
    .B1(net5313),
    .B2(\atari2600.ram[118][7] ),
    .A2(net5454),
    .A1(\atari2600.ram[117][7] ));
 sg13g2_a21oi_1 _19432_ (.A1(_11041_),
    .A2(_11042_),
    .Y(_11043_),
    .B1(net5520));
 sg13g2_a22oi_1 _19433_ (.Y(_11044_),
    .B1(net5362),
    .B2(\atari2600.ram[115][7] ),
    .A2(net5408),
    .A1(\atari2600.ram[112][7] ));
 sg13g2_a22oi_1 _19434_ (.Y(_11045_),
    .B1(net5313),
    .B2(\atari2600.ram[114][7] ),
    .A2(net5454),
    .A1(\atari2600.ram[113][7] ));
 sg13g2_a21oi_1 _19435_ (.A1(_11044_),
    .A2(_11045_),
    .Y(_11046_),
    .B1(net5506));
 sg13g2_a22oi_1 _19436_ (.Y(_11047_),
    .B1(net5350),
    .B2(\atari2600.ram[123][7] ),
    .A2(net5395),
    .A1(\atari2600.ram[120][7] ));
 sg13g2_a22oi_1 _19437_ (.Y(_11048_),
    .B1(net5317),
    .B2(\atari2600.ram[122][7] ),
    .A2(net5456),
    .A1(\atari2600.ram[121][7] ));
 sg13g2_a21oi_2 _19438_ (.B1(net5481),
    .Y(_11049_),
    .A2(_11048_),
    .A1(_11047_));
 sg13g2_nor4_2 _19439_ (.A(_11040_),
    .B(_11043_),
    .C(_11046_),
    .Y(_11050_),
    .D(_11049_));
 sg13g2_nor2_2 _19440_ (.A(_09361_),
    .B(_11050_),
    .Y(_11051_));
 sg13g2_o21ai_1 _19441_ (.B1(net5545),
    .Y(_11052_),
    .A1(net5266),
    .A2(_11037_));
 sg13g2_nor4_2 _19442_ (.A(_11010_),
    .B(_11024_),
    .C(_11051_),
    .Y(_11053_),
    .D(_11052_));
 sg13g2_nor2_1 _19443_ (.A(_10996_),
    .B(_11053_),
    .Y(_00008_));
 sg13g2_nand2_2 _19444_ (.Y(_11054_),
    .A(\flash_rom.fsm_state[1] ),
    .B(_08473_));
 sg13g2_nor2_2 _19445_ (.A(net6245),
    .B(_11054_),
    .Y(_11055_));
 sg13g2_nor2_2 _19446_ (.A(\flash_rom.fsm_state[1] ),
    .B(_08473_),
    .Y(_11056_));
 sg13g2_nand2_1 _19447_ (.Y(_11057_),
    .A(net7303),
    .B(_11056_));
 sg13g2_o21ai_1 _19448_ (.B1(net7444),
    .Y(_11058_),
    .A1(\flash_rom.nibbles_remaining[1] ),
    .A2(\flash_rom.nibbles_remaining[0] ));
 sg13g2_a21oi_1 _19449_ (.A1(\flash_rom.nibbles_remaining[1] ),
    .A2(_08474_),
    .Y(_11059_),
    .B1(\flash_rom.nibbles_remaining[2] ));
 sg13g2_nor2_1 _19450_ (.A(_11057_),
    .B(_11059_),
    .Y(_11060_));
 sg13g2_a22oi_1 _19451_ (.Y(uio_out[1]),
    .B1(_11058_),
    .B2(_11060_),
    .A2(_11055_),
    .A1(_08558_));
 sg13g2_and2_1 _19452_ (.A(\flash_rom.addr[21] ),
    .B(_11055_),
    .X(uio_out[2]));
 sg13g2_and2_1 _19453_ (.A(\flash_rom.addr[22] ),
    .B(_11055_),
    .X(uio_out[4]));
 sg13g2_and2_1 _19454_ (.A(\flash_rom.addr[23] ),
    .B(_11055_),
    .X(uio_out[5]));
 sg13g2_nand2_1 _19455_ (.Y(_00172_),
    .A(_08948_),
    .B(_08988_));
 sg13g2_nand4_1 _19456_ (.B(_08956_),
    .C(_08973_),
    .A(_08953_),
    .Y(_11061_),
    .D(_08979_));
 sg13g2_or4_1 _19457_ (.A(_08934_),
    .B(_09001_),
    .C(_09037_),
    .D(_11061_),
    .X(_00173_));
 sg13g2_nor4_1 _19458_ (.A(_08794_),
    .B(_08882_),
    .C(_08952_),
    .D(_08972_),
    .Y(_11062_));
 sg13g2_nand4_1 _19459_ (.B(_08998_),
    .C(_09028_),
    .A(_08964_),
    .Y(_11063_),
    .D(_11062_));
 sg13g2_nor4_1 _19460_ (.A(_08857_),
    .B(_08868_),
    .C(_08982_),
    .D(_11063_),
    .Y(_11064_));
 sg13g2_nor2_1 _19461_ (.A(_08938_),
    .B(_09009_),
    .Y(_11065_));
 sg13g2_nand4_1 _19462_ (.B(_08899_),
    .C(_11064_),
    .A(_08889_),
    .Y(_11066_),
    .D(_11065_));
 sg13g2_a221oi_1 _19463_ (.B2(net5823),
    .C1(_11066_),
    .B1(_08766_),
    .A1(_08721_),
    .Y(_11067_),
    .A2(net5851));
 sg13g2_nand2_1 _19464_ (.Y(_00174_),
    .A(_08912_),
    .B(_11067_));
 sg13g2_nand2b_1 _19465_ (.Y(_11068_),
    .B(_09030_),
    .A_N(_08791_));
 sg13g2_nor3_1 _19466_ (.A(_08865_),
    .B(_08970_),
    .C(_11068_),
    .Y(_11069_));
 sg13g2_nor2_1 _19467_ (.A(_08860_),
    .B(_08984_),
    .Y(_11070_));
 sg13g2_nand4_1 _19468_ (.B(_09014_),
    .C(_11069_),
    .A(_08960_),
    .Y(_11071_),
    .D(_11070_));
 sg13g2_nand2_1 _19469_ (.Y(_11072_),
    .A(_08916_),
    .B(_08942_));
 sg13g2_nor4_1 _19470_ (.A(_08782_),
    .B(_08893_),
    .C(_11071_),
    .D(_11072_),
    .Y(_11073_));
 sg13g2_nand4_1 _19471_ (.B(_08901_),
    .C(_09006_),
    .A(_08842_),
    .Y(_11074_),
    .D(_11073_));
 sg13g2_nor3_1 _19472_ (.A(_08950_),
    .B(_08955_),
    .C(_11074_),
    .Y(_11075_));
 sg13g2_nand2_1 _19473_ (.Y(_00175_),
    .A(_08996_),
    .B(_11075_));
 sg13g2_and2_1 _19474_ (.A(net4937),
    .B(\atari2600.cpu.adc_sbc ),
    .X(_00022_));
 sg13g2_xor2_1 _19475_ (.B(net8),
    .A(net1),
    .X(_11076_));
 sg13g2_mux2_1 _19476_ (.A0(net2994),
    .A1(_11076_),
    .S(net6523),
    .X(_00177_));
 sg13g2_xor2_1 _19477_ (.B(net8),
    .A(net2),
    .X(_11077_));
 sg13g2_mux2_1 _19478_ (.A0(net4517),
    .A1(_11077_),
    .S(net6523),
    .X(_00178_));
 sg13g2_xor2_1 _19479_ (.B(net8),
    .A(net3),
    .X(_11078_));
 sg13g2_mux2_1 _19480_ (.A0(net7194),
    .A1(_11078_),
    .S(net6522),
    .X(_00179_));
 sg13g2_or2_1 _19481_ (.X(_11079_),
    .B(net8),
    .A(net4));
 sg13g2_a21oi_1 _19482_ (.A1(net4),
    .A2(net8),
    .Y(_03019_),
    .B1(net6544));
 sg13g2_a22oi_1 _19483_ (.Y(_03020_),
    .B1(_11079_),
    .B2(_03019_),
    .A2(net4425),
    .A1(net6545));
 sg13g2_inv_1 _19484_ (.Y(_00180_),
    .A(_03020_));
 sg13g2_nand2_2 _19485_ (.Y(_03021_),
    .A(_09262_),
    .B(_09345_));
 sg13g2_or2_1 _19486_ (.X(_03022_),
    .B(net5912),
    .A(\atari2600.address_bus_r[12] ));
 sg13g2_nor2b_2 _19487_ (.A(_09125_),
    .B_N(_03022_),
    .Y(_03023_));
 sg13g2_o21ai_1 _19488_ (.B1(_03022_),
    .Y(_03024_),
    .A1(net5869),
    .A2(_09124_));
 sg13g2_and2_1 _19489_ (.A(net5514),
    .B(net5536),
    .X(_03025_));
 sg13g2_and3_2 _19490_ (.X(_03026_),
    .A(_09113_),
    .B(_09276_),
    .C(_03025_));
 sg13g2_nand2_2 _19491_ (.Y(_03027_),
    .A(_09349_),
    .B(_03026_));
 sg13g2_nor2_1 _19492_ (.A(_03021_),
    .B(net5258),
    .Y(_03028_));
 sg13g2_nor2_1 _19493_ (.A(net4069),
    .B(net5202),
    .Y(_03029_));
 sg13g2_a21oi_1 _19494_ (.A1(net5774),
    .A2(net5202),
    .Y(_00181_),
    .B1(_03029_));
 sg13g2_nor2_1 _19495_ (.A(net4173),
    .B(net5202),
    .Y(_03030_));
 sg13g2_a21oi_1 _19496_ (.A1(net5794),
    .A2(net5202),
    .Y(_00182_),
    .B1(_03030_));
 sg13g2_nor2_1 _19497_ (.A(net3397),
    .B(net5202),
    .Y(_03031_));
 sg13g2_a21oi_1 _19498_ (.A1(net5724),
    .A2(net5202),
    .Y(_00183_),
    .B1(_03031_));
 sg13g2_nor2_1 _19499_ (.A(net3507),
    .B(net5202),
    .Y(_03032_));
 sg13g2_nor2_1 _19500_ (.A(net5936),
    .B(_09159_),
    .Y(_03033_));
 sg13g2_nor2_1 _19501_ (.A(_00136_),
    .B(_09179_),
    .Y(_03034_));
 sg13g2_a21oi_1 _19502_ (.A1(\atari2600.cpu.PC[11] ),
    .A2(_09181_),
    .Y(_03035_),
    .B1(_03034_));
 sg13g2_a22oi_1 _19503_ (.Y(_03036_),
    .B1(_09177_),
    .B2(_08597_),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[3] ));
 sg13g2_nand3_1 _19504_ (.B(_03035_),
    .C(_03036_),
    .A(net5936),
    .Y(_03037_));
 sg13g2_nor2b_1 _19505_ (.A(_03033_),
    .B_N(_03037_),
    .Y(_03038_));
 sg13g2_o21ai_1 _19506_ (.B1(_03037_),
    .Y(_03039_),
    .A1(net5936),
    .A2(_09159_));
 sg13g2_a21oi_1 _19507_ (.A1(_03028_),
    .A2(net5702),
    .Y(_00184_),
    .B1(_03032_));
 sg13g2_nor2_1 _19508_ (.A(net3424),
    .B(net5201),
    .Y(_03040_));
 sg13g2_nor2_1 _19509_ (.A(_09064_),
    .B(net5936),
    .Y(_03041_));
 sg13g2_o21ai_1 _19510_ (.B1(net6250),
    .Y(_03042_),
    .A1(_08814_),
    .A2(net6031));
 sg13g2_a22oi_1 _19511_ (.Y(_03043_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[12] ),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[4] ));
 sg13g2_nand4_1 _19512_ (.B(_09179_),
    .C(_03042_),
    .A(net5937),
    .Y(_03044_),
    .D(_03043_));
 sg13g2_nor2b_2 _19513_ (.A(_03041_),
    .B_N(_03044_),
    .Y(_03045_));
 sg13g2_o21ai_1 _19514_ (.B1(_03044_),
    .Y(_03046_),
    .A1(_09064_),
    .A2(net5936));
 sg13g2_a21oi_1 _19515_ (.A1(net5201),
    .A2(net5681),
    .Y(_00185_),
    .B1(_03040_));
 sg13g2_nor2_1 _19516_ (.A(net4110),
    .B(net5201),
    .Y(_03047_));
 sg13g2_a22oi_1 _19517_ (.Y(_03048_),
    .B1(net6031),
    .B2(net6249),
    .A2(_08814_),
    .A1(_08596_));
 sg13g2_a22oi_1 _19518_ (.Y(_03049_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[13] ),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[5] ));
 sg13g2_nand3_1 _19519_ (.B(_03048_),
    .C(_03049_),
    .A(_09179_),
    .Y(_03050_));
 sg13g2_nand2_2 _19520_ (.Y(_03051_),
    .A(_09098_),
    .B(_09110_));
 sg13g2_nor2b_1 _19521_ (.A(_03050_),
    .B_N(_03051_),
    .Y(_03052_));
 sg13g2_nand2b_2 _19522_ (.Y(_03053_),
    .B(_03051_),
    .A_N(_03050_));
 sg13g2_a21oi_1 _19523_ (.A1(net5201),
    .A2(net5604),
    .Y(_00186_),
    .B1(_03047_));
 sg13g2_nor2_1 _19524_ (.A(net4352),
    .B(net5201),
    .Y(_03054_));
 sg13g2_nor2_1 _19525_ (.A(net5936),
    .B(_09253_),
    .Y(_03055_));
 sg13g2_nand2b_1 _19526_ (.Y(_03056_),
    .B(_09177_),
    .A_N(_00092_));
 sg13g2_a22oi_1 _19527_ (.Y(_03057_),
    .B1(_09181_),
    .B2(\atari2600.cpu.PC[14] ),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[6] ));
 sg13g2_or2_1 _19528_ (.X(_03058_),
    .B(_09179_),
    .A(_00137_));
 sg13g2_nand4_1 _19529_ (.B(_03056_),
    .C(_03057_),
    .A(net5937),
    .Y(_03059_),
    .D(_03058_));
 sg13g2_nor2b_1 _19530_ (.A(_03055_),
    .B_N(_03059_),
    .Y(_03060_));
 sg13g2_o21ai_1 _19531_ (.B1(_03059_),
    .Y(_03061_),
    .A1(net5936),
    .A2(_09253_));
 sg13g2_a21oi_1 _19532_ (.A1(net5201),
    .A2(net5658),
    .Y(_00187_),
    .B1(_03054_));
 sg13g2_nor2_1 _19533_ (.A(net3708),
    .B(net5201),
    .Y(_03062_));
 sg13g2_nand3_1 _19534_ (.B(_09114_),
    .C(_09115_),
    .A(_09110_),
    .Y(_03063_));
 sg13g2_or2_1 _19535_ (.X(_03064_),
    .B(_09179_),
    .A(_00138_));
 sg13g2_nand2_1 _19536_ (.Y(_03065_),
    .A(\atari2600.cpu.PC[15] ),
    .B(_09181_));
 sg13g2_a22oi_1 _19537_ (.Y(_03066_),
    .B1(_09177_),
    .B2(_08599_),
    .A2(net5989),
    .A1(\atari2600.cpu.PC[7] ));
 sg13g2_nand4_1 _19538_ (.B(_03064_),
    .C(_03065_),
    .A(net5937),
    .Y(_03067_),
    .D(_03066_));
 sg13g2_and2_1 _19539_ (.A(_03063_),
    .B(_03067_),
    .X(_03068_));
 sg13g2_nand2_1 _19540_ (.Y(_03069_),
    .A(_03063_),
    .B(_03067_));
 sg13g2_a21oi_1 _19541_ (.A1(net5201),
    .A2(net5636),
    .Y(_00188_),
    .B1(_03062_));
 sg13g2_nor2_1 _19542_ (.A(net5203),
    .B(net5259),
    .Y(_03070_));
 sg13g2_nor2_1 _19543_ (.A(net3211),
    .B(net5077),
    .Y(_03071_));
 sg13g2_nor2_2 _19544_ (.A(_09350_),
    .B(net5203),
    .Y(_03072_));
 sg13g2_nand2_2 _19545_ (.Y(_03073_),
    .A(_09349_),
    .B(_09413_));
 sg13g2_a21oi_1 _19546_ (.A1(net5762),
    .A2(net5077),
    .Y(_00189_),
    .B1(_03071_));
 sg13g2_nor2_1 _19547_ (.A(net4131),
    .B(net5077),
    .Y(_03074_));
 sg13g2_a21oi_1 _19548_ (.A1(net5782),
    .A2(net5077),
    .Y(_00190_),
    .B1(_03074_));
 sg13g2_nor2_1 _19549_ (.A(net3951),
    .B(net5077),
    .Y(_03075_));
 sg13g2_a21oi_1 _19550_ (.A1(net5712),
    .A2(net5077),
    .Y(_00191_),
    .B1(_03075_));
 sg13g2_nor2_1 _19551_ (.A(net4309),
    .B(net5076),
    .Y(_03076_));
 sg13g2_a21oi_1 _19552_ (.A1(net5690),
    .A2(net5076),
    .Y(_00192_),
    .B1(_03076_));
 sg13g2_nor2_1 _19553_ (.A(net3409),
    .B(net5077),
    .Y(_03077_));
 sg13g2_a21oi_1 _19554_ (.A1(net5668),
    .A2(net5077),
    .Y(_00193_),
    .B1(_03077_));
 sg13g2_nor2_1 _19555_ (.A(net3664),
    .B(net5076),
    .Y(_03078_));
 sg13g2_a21oi_1 _19556_ (.A1(net5591),
    .A2(net5076),
    .Y(_00194_),
    .B1(_03078_));
 sg13g2_nor2_1 _19557_ (.A(net4373),
    .B(net5076),
    .Y(_03079_));
 sg13g2_a21oi_1 _19558_ (.A1(net5650),
    .A2(net5076),
    .Y(_00195_),
    .B1(_03079_));
 sg13g2_nor2_1 _19559_ (.A(net4523),
    .B(net5076),
    .Y(_03080_));
 sg13g2_a21oi_1 _19560_ (.A1(net5629),
    .A2(net5076),
    .Y(_00196_),
    .B1(_03080_));
 sg13g2_nand2b_2 _19561_ (.Y(_03081_),
    .B(_03026_),
    .A_N(_09376_));
 sg13g2_nor2_1 _19562_ (.A(_03021_),
    .B(_03081_),
    .Y(_03082_));
 sg13g2_nor2_1 _19563_ (.A(net3165),
    .B(net5199),
    .Y(_03083_));
 sg13g2_a21oi_1 _19564_ (.A1(net5774),
    .A2(net5199),
    .Y(_00197_),
    .B1(_03083_));
 sg13g2_nor2_1 _19565_ (.A(net3769),
    .B(net5199),
    .Y(_03084_));
 sg13g2_a21oi_1 _19566_ (.A1(net5794),
    .A2(net5199),
    .Y(_00198_),
    .B1(_03084_));
 sg13g2_nor2_1 _19567_ (.A(net3287),
    .B(net5199),
    .Y(_03085_));
 sg13g2_a21oi_1 _19568_ (.A1(net5724),
    .A2(net5199),
    .Y(_00199_),
    .B1(_03085_));
 sg13g2_nor2_1 _19569_ (.A(net3589),
    .B(net5199),
    .Y(_03086_));
 sg13g2_a21oi_1 _19570_ (.A1(net5700),
    .A2(net5199),
    .Y(_00200_),
    .B1(_03086_));
 sg13g2_nor2_1 _19571_ (.A(net3312),
    .B(net5200),
    .Y(_03087_));
 sg13g2_a21oi_1 _19572_ (.A1(net5681),
    .A2(net5200),
    .Y(_00201_),
    .B1(_03087_));
 sg13g2_nor2_1 _19573_ (.A(net3261),
    .B(net5200),
    .Y(_03088_));
 sg13g2_a21oi_1 _19574_ (.A1(net5601),
    .A2(net5200),
    .Y(_00202_),
    .B1(_03088_));
 sg13g2_nor2_1 _19575_ (.A(net3369),
    .B(net5200),
    .Y(_03089_));
 sg13g2_a21oi_1 _19576_ (.A1(net5658),
    .A2(net5200),
    .Y(_00203_),
    .B1(_03089_));
 sg13g2_nor2_1 _19577_ (.A(net3181),
    .B(net5200),
    .Y(_03090_));
 sg13g2_a21oi_1 _19578_ (.A1(net5637),
    .A2(net5200),
    .Y(_00204_),
    .B1(_03090_));
 sg13g2_nand3_1 _19579_ (.B(net5555),
    .C(net5545),
    .A(_09105_),
    .Y(_03091_));
 sg13g2_nor2b_1 _19580_ (.A(net5567),
    .B_N(_03026_),
    .Y(_03092_));
 sg13g2_nand2_2 _19581_ (.Y(_03093_),
    .A(_09312_),
    .B(_03092_));
 sg13g2_nor2_1 _19582_ (.A(_03091_),
    .B(net5239),
    .Y(_03094_));
 sg13g2_nor2_1 _19583_ (.A(net4133),
    .B(net5197),
    .Y(_03095_));
 sg13g2_a21oi_1 _19584_ (.A1(net5772),
    .A2(net5197),
    .Y(_00205_),
    .B1(_03095_));
 sg13g2_nor2_1 _19585_ (.A(net3906),
    .B(net5198),
    .Y(_03096_));
 sg13g2_a21oi_1 _19586_ (.A1(net5792),
    .A2(net5198),
    .Y(_00206_),
    .B1(_03096_));
 sg13g2_nor2_1 _19587_ (.A(net3130),
    .B(net5198),
    .Y(_03097_));
 sg13g2_a21oi_1 _19588_ (.A1(net5722),
    .A2(net5198),
    .Y(_00207_),
    .B1(_03097_));
 sg13g2_nor2_1 _19589_ (.A(net3884),
    .B(net5198),
    .Y(_03098_));
 sg13g2_a21oi_1 _19590_ (.A1(net5699),
    .A2(net5198),
    .Y(_00208_),
    .B1(_03098_));
 sg13g2_nor2_1 _19591_ (.A(net3282),
    .B(net5198),
    .Y(_03099_));
 sg13g2_a21oi_1 _19592_ (.A1(net5679),
    .A2(net5197),
    .Y(_00209_),
    .B1(_03099_));
 sg13g2_nor2_1 _19593_ (.A(net3325),
    .B(net5197),
    .Y(_03100_));
 sg13g2_a21oi_1 _19594_ (.A1(net5596),
    .A2(net5197),
    .Y(_00210_),
    .B1(_03100_));
 sg13g2_nor2_1 _19595_ (.A(net3010),
    .B(_03094_),
    .Y(_03101_));
 sg13g2_a21oi_1 _19596_ (.A1(net5661),
    .A2(net5197),
    .Y(_00211_),
    .B1(_03101_));
 sg13g2_nor2_1 _19597_ (.A(net3108),
    .B(net5197),
    .Y(_03102_));
 sg13g2_a21oi_1 _19598_ (.A1(net5632),
    .A2(net5197),
    .Y(_00212_),
    .B1(_03102_));
 sg13g2_nand2_2 _19599_ (.Y(_03103_),
    .A(_09353_),
    .B(_03026_));
 sg13g2_nor2_1 _19600_ (.A(_03021_),
    .B(_03103_),
    .Y(_03104_));
 sg13g2_nor2_1 _19601_ (.A(net3128),
    .B(net5195),
    .Y(_03105_));
 sg13g2_a21oi_1 _19602_ (.A1(net5774),
    .A2(net5195),
    .Y(_00213_),
    .B1(_03105_));
 sg13g2_nor2_1 _19603_ (.A(net3598),
    .B(net5195),
    .Y(_03106_));
 sg13g2_a21oi_1 _19604_ (.A1(net5794),
    .A2(net5195),
    .Y(_00214_),
    .B1(_03106_));
 sg13g2_nor2_1 _19605_ (.A(net3189),
    .B(net5195),
    .Y(_03107_));
 sg13g2_a21oi_1 _19606_ (.A1(net5724),
    .A2(net5195),
    .Y(_00215_),
    .B1(_03107_));
 sg13g2_nor2_1 _19607_ (.A(net3910),
    .B(net5195),
    .Y(_03108_));
 sg13g2_a21oi_1 _19608_ (.A1(net5700),
    .A2(net5195),
    .Y(_00216_),
    .B1(_03108_));
 sg13g2_nor2_1 _19609_ (.A(net3192),
    .B(net5196),
    .Y(_03109_));
 sg13g2_a21oi_1 _19610_ (.A1(net5681),
    .A2(net5196),
    .Y(_00217_),
    .B1(_03109_));
 sg13g2_nor2_1 _19611_ (.A(net3081),
    .B(net5196),
    .Y(_03110_));
 sg13g2_a21oi_1 _19612_ (.A1(net5601),
    .A2(net5196),
    .Y(_00218_),
    .B1(_03110_));
 sg13g2_nor2_1 _19613_ (.A(net3326),
    .B(net5196),
    .Y(_03111_));
 sg13g2_a21oi_1 _19614_ (.A1(net5659),
    .A2(net5196),
    .Y(_00219_),
    .B1(_03111_));
 sg13g2_nor2_1 _19615_ (.A(net3908),
    .B(net5196),
    .Y(_03112_));
 sg13g2_a21oi_1 _19616_ (.A1(net5636),
    .A2(net5196),
    .Y(_00220_),
    .B1(_03112_));
 sg13g2_nor2_1 _19617_ (.A(net5256),
    .B(_03091_),
    .Y(_03113_));
 sg13g2_nor2_1 _19618_ (.A(net3868),
    .B(net5194),
    .Y(_03114_));
 sg13g2_a21oi_1 _19619_ (.A1(net5772),
    .A2(net5194),
    .Y(_00221_),
    .B1(_03114_));
 sg13g2_nor2_1 _19620_ (.A(net3250),
    .B(net5193),
    .Y(_03115_));
 sg13g2_a21oi_1 _19621_ (.A1(net5792),
    .A2(net5193),
    .Y(_00222_),
    .B1(_03115_));
 sg13g2_nor2_1 _19622_ (.A(net4251),
    .B(net5193),
    .Y(_03116_));
 sg13g2_a21oi_1 _19623_ (.A1(net5722),
    .A2(net5193),
    .Y(_00223_),
    .B1(_03116_));
 sg13g2_nor2_1 _19624_ (.A(net4315),
    .B(net5193),
    .Y(_03117_));
 sg13g2_a21oi_1 _19625_ (.A1(net5699),
    .A2(net5193),
    .Y(_00224_),
    .B1(_03117_));
 sg13g2_nor2_1 _19626_ (.A(net4289),
    .B(net5193),
    .Y(_03118_));
 sg13g2_a21oi_1 _19627_ (.A1(net5679),
    .A2(net5193),
    .Y(_00225_),
    .B1(_03118_));
 sg13g2_nor2_1 _19628_ (.A(net4012),
    .B(net5194),
    .Y(_03119_));
 sg13g2_a21oi_1 _19629_ (.A1(net5598),
    .A2(net5194),
    .Y(_00226_),
    .B1(_03119_));
 sg13g2_nor2_1 _19630_ (.A(net3645),
    .B(net5194),
    .Y(_03120_));
 sg13g2_a21oi_1 _19631_ (.A1(net5661),
    .A2(net5194),
    .Y(_00227_),
    .B1(_03120_));
 sg13g2_nor2_1 _19632_ (.A(net4219),
    .B(net5194),
    .Y(_03121_));
 sg13g2_a21oi_1 _19633_ (.A1(net5632),
    .A2(net5194),
    .Y(_00228_),
    .B1(_03121_));
 sg13g2_nor2_2 _19634_ (.A(net5555),
    .B(_09260_),
    .Y(_03122_));
 sg13g2_nand2_2 _19635_ (.Y(_03123_),
    .A(net5551),
    .B(net5546));
 sg13g2_nand2_2 _19636_ (.Y(_03124_),
    .A(_09105_),
    .B(_03122_));
 sg13g2_and3_2 _19637_ (.X(_03125_),
    .A(net5561),
    .B(net5357),
    .C(_03026_));
 sg13g2_nand3_1 _19638_ (.B(_03122_),
    .C(_03125_),
    .A(_09105_),
    .Y(_03126_));
 sg13g2_mux2_1 _19639_ (.A0(net5742),
    .A1(net7171),
    .S(_03126_),
    .X(_00229_));
 sg13g2_mux2_1 _19640_ (.A0(net5747),
    .A1(net4601),
    .S(_03126_),
    .X(_00230_));
 sg13g2_mux2_1 _19641_ (.A0(net5618),
    .A1(net6591),
    .S(_03126_),
    .X(_00231_));
 sg13g2_mux2_1 _19642_ (.A0(net5612),
    .A1(net6670),
    .S(_03126_),
    .X(_00232_));
 sg13g2_mux2_1 _19643_ (.A0(net5609),
    .A1(net6754),
    .S(_03126_),
    .X(_00233_));
 sg13g2_mux2_1 _19644_ (.A0(net5584),
    .A1(net4762),
    .S(_03126_),
    .X(_00234_));
 sg13g2_mux2_1 _19645_ (.A0(net5579),
    .A1(net6955),
    .S(_03126_),
    .X(_00235_));
 sg13g2_mux2_1 _19646_ (.A0(net5643),
    .A1(net7048),
    .S(_03126_),
    .X(_00236_));
 sg13g2_and2_1 _19647_ (.A(_10001_),
    .B(net6072),
    .X(_03127_));
 sg13g2_nand2_2 _19648_ (.Y(_03128_),
    .A(_10001_),
    .B(net6072));
 sg13g2_nor2_2 _19649_ (.A(_08626_),
    .B(net6503),
    .Y(_03129_));
 sg13g2_nand2_2 _19650_ (.Y(_03130_),
    .A(net6501),
    .B(net6124));
 sg13g2_nor2_2 _19651_ (.A(_10124_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_nand2_2 _19652_ (.Y(_03132_),
    .A(_10123_),
    .B(_03129_));
 sg13g2_nand2_2 _19653_ (.Y(_03133_),
    .A(net6028),
    .B(_03131_));
 sg13g2_mux2_1 _19654_ (.A0(net6456),
    .A1(net7055),
    .S(_03133_),
    .X(_00237_));
 sg13g2_mux2_1 _19655_ (.A0(net6426),
    .A1(net4727),
    .S(_03133_),
    .X(_00238_));
 sg13g2_mux2_1 _19656_ (.A0(net6398),
    .A1(net4843),
    .S(_03133_),
    .X(_00239_));
 sg13g2_mux2_1 _19657_ (.A0(net6368),
    .A1(net7071),
    .S(_03133_),
    .X(_00240_));
 sg13g2_mux2_1 _19658_ (.A0(net6336),
    .A1(net6991),
    .S(_03133_),
    .X(_00241_));
 sg13g2_mux2_1 _19659_ (.A0(net6310),
    .A1(net6793),
    .S(_03133_),
    .X(_00242_));
 sg13g2_mux2_1 _19660_ (.A0(net6279),
    .A1(net4520),
    .S(_03133_),
    .X(_00243_));
 sg13g2_nand2_2 _19661_ (.Y(_03134_),
    .A(net5550),
    .B(_09321_));
 sg13g2_nor2_1 _19662_ (.A(net5257),
    .B(_03134_),
    .Y(_03135_));
 sg13g2_nor2_1 _19663_ (.A(net3952),
    .B(net5075),
    .Y(_03136_));
 sg13g2_a21oi_1 _19664_ (.A1(net5769),
    .A2(net5075),
    .Y(_00244_),
    .B1(_03136_));
 sg13g2_nor2_1 _19665_ (.A(net3949),
    .B(net5073),
    .Y(_03137_));
 sg13g2_a21oi_1 _19666_ (.A1(net5789),
    .A2(net5073),
    .Y(_00245_),
    .B1(_03137_));
 sg13g2_nor2_1 _19667_ (.A(net4332),
    .B(net5075),
    .Y(_03138_));
 sg13g2_a21oi_1 _19668_ (.A1(net5719),
    .A2(net5075),
    .Y(_00246_),
    .B1(_03138_));
 sg13g2_nor2_1 _19669_ (.A(net3435),
    .B(net5074),
    .Y(_03139_));
 sg13g2_a21oi_1 _19670_ (.A1(net5695),
    .A2(net5074),
    .Y(_00247_),
    .B1(_03139_));
 sg13g2_nor2_1 _19671_ (.A(net3641),
    .B(net5073),
    .Y(_03140_));
 sg13g2_a21oi_1 _19672_ (.A1(net5672),
    .A2(net5073),
    .Y(_00248_),
    .B1(_03140_));
 sg13g2_nor2_1 _19673_ (.A(net3444),
    .B(net5074),
    .Y(_03141_));
 sg13g2_a21oi_1 _19674_ (.A1(net5593),
    .A2(net5074),
    .Y(_00249_),
    .B1(_03141_));
 sg13g2_nor2_1 _19675_ (.A(net3344),
    .B(net5073),
    .Y(_03142_));
 sg13g2_a21oi_1 _19676_ (.A1(net5656),
    .A2(net5073),
    .Y(_00250_),
    .B1(_03142_));
 sg13g2_nor2_1 _19677_ (.A(net4185),
    .B(net5073),
    .Y(_03143_));
 sg13g2_a21oi_1 _19678_ (.A1(net5630),
    .A2(net5073),
    .Y(_00251_),
    .B1(_03143_));
 sg13g2_nor2_1 _19679_ (.A(_09441_),
    .B(_03027_),
    .Y(_03144_));
 sg13g2_nor2_1 _19680_ (.A(net3797),
    .B(_03144_),
    .Y(_03145_));
 sg13g2_a21oi_1 _19681_ (.A1(net5768),
    .A2(net5072),
    .Y(_00252_),
    .B1(_03145_));
 sg13g2_nor2_1 _19682_ (.A(net4075),
    .B(net5072),
    .Y(_03146_));
 sg13g2_a21oi_1 _19683_ (.A1(net5788),
    .A2(net5072),
    .Y(_00253_),
    .B1(_03146_));
 sg13g2_nor2_1 _19684_ (.A(net3553),
    .B(net5071),
    .Y(_03147_));
 sg13g2_a21oi_1 _19685_ (.A1(net5718),
    .A2(net5071),
    .Y(_00254_),
    .B1(_03147_));
 sg13g2_nor2_1 _19686_ (.A(net3573),
    .B(net5071),
    .Y(_03148_));
 sg13g2_a21oi_1 _19687_ (.A1(net5695),
    .A2(net5071),
    .Y(_00255_),
    .B1(_03148_));
 sg13g2_nor2_1 _19688_ (.A(net4236),
    .B(net5072),
    .Y(_03149_));
 sg13g2_a21oi_1 _19689_ (.A1(net5674),
    .A2(net5072),
    .Y(_00256_),
    .B1(_03149_));
 sg13g2_nor2_1 _19690_ (.A(net4192),
    .B(net5072),
    .Y(_03150_));
 sg13g2_a21oi_1 _19691_ (.A1(net5593),
    .A2(net5072),
    .Y(_00257_),
    .B1(_03150_));
 sg13g2_nor2_1 _19692_ (.A(net4330),
    .B(net5071),
    .Y(_03151_));
 sg13g2_a21oi_1 _19693_ (.A1(net5657),
    .A2(net5071),
    .Y(_00258_),
    .B1(_03151_));
 sg13g2_nor2_1 _19694_ (.A(net4071),
    .B(net5071),
    .Y(_03152_));
 sg13g2_a21oi_1 _19695_ (.A1(net5635),
    .A2(net5071),
    .Y(_00259_),
    .B1(_03152_));
 sg13g2_nand2_1 _19696_ (.Y(_03153_),
    .A(net3336),
    .B(net6544));
 sg13g2_xnor2_1 _19697_ (.Y(_03154_),
    .A(_08615_),
    .B(_09283_));
 sg13g2_xnor2_1 _19698_ (.Y(_03155_),
    .A(\rom_next_addr_in_queue[6] ),
    .B(net5544));
 sg13g2_xnor2_1 _19699_ (.Y(_03156_),
    .A(\rom_next_addr_in_queue[3] ),
    .B(net5556));
 sg13g2_nor2_1 _19700_ (.A(\rom_next_addr_in_queue[5] ),
    .B(net5570),
    .Y(_03157_));
 sg13g2_xnor2_1 _19701_ (.Y(_03158_),
    .A(\rom_next_addr_in_queue[2] ),
    .B(net5563));
 sg13g2_xnor2_1 _19702_ (.Y(_03159_),
    .A(\rom_next_addr_in_queue[11] ),
    .B(net5541));
 sg13g2_xnor2_1 _19703_ (.Y(_03160_),
    .A(\rom_last_read_addr[11] ),
    .B(net5541));
 sg13g2_nor2_1 _19704_ (.A(\rom_last_read_addr[8] ),
    .B(_09272_),
    .Y(_03161_));
 sg13g2_xnor2_1 _19705_ (.Y(_03162_),
    .A(\rom_last_read_addr[4] ),
    .B(net5280));
 sg13g2_xnor2_1 _19706_ (.Y(_03163_),
    .A(\rom_last_read_addr[3] ),
    .B(net5548));
 sg13g2_xor2_1 _19707_ (.B(_09135_),
    .A(\rom_last_read_addr[1] ),
    .X(_03164_));
 sg13g2_xor2_1 _19708_ (.B(_09283_),
    .A(\rom_last_read_addr[10] ),
    .X(_03165_));
 sg13g2_xnor2_1 _19709_ (.Y(_03166_),
    .A(_08602_),
    .B(net5514));
 sg13g2_xnor2_1 _19710_ (.Y(_03167_),
    .A(\rom_last_read_addr[2] ),
    .B(net5560));
 sg13g2_xnor2_1 _19711_ (.Y(_03168_),
    .A(\rom_last_read_addr[5] ),
    .B(net5570));
 sg13g2_nor4_1 _19712_ (.A(_03163_),
    .B(_03166_),
    .C(_03167_),
    .D(_03168_),
    .Y(_03169_));
 sg13g2_a22oi_1 _19713_ (.Y(_03170_),
    .B1(_09277_),
    .B2(_08604_),
    .A2(_09272_),
    .A1(\rom_last_read_addr[8] ));
 sg13g2_a22oi_1 _19714_ (.Y(_03171_),
    .B1(_09278_),
    .B2(\rom_last_read_addr[9] ),
    .A2(net5529),
    .A1(_08600_));
 sg13g2_a221oi_1 _19715_ (.B2(\rom_last_read_addr[6] ),
    .C1(_03161_),
    .B1(net5543),
    .A1(\rom_last_read_addr[0] ),
    .Y(_03172_),
    .A2(net5532));
 sg13g2_and4_1 _19716_ (.A(_03160_),
    .B(_03170_),
    .C(_03171_),
    .D(_03172_),
    .X(_03173_));
 sg13g2_o21ai_1 _19717_ (.B1(_03165_),
    .Y(_03174_),
    .A1(\rom_last_read_addr[6] ),
    .A2(net5543));
 sg13g2_nor3_1 _19718_ (.A(_03162_),
    .B(_03164_),
    .C(_03174_),
    .Y(_03175_));
 sg13g2_nand3_1 _19719_ (.B(_03173_),
    .C(_03175_),
    .A(_03169_),
    .Y(_03176_));
 sg13g2_xnor2_1 _19720_ (.Y(_03177_),
    .A(\rom_next_addr_in_queue[1] ),
    .B(net5564));
 sg13g2_xnor2_1 _19721_ (.Y(_03178_),
    .A(_08614_),
    .B(_09272_));
 sg13g2_nand3_1 _19722_ (.B(_03177_),
    .C(_03178_),
    .A(_03158_),
    .Y(_03179_));
 sg13g2_xnor2_1 _19723_ (.Y(_03180_),
    .A(\rom_next_addr_in_queue[4] ),
    .B(net5280));
 sg13g2_xnor2_1 _19724_ (.Y(_03181_),
    .A(_08613_),
    .B(net5514));
 sg13g2_a21oi_1 _19725_ (.A1(_00093_),
    .A2(net5529),
    .Y(_03182_),
    .B1(_03157_));
 sg13g2_nand3_1 _19726_ (.B(_03159_),
    .C(_03182_),
    .A(_03155_),
    .Y(_03183_));
 sg13g2_nor4_1 _19727_ (.A(_03179_),
    .B(_03180_),
    .C(_03181_),
    .D(_03183_),
    .Y(_03184_));
 sg13g2_xor2_1 _19728_ (.B(_09277_),
    .A(\rom_next_addr_in_queue[9] ),
    .X(_03185_));
 sg13g2_a221oi_1 _19729_ (.B2(_08608_),
    .C1(_03185_),
    .B1(net5532),
    .A1(\rom_next_addr_in_queue[5] ),
    .Y(_03186_),
    .A2(net5570));
 sg13g2_nand4_1 _19730_ (.B(_03156_),
    .C(_03184_),
    .A(_03154_),
    .Y(_03187_),
    .D(_03186_));
 sg13g2_nand4_1 _19731_ (.B(_03023_),
    .C(_03176_),
    .A(net5857),
    .Y(_03188_),
    .D(_03187_));
 sg13g2_a21oi_1 _19732_ (.A1(_03153_),
    .A2(_03188_),
    .Y(_00260_),
    .B1(\flash_rom.spi_select ));
 sg13g2_or4_1 _19733_ (.A(_08625_),
    .B(net5853),
    .C(net5536),
    .D(_03187_),
    .X(_03189_));
 sg13g2_o21ai_1 _19734_ (.B1(_03189_),
    .Y(_03190_),
    .A1(net7362),
    .A2(rom_data_pending));
 sg13g2_inv_1 _19735_ (.Y(_00261_),
    .A(_03190_));
 sg13g2_and2_1 _19736_ (.A(net7561),
    .B(net7468),
    .X(_03191_));
 sg13g2_nand3_1 _19737_ (.B(net6209),
    .C(_03191_),
    .A(net6154),
    .Y(_03192_));
 sg13g2_nor2b_2 _19738_ (.A(net6133),
    .B_N(net6134),
    .Y(_03193_));
 sg13g2_nand2b_1 _19739_ (.Y(_03194_),
    .B(net6134),
    .A_N(net6133));
 sg13g2_nand2_2 _19740_ (.Y(_03195_),
    .A(net6115),
    .B(net6113));
 sg13g2_nand3_1 _19741_ (.B(net6126),
    .C(net6061),
    .A(\hvsync_gen.hpos[9] ),
    .Y(_03196_));
 sg13g2_nor3_2 _19742_ (.A(_03192_),
    .B(net6025),
    .C(_03196_),
    .Y(_03197_));
 sg13g2_nor2_2 _19743_ (.A(net6540),
    .B(_03197_),
    .Y(_03198_));
 sg13g2_nand2b_2 _19744_ (.Y(_03199_),
    .B(net6575),
    .A_N(_03197_));
 sg13g2_and2_1 _19745_ (.A(net2930),
    .B(_03198_),
    .X(_00262_));
 sg13g2_nor2_1 _19746_ (.A(\hvsync_gen.hpos[0] ),
    .B(net7468),
    .Y(_03200_));
 sg13g2_nor3_1 _19747_ (.A(_03191_),
    .B(_03199_),
    .C(net7469),
    .Y(_00263_));
 sg13g2_nor2_1 _19748_ (.A(_08625_),
    .B(spi_data_ready_last),
    .Y(_03201_));
 sg13g2_nand2b_1 _19749_ (.Y(_03202_),
    .B(net2932),
    .A_N(spi_data_ready_last));
 sg13g2_nor2b_1 _19750_ (.A(spi_restart),
    .B_N(_03188_),
    .Y(_03203_));
 sg13g2_nor2_1 _19751_ (.A(_09038_),
    .B(_03203_),
    .Y(_03204_));
 sg13g2_inv_1 _19752_ (.Y(_03205_),
    .A(net4989));
 sg13g2_nand3_1 _19753_ (.B(net6055),
    .C(net4987),
    .A(net5529),
    .Y(_03206_));
 sg13g2_nor3_1 _19754_ (.A(net6523),
    .B(net6022),
    .C(net4986),
    .Y(_03207_));
 sg13g2_nand3_1 _19755_ (.B(net6055),
    .C(net4982),
    .A(net6544),
    .Y(_03208_));
 sg13g2_nand2_1 _19756_ (.Y(_03209_),
    .A(net7165),
    .B(net6023));
 sg13g2_nor2b_1 _19757_ (.A(net4979),
    .B_N(_03209_),
    .Y(_03210_));
 sg13g2_a22oi_1 _19758_ (.Y(_00264_),
    .B1(_03210_),
    .B2(_03206_),
    .A2(net4979),
    .A1(_08600_));
 sg13g2_nand2_1 _19759_ (.Y(_03211_),
    .A(net7075),
    .B(net4979));
 sg13g2_nand2_1 _19760_ (.Y(_03212_),
    .A(\rom_next_addr_in_queue[1] ),
    .B(net6023));
 sg13g2_nand3_1 _19761_ (.B(net6055),
    .C(net4987),
    .A(net5564),
    .Y(_03213_));
 sg13g2_nand3_1 _19762_ (.B(_03212_),
    .C(_03213_),
    .A(_03211_),
    .Y(_00265_));
 sg13g2_a21oi_1 _19763_ (.A1(net5563),
    .A2(net4987),
    .Y(_03214_),
    .B1(net6023));
 sg13g2_a21oi_1 _19764_ (.A1(_08609_),
    .A2(net6023),
    .Y(_03215_),
    .B1(_03214_));
 sg13g2_a21o_1 _19765_ (.A2(net4979),
    .A1(net4509),
    .B1(_03215_),
    .X(_00266_));
 sg13g2_nor3_1 _19766_ (.A(net5548),
    .B(net6023),
    .C(net4983),
    .Y(_03216_));
 sg13g2_a21o_1 _19767_ (.A2(net6023),
    .A1(\rom_next_addr_in_queue[3] ),
    .B1(_03216_),
    .X(_03217_));
 sg13g2_a21o_1 _19768_ (.A2(net4979),
    .A1(net4670),
    .B1(_03217_),
    .X(_00267_));
 sg13g2_nand2_1 _19769_ (.Y(_03218_),
    .A(net5275),
    .B(net4987));
 sg13g2_nor2_1 _19770_ (.A(net6022),
    .B(_03218_),
    .Y(_03219_));
 sg13g2_a21oi_1 _19771_ (.A1(\rom_next_addr_in_queue[4] ),
    .A2(net6022),
    .Y(_03220_),
    .B1(_03219_));
 sg13g2_nor2_1 _19772_ (.A(net6626),
    .B(net4976),
    .Y(_03221_));
 sg13g2_a21oi_1 _19773_ (.A1(net4976),
    .A2(_03220_),
    .Y(_00268_),
    .B1(_03221_));
 sg13g2_nor3_1 _19774_ (.A(net5570),
    .B(net6024),
    .C(net4982),
    .Y(_03222_));
 sg13g2_a21oi_1 _19775_ (.A1(\rom_next_addr_in_queue[5] ),
    .A2(net6022),
    .Y(_03223_),
    .B1(_03222_));
 sg13g2_nor2_1 _19776_ (.A(net4336),
    .B(net4976),
    .Y(_03224_));
 sg13g2_a21oi_1 _19777_ (.A1(net4976),
    .A2(_03223_),
    .Y(_00269_),
    .B1(_03224_));
 sg13g2_nand2_1 _19778_ (.Y(_03225_),
    .A(net5544),
    .B(net4986));
 sg13g2_nand3_1 _19779_ (.B(net6055),
    .C(net4986),
    .A(net5544),
    .Y(_03226_));
 sg13g2_a21oi_1 _19780_ (.A1(\rom_next_addr_in_queue[6] ),
    .A2(net6022),
    .Y(_03227_),
    .B1(net4978));
 sg13g2_a22oi_1 _19781_ (.Y(_00270_),
    .B1(_03226_),
    .B2(_03227_),
    .A2(net4977),
    .A1(_08601_));
 sg13g2_nand2_1 _19782_ (.Y(_03228_),
    .A(net5514),
    .B(net4986));
 sg13g2_nand3_1 _19783_ (.B(net6055),
    .C(net4987),
    .A(net5514),
    .Y(_03229_));
 sg13g2_a21oi_1 _19784_ (.A1(\rom_next_addr_in_queue[7] ),
    .A2(net6022),
    .Y(_03230_),
    .B1(net4980));
 sg13g2_a22oi_1 _19785_ (.Y(_00271_),
    .B1(_03229_),
    .B2(_03230_),
    .A2(net4980),
    .A1(_08602_));
 sg13g2_nor3_1 _19786_ (.A(_09272_),
    .B(net6021),
    .C(net4982),
    .Y(_03231_));
 sg13g2_a21oi_1 _19787_ (.A1(\rom_next_addr_in_queue[8] ),
    .A2(net6021),
    .Y(_03232_),
    .B1(_03231_));
 sg13g2_nor2_1 _19788_ (.A(net4919),
    .B(net4975),
    .Y(_03233_));
 sg13g2_a21oi_1 _19789_ (.A1(net4975),
    .A2(_03232_),
    .Y(_00272_),
    .B1(_03233_));
 sg13g2_nand2_1 _19790_ (.Y(_03234_),
    .A(_09277_),
    .B(net4988));
 sg13g2_nand3_1 _19791_ (.B(net6055),
    .C(net4986),
    .A(_09277_),
    .Y(_03235_));
 sg13g2_a21oi_1 _19792_ (.A1(\rom_next_addr_in_queue[9] ),
    .A2(net6021),
    .Y(_03236_),
    .B1(net4977));
 sg13g2_a22oi_1 _19793_ (.Y(_00273_),
    .B1(_03235_),
    .B2(_03236_),
    .A2(net4977),
    .A1(_08604_));
 sg13g2_nor3_1 _19794_ (.A(_09283_),
    .B(net6021),
    .C(net4982),
    .Y(_03237_));
 sg13g2_a21oi_1 _19795_ (.A1(\rom_next_addr_in_queue[10] ),
    .A2(net6021),
    .Y(_03238_),
    .B1(_03237_));
 sg13g2_nor2_1 _19796_ (.A(net4370),
    .B(net4975),
    .Y(_03239_));
 sg13g2_a21oi_1 _19797_ (.A1(net4975),
    .A2(_03238_),
    .Y(_00274_),
    .B1(_03239_));
 sg13g2_nand2_1 _19798_ (.Y(_03240_),
    .A(net5541),
    .B(net4984));
 sg13g2_nand3_1 _19799_ (.B(net6055),
    .C(net4984),
    .A(net5541),
    .Y(_03241_));
 sg13g2_a21oi_1 _19800_ (.A1(\rom_next_addr_in_queue[11] ),
    .A2(net6021),
    .Y(_03242_),
    .B1(net4977));
 sg13g2_a22oi_1 _19801_ (.Y(_00275_),
    .B1(_03241_),
    .B2(_03242_),
    .A2(net4977),
    .A1(_08606_));
 sg13g2_nand2_2 _19802_ (.Y(_03243_),
    .A(_09413_),
    .B(net5252));
 sg13g2_mux2_1 _19803_ (.A0(net5740),
    .A1(net4798),
    .S(_03243_),
    .X(_00276_));
 sg13g2_mux2_1 _19804_ (.A0(net5745),
    .A1(net4616),
    .S(_03243_),
    .X(_00277_));
 sg13g2_mux2_1 _19805_ (.A0(net5621),
    .A1(net6928),
    .S(_03243_),
    .X(_00278_));
 sg13g2_mux2_1 _19806_ (.A0(net5615),
    .A1(net4557),
    .S(_03243_),
    .X(_00279_));
 sg13g2_mux2_1 _19807_ (.A0(net5607),
    .A1(net6618),
    .S(_03243_),
    .X(_00280_));
 sg13g2_mux2_1 _19808_ (.A0(net5582),
    .A1(net4954),
    .S(_03243_),
    .X(_00281_));
 sg13g2_mux2_1 _19809_ (.A0(net5575),
    .A1(net6939),
    .S(_03243_),
    .X(_00282_));
 sg13g2_mux2_1 _19810_ (.A0(net5641),
    .A1(net6643),
    .S(_03243_),
    .X(_00283_));
 sg13g2_a21oi_1 _19811_ (.A1(_00093_),
    .A2(net6023),
    .Y(_03244_),
    .B1(net4979));
 sg13g2_a22oi_1 _19812_ (.Y(_00284_),
    .B1(_03244_),
    .B2(_03206_),
    .A2(net4979),
    .A1(_08607_));
 sg13g2_nand2_1 _19813_ (.Y(_03245_),
    .A(net7223),
    .B(net4979));
 sg13g2_and3_1 _19814_ (.X(_03246_),
    .A(_03209_),
    .B(_03212_),
    .C(_03213_));
 sg13g2_nand3_1 _19815_ (.B(\rom_next_addr_in_queue[1] ),
    .C(net6023),
    .A(net7165),
    .Y(_03247_));
 sg13g2_nand2_1 _19816_ (.Y(_03248_),
    .A(net4976),
    .B(_03247_));
 sg13g2_o21ai_1 _19817_ (.B1(_03245_),
    .Y(_00285_),
    .A1(_03246_),
    .A2(_03248_));
 sg13g2_nor2_1 _19818_ (.A(_03215_),
    .B(_03248_),
    .Y(_03249_));
 sg13g2_nor2_1 _19819_ (.A(net7369),
    .B(net4976),
    .Y(_03250_));
 sg13g2_nor2_1 _19820_ (.A(_08609_),
    .B(_03247_),
    .Y(_03251_));
 sg13g2_nor3_1 _19821_ (.A(_03249_),
    .B(_03250_),
    .C(_03251_),
    .Y(_00286_));
 sg13g2_and4_1 _19822_ (.A(\rom_next_addr_in_queue[0] ),
    .B(\rom_next_addr_in_queue[1] ),
    .C(\rom_next_addr_in_queue[2] ),
    .D(\rom_next_addr_in_queue[3] ),
    .X(_03252_));
 sg13g2_nand2b_1 _19823_ (.Y(_03253_),
    .B(_03252_),
    .A_N(_03216_));
 sg13g2_o21ai_1 _19824_ (.B1(_03253_),
    .Y(_03254_),
    .A1(_03217_),
    .A2(_03251_));
 sg13g2_o21ai_1 _19825_ (.B1(_03254_),
    .Y(_00287_),
    .A1(_08610_),
    .A2(net4975));
 sg13g2_and2_1 _19826_ (.A(\rom_next_addr_in_queue[4] ),
    .B(_03252_),
    .X(_03255_));
 sg13g2_o21ai_1 _19827_ (.B1(net6022),
    .Y(_03256_),
    .A1(\rom_next_addr_in_queue[4] ),
    .A2(_03252_));
 sg13g2_nor2_1 _19828_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 sg13g2_nor3_1 _19829_ (.A(net4980),
    .B(_03219_),
    .C(_03257_),
    .Y(_03258_));
 sg13g2_a21oi_1 _19830_ (.A1(_08611_),
    .A2(net4980),
    .Y(_00288_),
    .B1(_03258_));
 sg13g2_and2_1 _19831_ (.A(\rom_next_addr_in_queue[5] ),
    .B(_03255_),
    .X(_03259_));
 sg13g2_o21ai_1 _19832_ (.B1(net6022),
    .Y(_03260_),
    .A1(\rom_next_addr_in_queue[5] ),
    .A2(_03255_));
 sg13g2_nor2_1 _19833_ (.A(_03259_),
    .B(_03260_),
    .Y(_03261_));
 sg13g2_nor3_1 _19834_ (.A(net4980),
    .B(_03222_),
    .C(_03261_),
    .Y(_03262_));
 sg13g2_a21oi_1 _19835_ (.A1(_08612_),
    .A2(net4980),
    .Y(_00289_),
    .B1(_03262_));
 sg13g2_a21oi_1 _19836_ (.A1(\rom_next_addr_in_queue[6] ),
    .A2(_03259_),
    .Y(_03263_),
    .B1(net6055));
 sg13g2_o21ai_1 _19837_ (.B1(_03263_),
    .Y(_03264_),
    .A1(\rom_next_addr_in_queue[6] ),
    .A2(_03259_));
 sg13g2_nand3_1 _19838_ (.B(_03226_),
    .C(_03264_),
    .A(net4975),
    .Y(_03265_));
 sg13g2_o21ai_1 _19839_ (.B1(_03265_),
    .Y(_03266_),
    .A1(net7478),
    .A2(net4975));
 sg13g2_inv_1 _19840_ (.Y(_00290_),
    .A(_03266_));
 sg13g2_a21oi_1 _19841_ (.A1(\rom_next_addr_in_queue[6] ),
    .A2(_03259_),
    .Y(_03267_),
    .B1(net7422));
 sg13g2_and3_1 _19842_ (.X(_03268_),
    .A(\rom_next_addr_in_queue[6] ),
    .B(\rom_next_addr_in_queue[7] ),
    .C(_03259_));
 sg13g2_nor3_1 _19843_ (.A(_03202_),
    .B(_03267_),
    .C(_03268_),
    .Y(_03269_));
 sg13g2_nor2_1 _19844_ (.A(net4980),
    .B(_03269_),
    .Y(_03270_));
 sg13g2_a22oi_1 _19845_ (.Y(_00291_),
    .B1(_03229_),
    .B2(_03270_),
    .A2(net4980),
    .A1(_08613_));
 sg13g2_and2_1 _19846_ (.A(\rom_next_addr_in_queue[8] ),
    .B(_03268_),
    .X(_03271_));
 sg13g2_o21ai_1 _19847_ (.B1(net6024),
    .Y(_03272_),
    .A1(net7316),
    .A2(_03268_));
 sg13g2_nor2_1 _19848_ (.A(_03271_),
    .B(_03272_),
    .Y(_03273_));
 sg13g2_nor3_1 _19849_ (.A(net4978),
    .B(_03231_),
    .C(_03273_),
    .Y(_03274_));
 sg13g2_a21oi_1 _19850_ (.A1(_08614_),
    .A2(net4978),
    .Y(_00292_),
    .B1(_03274_));
 sg13g2_and2_1 _19851_ (.A(\rom_next_addr_in_queue[9] ),
    .B(_03271_),
    .X(_03275_));
 sg13g2_o21ai_1 _19852_ (.B1(net6021),
    .Y(_03276_),
    .A1(\rom_next_addr_in_queue[9] ),
    .A2(_03271_));
 sg13g2_o21ai_1 _19853_ (.B1(_03235_),
    .Y(_03277_),
    .A1(_03275_),
    .A2(_03276_));
 sg13g2_mux2_1 _19854_ (.A0(net7350),
    .A1(_03277_),
    .S(net4975),
    .X(_00293_));
 sg13g2_nand2_1 _19855_ (.Y(_03278_),
    .A(\rom_next_addr_in_queue[10] ),
    .B(_03275_));
 sg13g2_o21ai_1 _19856_ (.B1(net6021),
    .Y(_03279_),
    .A1(net7323),
    .A2(_03275_));
 sg13g2_nor2b_1 _19857_ (.A(_03279_),
    .B_N(_03278_),
    .Y(_03280_));
 sg13g2_nor3_1 _19858_ (.A(net4977),
    .B(_03237_),
    .C(_03280_),
    .Y(_03281_));
 sg13g2_a21oi_1 _19859_ (.A1(_08615_),
    .A2(net4977),
    .Y(_00294_),
    .B1(_03281_));
 sg13g2_xnor2_1 _19860_ (.Y(_03282_),
    .A(net7406),
    .B(_03278_));
 sg13g2_a21oi_1 _19861_ (.A1(net6024),
    .A2(_03282_),
    .Y(_03283_),
    .B1(net4978));
 sg13g2_a22oi_1 _19862_ (.Y(_00295_),
    .B1(_03241_),
    .B2(_03283_),
    .A2(net4977),
    .A1(_08616_));
 sg13g2_nand3_1 _19863_ (.B(net6508),
    .C(net7374),
    .A(net7331),
    .Y(_03284_));
 sg13g2_a21o_1 _19864_ (.A2(net6508),
    .A1(net7331),
    .B1(net7374),
    .X(_03285_));
 sg13g2_nand2_1 _19865_ (.Y(_03286_),
    .A(_03284_),
    .B(_03285_));
 sg13g2_nand2_1 _19866_ (.Y(_03287_),
    .A(net7279),
    .B(\atari2600.tia.audio_l ));
 sg13g2_o21ai_1 _19867_ (.B1(net6572),
    .Y(_03288_),
    .A1(_03286_),
    .A2(_03287_));
 sg13g2_a21oi_1 _19868_ (.A1(_03286_),
    .A2(_03287_),
    .Y(_00296_),
    .B1(_03288_));
 sg13g2_o21ai_1 _19869_ (.B1(_03284_),
    .Y(_03289_),
    .A1(_03286_),
    .A2(_03287_));
 sg13g2_nand2_1 _19870_ (.Y(_03290_),
    .A(net7111),
    .B(\atari2600.tia.audio_l ));
 sg13g2_nand3_1 _19871_ (.B(net6509),
    .C(\audio_pwm_accumulator[1] ),
    .A(\atari2600.tia.audv1[1] ),
    .Y(_03291_));
 sg13g2_a21o_1 _19872_ (.A2(net6509),
    .A1(\atari2600.tia.audv1[1] ),
    .B1(\audio_pwm_accumulator[1] ),
    .X(_03292_));
 sg13g2_nand2_1 _19873_ (.Y(_03293_),
    .A(_03291_),
    .B(_03292_));
 sg13g2_xor2_1 _19874_ (.B(_03293_),
    .A(_03290_),
    .X(_03294_));
 sg13g2_or2_1 _19875_ (.X(_03295_),
    .B(_03294_),
    .A(_03289_));
 sg13g2_nand2_1 _19876_ (.Y(_03296_),
    .A(_03289_),
    .B(_03294_));
 sg13g2_and3_1 _19877_ (.X(_00297_),
    .A(net6572),
    .B(_03295_),
    .C(_03296_));
 sg13g2_nand2_1 _19878_ (.Y(_03297_),
    .A(\atari2600.tia.audv0[2] ),
    .B(\atari2600.tia.audio_l ));
 sg13g2_and3_1 _19879_ (.X(_03298_),
    .A(\atari2600.tia.audv1[2] ),
    .B(net6508),
    .C(\audio_pwm_accumulator[2] ));
 sg13g2_nand3_1 _19880_ (.B(net6508),
    .C(\audio_pwm_accumulator[2] ),
    .A(\atari2600.tia.audv1[2] ),
    .Y(_03299_));
 sg13g2_a21oi_1 _19881_ (.A1(\atari2600.tia.audv1[2] ),
    .A2(net6508),
    .Y(_03300_),
    .B1(\audio_pwm_accumulator[2] ));
 sg13g2_nor2_1 _19882_ (.A(_03298_),
    .B(_03300_),
    .Y(_03301_));
 sg13g2_xnor2_1 _19883_ (.Y(_03302_),
    .A(_03297_),
    .B(_03301_));
 sg13g2_o21ai_1 _19884_ (.B1(_03291_),
    .Y(_03303_),
    .A1(_03290_),
    .A2(_03293_));
 sg13g2_nand2_1 _19885_ (.Y(_03304_),
    .A(_03302_),
    .B(_03303_));
 sg13g2_xnor2_1 _19886_ (.Y(_03305_),
    .A(_03302_),
    .B(_03303_));
 sg13g2_or2_1 _19887_ (.X(_03306_),
    .B(_03305_),
    .A(_03296_));
 sg13g2_nand2_1 _19888_ (.Y(_03307_),
    .A(net6572),
    .B(_03306_));
 sg13g2_a21oi_1 _19889_ (.A1(_03296_),
    .A2(_03305_),
    .Y(_00298_),
    .B1(_03307_));
 sg13g2_nand2_1 _19890_ (.Y(_03308_),
    .A(_03304_),
    .B(_03306_));
 sg13g2_nand2_2 _19891_ (.Y(_03309_),
    .A(\atari2600.tia.audv0[3] ),
    .B(\atari2600.tia.audio_l ));
 sg13g2_and3_1 _19892_ (.X(_03310_),
    .A(\atari2600.tia.audv1[3] ),
    .B(net6508),
    .C(\audio_pwm_accumulator[3] ));
 sg13g2_nand3_1 _19893_ (.B(net6508),
    .C(\audio_pwm_accumulator[3] ),
    .A(\atari2600.tia.audv1[3] ),
    .Y(_03311_));
 sg13g2_a21oi_1 _19894_ (.A1(\atari2600.tia.audv1[3] ),
    .A2(net6508),
    .Y(_03312_),
    .B1(\audio_pwm_accumulator[3] ));
 sg13g2_nor2_1 _19895_ (.A(_03310_),
    .B(_03312_),
    .Y(_03313_));
 sg13g2_xnor2_1 _19896_ (.Y(_03314_),
    .A(_03309_),
    .B(_03313_));
 sg13g2_o21ai_1 _19897_ (.B1(_03299_),
    .Y(_03315_),
    .A1(_03297_),
    .A2(_03300_));
 sg13g2_nand2_1 _19898_ (.Y(_03316_),
    .A(_03314_),
    .B(_03315_));
 sg13g2_xor2_1 _19899_ (.B(_03315_),
    .A(_03314_),
    .X(_03317_));
 sg13g2_nand2_1 _19900_ (.Y(_03318_),
    .A(_03308_),
    .B(_03317_));
 sg13g2_o21ai_1 _19901_ (.B1(net6570),
    .Y(_03319_),
    .A1(_03308_),
    .A2(_03317_));
 sg13g2_nor2b_1 _19902_ (.A(_03319_),
    .B_N(_03318_),
    .Y(_00299_));
 sg13g2_o21ai_1 _19903_ (.B1(_03311_),
    .Y(_03320_),
    .A1(_03309_),
    .A2(_03312_));
 sg13g2_nand2_1 _19904_ (.Y(_03321_),
    .A(net7566),
    .B(_03320_));
 sg13g2_xnor2_1 _19905_ (.Y(_03322_),
    .A(net7566),
    .B(_03320_));
 sg13g2_nand3_1 _19906_ (.B(_03318_),
    .C(_03322_),
    .A(_03316_),
    .Y(_03323_));
 sg13g2_a21o_1 _19907_ (.A2(_03318_),
    .A1(_03316_),
    .B1(_03322_),
    .X(_03324_));
 sg13g2_and3_1 _19908_ (.X(_00300_),
    .A(net6571),
    .B(_03323_),
    .C(_03324_));
 sg13g2_a21oi_2 _19909_ (.B1(net6530),
    .Y(_00301_),
    .A2(_03324_),
    .A1(_03321_));
 sg13g2_nor3_1 _19910_ (.A(net6153),
    .B(net6208),
    .C(net6125),
    .Y(_03325_));
 sg13g2_and4_2 _19911_ (.A(_09226_),
    .B(_09231_),
    .C(_03200_),
    .D(_03325_),
    .X(_03326_));
 sg13g2_nand4_1 _19912_ (.B(_09231_),
    .C(_03200_),
    .A(_09226_),
    .Y(_03327_),
    .D(_03325_));
 sg13g2_xnor2_1 _19913_ (.Y(_03328_),
    .A(\frame_counter[2] ),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_xnor2_1 _19914_ (.Y(_03329_),
    .A(\frame_counter[1] ),
    .B(\hvsync_gen.hpos[0] ));
 sg13g2_nand2_2 _19915_ (.Y(_03330_),
    .A(_03328_),
    .B(_03329_));
 sg13g2_and3_1 _19916_ (.X(_00302_),
    .A(net2988),
    .B(net5981),
    .C(net6017));
 sg13g2_mux4_1 _19917_ (.S0(net6192),
    .A0(\scanline[128][3] ),
    .A1(\scanline[129][3] ),
    .A2(\scanline[130][3] ),
    .A3(\scanline[131][3] ),
    .S1(net6140),
    .X(_03331_));
 sg13g2_nor3_2 _19918_ (.A(net6130),
    .B(net6074),
    .C(_03331_),
    .Y(_03332_));
 sg13g2_nor2_1 _19919_ (.A(_09220_),
    .B(_03332_),
    .Y(_03333_));
 sg13g2_mux4_1 _19920_ (.S0(net6206),
    .A0(\scanline[148][3] ),
    .A1(\scanline[149][3] ),
    .A2(\scanline[150][3] ),
    .A3(\scanline[151][3] ),
    .S1(net6151),
    .X(_03334_));
 sg13g2_nor2_1 _19921_ (.A(net6057),
    .B(_03334_),
    .Y(_03335_));
 sg13g2_mux4_1 _19922_ (.S0(net6203),
    .A0(\scanline[156][3] ),
    .A1(\scanline[157][3] ),
    .A2(\scanline[158][3] ),
    .A3(\scanline[159][3] ),
    .S1(net6148),
    .X(_03336_));
 sg13g2_nor2_1 _19923_ (.A(net6090),
    .B(_03336_),
    .Y(_03337_));
 sg13g2_nor2b_1 _19924_ (.A(net6134),
    .B_N(net6133),
    .Y(_03338_));
 sg13g2_nand2b_1 _19925_ (.Y(_03339_),
    .B(net6133),
    .A_N(net6134));
 sg13g2_mux4_1 _19926_ (.S0(net6206),
    .A0(\scanline[152][3] ),
    .A1(\scanline[153][3] ),
    .A2(\scanline[154][3] ),
    .A3(\scanline[155][3] ),
    .S1(net6151),
    .X(_03340_));
 sg13g2_nor2_1 _19927_ (.A(net6046),
    .B(_03340_),
    .Y(_03341_));
 sg13g2_mux4_1 _19928_ (.S0(net6209),
    .A0(\scanline[144][3] ),
    .A1(\scanline[145][3] ),
    .A2(\scanline[146][3] ),
    .A3(\scanline[147][3] ),
    .S1(net6153),
    .X(_03342_));
 sg13g2_o21ai_1 _19929_ (.B1(net6128),
    .Y(_03343_),
    .A1(net6073),
    .A2(_03342_));
 sg13g2_nor4_1 _19930_ (.A(_03335_),
    .B(_03337_),
    .C(_03341_),
    .D(_03343_),
    .Y(_03344_));
 sg13g2_mux4_1 _19931_ (.S0(net6191),
    .A0(\scanline[136][3] ),
    .A1(\scanline[137][3] ),
    .A2(\scanline[138][3] ),
    .A3(\scanline[139][3] ),
    .S1(net6139),
    .X(_03345_));
 sg13g2_nor2_1 _19932_ (.A(net6044),
    .B(_03345_),
    .Y(_03346_));
 sg13g2_mux4_1 _19933_ (.S0(net6189),
    .A0(\scanline[132][3] ),
    .A1(\scanline[133][3] ),
    .A2(\scanline[134][3] ),
    .A3(\scanline[135][3] ),
    .S1(net6137),
    .X(_03347_));
 sg13g2_nor2_1 _19934_ (.A(net6056),
    .B(_03347_),
    .Y(_03348_));
 sg13g2_mux4_1 _19935_ (.S0(net6203),
    .A0(\scanline[140][3] ),
    .A1(\scanline[141][3] ),
    .A2(\scanline[142][3] ),
    .A3(\scanline[143][3] ),
    .S1(net6148),
    .X(_03349_));
 sg13g2_o21ai_1 _19936_ (.B1(net6117),
    .Y(_03350_),
    .A1(net6090),
    .A2(_03349_));
 sg13g2_nor3_2 _19937_ (.A(_03346_),
    .B(_03348_),
    .C(_03350_),
    .Y(_03351_));
 sg13g2_o21ai_1 _19938_ (.B1(_03333_),
    .Y(_03352_),
    .A1(_03344_),
    .A2(_03351_));
 sg13g2_mux4_1 _19939_ (.S0(net6200),
    .A0(\scanline[60][3] ),
    .A1(\scanline[61][3] ),
    .A2(\scanline[62][3] ),
    .A3(\scanline[63][3] ),
    .S1(net6145),
    .X(_03353_));
 sg13g2_and2_1 _19940_ (.A(net6093),
    .B(_03353_),
    .X(_03354_));
 sg13g2_mux4_1 _19941_ (.S0(net6201),
    .A0(\scanline[52][3] ),
    .A1(\scanline[53][3] ),
    .A2(\scanline[54][3] ),
    .A3(\scanline[55][3] ),
    .S1(net6145),
    .X(_03355_));
 sg13g2_nand2b_1 _19942_ (.Y(_03356_),
    .B(\scanline[56][3] ),
    .A_N(net6199));
 sg13g2_a21oi_1 _19943_ (.A1(net6199),
    .A2(\scanline[57][3] ),
    .Y(_03357_),
    .B1(net6146));
 sg13g2_nand2_1 _19944_ (.Y(_03358_),
    .A(net6209),
    .B(\scanline[59][3] ));
 sg13g2_nand2b_1 _19945_ (.Y(_03359_),
    .B(\scanline[58][3] ),
    .A_N(net6209));
 sg13g2_nand3_1 _19946_ (.B(_03358_),
    .C(_03359_),
    .A(net6153),
    .Y(_03360_));
 sg13g2_a21oi_1 _19947_ (.A1(_03356_),
    .A2(_03357_),
    .Y(_03361_),
    .B1(net6044));
 sg13g2_mux4_1 _19948_ (.S0(net6198),
    .A0(\scanline[48][3] ),
    .A1(\scanline[49][3] ),
    .A2(\scanline[50][3] ),
    .A3(\scanline[51][3] ),
    .S1(net6144),
    .X(_03362_));
 sg13g2_a21oi_2 _19949_ (.B1(net6117),
    .Y(_03363_),
    .A2(_03361_),
    .A1(_03360_));
 sg13g2_a221oi_1 _19950_ (.B2(net6078),
    .C1(_03354_),
    .B1(_03362_),
    .A1(net6060),
    .Y(_03364_),
    .A2(_03355_));
 sg13g2_mux4_1 _19951_ (.S0(net6196),
    .A0(\scanline[40][3] ),
    .A1(\scanline[41][3] ),
    .A2(\scanline[42][3] ),
    .A3(\scanline[43][3] ),
    .S1(net6143),
    .X(_03365_));
 sg13g2_nand2_1 _19952_ (.Y(_03366_),
    .A(net6219),
    .B(\scanline[35][3] ));
 sg13g2_nand2b_1 _19953_ (.Y(_03367_),
    .B(\scanline[34][3] ),
    .A_N(net6216));
 sg13g2_nand3_1 _19954_ (.B(_03366_),
    .C(_03367_),
    .A(net6160),
    .Y(_03368_));
 sg13g2_nand2b_1 _19955_ (.Y(_03369_),
    .B(\scanline[32][3] ),
    .A_N(net6216));
 sg13g2_a21oi_1 _19956_ (.A1(net6215),
    .A2(\scanline[33][3] ),
    .Y(_03370_),
    .B1(net6161));
 sg13g2_a21oi_1 _19957_ (.A1(_03369_),
    .A2(_03370_),
    .Y(_03371_),
    .B1(net6075));
 sg13g2_mux4_1 _19958_ (.S0(net6211),
    .A0(\scanline[36][3] ),
    .A1(\scanline[37][3] ),
    .A2(\scanline[38][3] ),
    .A3(\scanline[39][3] ),
    .S1(net6156),
    .X(_03372_));
 sg13g2_mux4_1 _19959_ (.S0(net6211),
    .A0(\scanline[44][3] ),
    .A1(\scanline[45][3] ),
    .A2(\scanline[46][3] ),
    .A3(\scanline[47][3] ),
    .S1(net6156),
    .X(_03373_));
 sg13g2_a22oi_1 _19960_ (.Y(_03374_),
    .B1(_03373_),
    .B2(net6093),
    .A2(_03365_),
    .A1(net6047));
 sg13g2_a221oi_1 _19961_ (.B2(net6060),
    .C1(net6131),
    .B1(_03372_),
    .A1(_03368_),
    .Y(_03375_),
    .A2(_03371_));
 sg13g2_a221oi_1 _19962_ (.B2(_03375_),
    .C1(net6113),
    .B1(_03374_),
    .A1(_03363_),
    .Y(_03376_),
    .A2(_03364_));
 sg13g2_nand2_1 _19963_ (.Y(_03377_),
    .A(net6131),
    .B(net6114));
 sg13g2_mux4_1 _19964_ (.S0(net6221),
    .A0(\scanline[20][3] ),
    .A1(\scanline[21][3] ),
    .A2(\scanline[22][3] ),
    .A3(\scanline[23][3] ),
    .S1(net6164),
    .X(_03378_));
 sg13g2_mux4_1 _19965_ (.S0(net6213),
    .A0(\scanline[28][3] ),
    .A1(\scanline[29][3] ),
    .A2(\scanline[30][3] ),
    .A3(\scanline[31][3] ),
    .S1(net6158),
    .X(_03379_));
 sg13g2_mux4_1 _19966_ (.S0(net6221),
    .A0(\scanline[24][3] ),
    .A1(\scanline[25][3] ),
    .A2(\scanline[26][3] ),
    .A3(\scanline[27][3] ),
    .S1(net6164),
    .X(_03380_));
 sg13g2_mux4_1 _19967_ (.S0(net6212),
    .A0(\scanline[16][3] ),
    .A1(\scanline[17][3] ),
    .A2(\scanline[18][3] ),
    .A3(\scanline[19][3] ),
    .S1(net6157),
    .X(_03381_));
 sg13g2_a22oi_1 _19968_ (.Y(_03382_),
    .B1(_03381_),
    .B2(net6079),
    .A2(_03379_),
    .A1(net6095));
 sg13g2_a22oi_1 _19969_ (.Y(_03383_),
    .B1(_03380_),
    .B2(net6050),
    .A2(_03378_),
    .A1(net6062));
 sg13g2_a21oi_2 _19970_ (.B1(net6011),
    .Y(_03384_),
    .A2(_03383_),
    .A1(_03382_));
 sg13g2_mux4_1 _19971_ (.S0(net6193),
    .A0(\scanline[8][3] ),
    .A1(\scanline[9][3] ),
    .A2(\scanline[10][3] ),
    .A3(\scanline[11][3] ),
    .S1(net6141),
    .X(_03385_));
 sg13g2_mux4_1 _19972_ (.S0(net6186),
    .A0(\scanline[12][3] ),
    .A1(\scanline[13][3] ),
    .A2(\scanline[14][3] ),
    .A3(\scanline[15][3] ),
    .S1(net6135),
    .X(_03386_));
 sg13g2_mux4_1 _19973_ (.S0(net6193),
    .A0(\scanline[0][3] ),
    .A1(\scanline[1][3] ),
    .A2(\scanline[2][3] ),
    .A3(\scanline[3][3] ),
    .S1(net6141),
    .X(_03387_));
 sg13g2_mux4_1 _19974_ (.S0(net6187),
    .A0(\scanline[4][3] ),
    .A1(\scanline[5][3] ),
    .A2(\scanline[6][3] ),
    .A3(\scanline[7][3] ),
    .S1(net6136),
    .X(_03388_));
 sg13g2_a22oi_1 _19975_ (.Y(_03389_),
    .B1(_03388_),
    .B2(net6059),
    .A2(_03386_),
    .A1(net6094));
 sg13g2_a22oi_1 _19976_ (.Y(_03390_),
    .B1(_03387_),
    .B2(net6076),
    .A2(_03385_),
    .A1(net6048));
 sg13g2_a21oi_2 _19977_ (.B1(net6025),
    .Y(_03391_),
    .A2(_03390_),
    .A1(_03389_));
 sg13g2_or3_2 _19978_ (.A(net6127),
    .B(_03384_),
    .C(_03391_),
    .X(_03392_));
 sg13g2_nand2b_1 _19979_ (.Y(_03393_),
    .B(\scanline[124][3] ),
    .A_N(net6227));
 sg13g2_a21oi_1 _19980_ (.A1(net6224),
    .A2(\scanline[125][3] ),
    .Y(_03394_),
    .B1(net6162));
 sg13g2_nand2_1 _19981_ (.Y(_03395_),
    .A(net6218),
    .B(\scanline[127][3] ));
 sg13g2_nand2b_1 _19982_ (.Y(_03396_),
    .B(\scanline[126][3] ),
    .A_N(net6217));
 sg13g2_nand3_1 _19983_ (.B(_03395_),
    .C(_03396_),
    .A(net6163),
    .Y(_03397_));
 sg13g2_a21oi_1 _19984_ (.A1(_03393_),
    .A2(_03394_),
    .Y(_03398_),
    .B1(net6092));
 sg13g2_mux4_1 _19985_ (.S0(net6233),
    .A0(\scanline[120][3] ),
    .A1(\scanline[121][3] ),
    .A2(\scanline[122][3] ),
    .A3(\scanline[123][3] ),
    .S1(net6175),
    .X(_03399_));
 sg13g2_mux4_1 _19986_ (.S0(net6230),
    .A0(\scanline[112][3] ),
    .A1(\scanline[113][3] ),
    .A2(\scanline[114][3] ),
    .A3(\scanline[115][3] ),
    .S1(net6171),
    .X(_03400_));
 sg13g2_mux4_1 _19987_ (.S0(net6233),
    .A0(\scanline[116][3] ),
    .A1(\scanline[117][3] ),
    .A2(\scanline[118][3] ),
    .A3(\scanline[119][3] ),
    .S1(net6175),
    .X(_03401_));
 sg13g2_a22oi_1 _19988_ (.Y(_03402_),
    .B1(_03401_),
    .B2(net6065),
    .A2(_03399_),
    .A1(net6049));
 sg13g2_a221oi_1 _19989_ (.B2(net6080),
    .C1(net6116),
    .B1(_03400_),
    .A1(_03397_),
    .Y(_03403_),
    .A2(_03398_));
 sg13g2_nand2b_1 _19990_ (.Y(_03404_),
    .B(\scanline[100][3] ),
    .A_N(net6230));
 sg13g2_a21oi_1 _19991_ (.A1(net6229),
    .A2(\scanline[101][3] ),
    .Y(_03405_),
    .B1(net6172));
 sg13g2_nand2_1 _19992_ (.Y(_03406_),
    .A(net6229),
    .B(\scanline[103][3] ));
 sg13g2_nand2b_1 _19993_ (.Y(_03407_),
    .B(\scanline[102][3] ),
    .A_N(net6229));
 sg13g2_nand3_1 _19994_ (.B(_03406_),
    .C(_03407_),
    .A(net6172),
    .Y(_03408_));
 sg13g2_a21oi_1 _19995_ (.A1(_03404_),
    .A2(_03405_),
    .Y(_03409_),
    .B1(net6058));
 sg13g2_a21oi_1 _19996_ (.A1(_03408_),
    .A2(_03409_),
    .Y(_03410_),
    .B1(net6132));
 sg13g2_mux4_1 _19997_ (.S0(net6234),
    .A0(\scanline[104][3] ),
    .A1(\scanline[105][3] ),
    .A2(\scanline[106][3] ),
    .A3(\scanline[107][3] ),
    .S1(net6176),
    .X(_03411_));
 sg13g2_mux4_1 _19998_ (.S0(net6234),
    .A0(\scanline[108][3] ),
    .A1(\scanline[109][3] ),
    .A2(\scanline[110][3] ),
    .A3(\scanline[111][3] ),
    .S1(net6176),
    .X(_03412_));
 sg13g2_mux4_1 _19999_ (.S0(net6238),
    .A0(\scanline[96][3] ),
    .A1(\scanline[97][3] ),
    .A2(\scanline[98][3] ),
    .A3(\scanline[99][3] ),
    .S1(net6178),
    .X(_03413_));
 sg13g2_and2_1 _20000_ (.A(net6081),
    .B(_03413_),
    .X(_03414_));
 sg13g2_a221oi_1 _20001_ (.B2(net6099),
    .C1(_03414_),
    .B1(_03412_),
    .A1(net6053),
    .Y(_03415_),
    .A2(_03411_));
 sg13g2_a221oi_1 _20002_ (.B2(_03415_),
    .C1(net6114),
    .B1(_03410_),
    .A1(_03402_),
    .Y(_03416_),
    .A2(_03403_));
 sg13g2_mux4_1 _20003_ (.S0(net6222),
    .A0(\scanline[68][3] ),
    .A1(\scanline[69][3] ),
    .A2(\scanline[70][3] ),
    .A3(\scanline[71][3] ),
    .S1(net6165),
    .X(_03417_));
 sg13g2_mux4_1 _20004_ (.S0(net6224),
    .A0(\scanline[76][3] ),
    .A1(\scanline[77][3] ),
    .A2(\scanline[78][3] ),
    .A3(\scanline[79][3] ),
    .S1(net6169),
    .X(_03418_));
 sg13g2_mux4_1 _20005_ (.S0(net6222),
    .A0(\scanline[72][3] ),
    .A1(\scanline[73][3] ),
    .A2(\scanline[74][3] ),
    .A3(\scanline[75][3] ),
    .S1(net6165),
    .X(_03419_));
 sg13g2_mux4_1 _20006_ (.S0(net6225),
    .A0(\scanline[64][3] ),
    .A1(\scanline[65][3] ),
    .A2(\scanline[66][3] ),
    .A3(\scanline[67][3] ),
    .S1(net6168),
    .X(_03420_));
 sg13g2_a22oi_1 _20007_ (.Y(_03421_),
    .B1(_03420_),
    .B2(net6081),
    .A2(_03418_),
    .A1(net6097));
 sg13g2_a22oi_1 _20008_ (.Y(_03422_),
    .B1(_03419_),
    .B2(net6050),
    .A2(_03417_),
    .A1(net6062));
 sg13g2_a21oi_2 _20009_ (.B1(net6026),
    .Y(_03423_),
    .A2(_03422_),
    .A1(_03421_));
 sg13g2_mux4_1 _20010_ (.S0(net6239),
    .A0(\scanline[80][3] ),
    .A1(\scanline[81][3] ),
    .A2(\scanline[82][3] ),
    .A3(\scanline[83][3] ),
    .S1(net6179),
    .X(_03424_));
 sg13g2_mux4_1 _20011_ (.S0(net6240),
    .A0(\scanline[92][3] ),
    .A1(\scanline[93][3] ),
    .A2(\scanline[94][3] ),
    .A3(\scanline[95][3] ),
    .S1(net6181),
    .X(_03425_));
 sg13g2_mux4_1 _20012_ (.S0(net6240),
    .A0(\scanline[84][3] ),
    .A1(\scanline[85][3] ),
    .A2(\scanline[86][3] ),
    .A3(\scanline[87][3] ),
    .S1(net6183),
    .X(_03426_));
 sg13g2_mux4_1 _20013_ (.S0(net6242),
    .A0(\scanline[88][3] ),
    .A1(\scanline[89][3] ),
    .A2(\scanline[90][3] ),
    .A3(\scanline[91][3] ),
    .S1(net6183),
    .X(_03427_));
 sg13g2_a22oi_1 _20014_ (.Y(_03428_),
    .B1(_03427_),
    .B2(net6054),
    .A2(_03425_),
    .A1(net6098));
 sg13g2_a22oi_1 _20015_ (.Y(_03429_),
    .B1(_03426_),
    .B2(net6066),
    .A2(_03424_),
    .A1(net6082));
 sg13g2_a21oi_1 _20016_ (.A1(_03428_),
    .A2(_03429_),
    .Y(_03430_),
    .B1(net6012));
 sg13g2_nor4_2 _20017_ (.A(_08656_),
    .B(_03416_),
    .C(_03423_),
    .Y(_03431_),
    .D(_03430_));
 sg13g2_o21ai_1 _20018_ (.B1(_08655_),
    .Y(_03432_),
    .A1(_03376_),
    .A2(_03392_));
 sg13g2_or2_1 _20019_ (.X(_03433_),
    .B(_03432_),
    .A(_03431_));
 sg13g2_o21ai_1 _20020_ (.B1(_03352_),
    .Y(_03434_),
    .A1(_03431_),
    .A2(_03432_));
 sg13g2_and2_1 _20021_ (.A(net6086),
    .B(_03434_),
    .X(_03435_));
 sg13g2_nand2_1 _20022_ (.Y(_03436_),
    .A(net6086),
    .B(_03434_));
 sg13g2_mux4_1 _20023_ (.S0(net6239),
    .A0(\scanline[80][1] ),
    .A1(\scanline[81][1] ),
    .A2(\scanline[82][1] ),
    .A3(\scanline[83][1] ),
    .S1(net6179),
    .X(_03437_));
 sg13g2_mux4_1 _20024_ (.S0(net6234),
    .A0(\scanline[84][1] ),
    .A1(\scanline[85][1] ),
    .A2(\scanline[86][1] ),
    .A3(\scanline[87][1] ),
    .S1(net6176),
    .X(_03438_));
 sg13g2_mux4_1 _20025_ (.S0(net6238),
    .A0(\scanline[92][1] ),
    .A1(\scanline[93][1] ),
    .A2(\scanline[94][1] ),
    .A3(\scanline[95][1] ),
    .S1(net6178),
    .X(_03439_));
 sg13g2_mux4_1 _20026_ (.S0(net6240),
    .A0(\scanline[88][1] ),
    .A1(\scanline[89][1] ),
    .A2(\scanline[90][1] ),
    .A3(\scanline[91][1] ),
    .S1(net6181),
    .X(_03440_));
 sg13g2_a22oi_1 _20027_ (.Y(_03441_),
    .B1(_03440_),
    .B2(net6052),
    .A2(_03438_),
    .A1(net6064));
 sg13g2_a22oi_1 _20028_ (.Y(_03442_),
    .B1(_03439_),
    .B2(net6098),
    .A2(_03437_),
    .A1(net6082));
 sg13g2_a21oi_1 _20029_ (.A1(_03441_),
    .A2(_03442_),
    .Y(_03443_),
    .B1(net6012));
 sg13g2_nand2_2 _20030_ (.Y(_03444_),
    .A(net6116),
    .B(\hvsync_gen.hpos[7] ));
 sg13g2_mux4_1 _20031_ (.S0(net6238),
    .A0(\scanline[108][1] ),
    .A1(\scanline[109][1] ),
    .A2(\scanline[110][1] ),
    .A3(\scanline[111][1] ),
    .S1(net6180),
    .X(_03445_));
 sg13g2_mux4_1 _20032_ (.S0(net6237),
    .A0(\scanline[96][1] ),
    .A1(\scanline[97][1] ),
    .A2(\scanline[98][1] ),
    .A3(\scanline[99][1] ),
    .S1(net6178),
    .X(_03446_));
 sg13g2_a22oi_1 _20033_ (.Y(_03447_),
    .B1(_03446_),
    .B2(net6080),
    .A2(_03445_),
    .A1(net6097));
 sg13g2_mux4_1 _20034_ (.S0(net6234),
    .A0(\scanline[104][1] ),
    .A1(\scanline[105][1] ),
    .A2(\scanline[106][1] ),
    .A3(\scanline[107][1] ),
    .S1(net6176),
    .X(_03448_));
 sg13g2_mux4_1 _20035_ (.S0(net6230),
    .A0(\scanline[100][1] ),
    .A1(\scanline[101][1] ),
    .A2(\scanline[102][1] ),
    .A3(\scanline[103][1] ),
    .S1(net6171),
    .X(_03449_));
 sg13g2_a22oi_1 _20036_ (.Y(_03450_),
    .B1(_03449_),
    .B2(net6064),
    .A2(_03448_),
    .A1(net6052));
 sg13g2_a21oi_1 _20037_ (.A1(_03447_),
    .A2(_03450_),
    .Y(_03451_),
    .B1(_03444_));
 sg13g2_mux4_1 _20038_ (.S0(net6222),
    .A0(\scanline[68][1] ),
    .A1(\scanline[69][1] ),
    .A2(\scanline[70][1] ),
    .A3(\scanline[71][1] ),
    .S1(net6165),
    .X(_03452_));
 sg13g2_mux4_1 _20039_ (.S0(net6224),
    .A0(\scanline[76][1] ),
    .A1(\scanline[77][1] ),
    .A2(\scanline[78][1] ),
    .A3(\scanline[79][1] ),
    .S1(net6169),
    .X(_03453_));
 sg13g2_mux4_1 _20040_ (.S0(net6223),
    .A0(\scanline[72][1] ),
    .A1(\scanline[73][1] ),
    .A2(\scanline[74][1] ),
    .A3(\scanline[75][1] ),
    .S1(net6166),
    .X(_03454_));
 sg13g2_mux4_1 _20041_ (.S0(net6226),
    .A0(\scanline[64][1] ),
    .A1(\scanline[65][1] ),
    .A2(\scanline[66][1] ),
    .A3(\scanline[67][1] ),
    .S1(net6168),
    .X(_03455_));
 sg13g2_a22oi_1 _20042_ (.Y(_03456_),
    .B1(_03455_),
    .B2(net6081),
    .A2(_03453_),
    .A1(net6096));
 sg13g2_a22oi_1 _20043_ (.Y(_03457_),
    .B1(_03454_),
    .B2(net6050),
    .A2(_03452_),
    .A1(net6062));
 sg13g2_a21oi_2 _20044_ (.B1(net6026),
    .Y(_03458_),
    .A2(_03457_),
    .A1(_03456_));
 sg13g2_mux4_1 _20045_ (.S0(net6231),
    .A0(\scanline[116][1] ),
    .A1(\scanline[117][1] ),
    .A2(\scanline[118][1] ),
    .A3(\scanline[119][1] ),
    .S1(net6173),
    .X(_03459_));
 sg13g2_mux4_1 _20046_ (.S0(net6233),
    .A0(\scanline[120][1] ),
    .A1(\scanline[121][1] ),
    .A2(\scanline[122][1] ),
    .A3(\scanline[123][1] ),
    .S1(net6175),
    .X(_03460_));
 sg13g2_a22oi_1 _20047_ (.Y(_03461_),
    .B1(_03460_),
    .B2(net6049),
    .A2(_03459_),
    .A1(net6065));
 sg13g2_mux4_1 _20048_ (.S0(net6219),
    .A0(\scanline[124][1] ),
    .A1(\scanline[125][1] ),
    .A2(\scanline[126][1] ),
    .A3(\scanline[127][1] ),
    .S1(net6163),
    .X(_03462_));
 sg13g2_mux4_1 _20049_ (.S0(net6231),
    .A0(\scanline[112][1] ),
    .A1(\scanline[113][1] ),
    .A2(\scanline[114][1] ),
    .A3(\scanline[115][1] ),
    .S1(net6173),
    .X(_03463_));
 sg13g2_a22oi_1 _20050_ (.Y(_03464_),
    .B1(_03463_),
    .B2(net6078),
    .A2(_03462_),
    .A1(net6099));
 sg13g2_a21oi_1 _20051_ (.A1(_03461_),
    .A2(_03464_),
    .Y(_03465_),
    .B1(_09223_));
 sg13g2_or4_2 _20052_ (.A(_03443_),
    .B(_03451_),
    .C(_03458_),
    .D(_03465_),
    .X(_03466_));
 sg13g2_mux4_1 _20053_ (.S0(net6215),
    .A0(\scanline[32][1] ),
    .A1(\scanline[33][1] ),
    .A2(\scanline[34][1] ),
    .A3(\scanline[35][1] ),
    .S1(net6161),
    .X(_03467_));
 sg13g2_mux4_1 _20054_ (.S0(net6195),
    .A0(\scanline[40][1] ),
    .A1(\scanline[41][1] ),
    .A2(\scanline[42][1] ),
    .A3(\scanline[43][1] ),
    .S1(net6142),
    .X(_03468_));
 sg13g2_mux4_1 _20055_ (.S0(net6216),
    .A0(\scanline[44][1] ),
    .A1(\scanline[45][1] ),
    .A2(\scanline[46][1] ),
    .A3(\scanline[47][1] ),
    .S1(net6161),
    .X(_03469_));
 sg13g2_mux4_1 _20056_ (.S0(net6211),
    .A0(\scanline[36][1] ),
    .A1(\scanline[37][1] ),
    .A2(\scanline[38][1] ),
    .A3(\scanline[39][1] ),
    .S1(net6156),
    .X(_03470_));
 sg13g2_a22oi_1 _20057_ (.Y(_03471_),
    .B1(_03470_),
    .B2(net6063),
    .A2(_03468_),
    .A1(net6047));
 sg13g2_a22oi_1 _20058_ (.Y(_03472_),
    .B1(_03469_),
    .B2(net6099),
    .A2(_03467_),
    .A1(net6078));
 sg13g2_a21o_1 _20059_ (.A2(_03472_),
    .A1(_03471_),
    .B1(_03444_),
    .X(_03473_));
 sg13g2_mux4_1 _20060_ (.S0(net6200),
    .A0(\scanline[60][1] ),
    .A1(\scanline[61][1] ),
    .A2(\scanline[62][1] ),
    .A3(\scanline[63][1] ),
    .S1(net6145),
    .X(_03474_));
 sg13g2_mux4_1 _20061_ (.S0(net6208),
    .A0(\scanline[52][1] ),
    .A1(\scanline[53][1] ),
    .A2(\scanline[54][1] ),
    .A3(\scanline[55][1] ),
    .S1(net6154),
    .X(_03475_));
 sg13g2_a22oi_1 _20062_ (.Y(_03476_),
    .B1(_03475_),
    .B2(net6061),
    .A2(_03474_),
    .A1(net6101));
 sg13g2_mux4_1 _20063_ (.S0(net6199),
    .A0(\scanline[56][1] ),
    .A1(\scanline[57][1] ),
    .A2(\scanline[58][1] ),
    .A3(\scanline[59][1] ),
    .S1(net6144),
    .X(_03477_));
 sg13g2_mux4_1 _20064_ (.S0(net6199),
    .A0(\scanline[48][1] ),
    .A1(\scanline[49][1] ),
    .A2(\scanline[50][1] ),
    .A3(\scanline[51][1] ),
    .S1(net6146),
    .X(_03478_));
 sg13g2_a22oi_1 _20065_ (.Y(_03479_),
    .B1(_03478_),
    .B2(net6078),
    .A2(_03477_),
    .A1(net6048));
 sg13g2_a21o_1 _20066_ (.A2(_03479_),
    .A1(_03476_),
    .B1(_09223_),
    .X(_03480_));
 sg13g2_a21oi_1 _20067_ (.A1(_03473_),
    .A2(_03480_),
    .Y(_03481_),
    .B1(net6126));
 sg13g2_nor2b_1 _20068_ (.A(net6187),
    .B_N(\scanline[8][1] ),
    .Y(_03482_));
 sg13g2_a21oi_1 _20069_ (.A1(net6187),
    .A2(\scanline[9][1] ),
    .Y(_03483_),
    .B1(_03482_));
 sg13g2_nand2b_1 _20070_ (.Y(_03484_),
    .B(\scanline[10][1] ),
    .A_N(net6193));
 sg13g2_a21oi_1 _20071_ (.A1(net6193),
    .A2(\scanline[11][1] ),
    .Y(_03485_),
    .B1(_08652_));
 sg13g2_a221oi_1 _20072_ (.B2(_03485_),
    .C1(net6045),
    .B1(_03484_),
    .A1(_08652_),
    .Y(_03486_),
    .A2(_03483_));
 sg13g2_mux4_1 _20073_ (.S0(net6187),
    .A0(\scanline[0][1] ),
    .A1(\scanline[1][1] ),
    .A2(\scanline[2][1] ),
    .A3(\scanline[3][1] ),
    .S1(net6136),
    .X(_03487_));
 sg13g2_mux4_1 _20074_ (.S0(net6189),
    .A0(\scanline[12][1] ),
    .A1(\scanline[13][1] ),
    .A2(\scanline[14][1] ),
    .A3(\scanline[15][1] ),
    .S1(net6137),
    .X(_03488_));
 sg13g2_nand2_1 _20075_ (.Y(_03489_),
    .A(net6094),
    .B(_03488_));
 sg13g2_mux4_1 _20076_ (.S0(net6188),
    .A0(\scanline[4][1] ),
    .A1(\scanline[5][1] ),
    .A2(\scanline[6][1] ),
    .A3(\scanline[7][1] ),
    .S1(net6136),
    .X(_03490_));
 sg13g2_a221oi_1 _20077_ (.B2(net6059),
    .C1(net6130),
    .B1(_03490_),
    .A1(net6076),
    .Y(_03491_),
    .A2(_03487_));
 sg13g2_nand3b_1 _20078_ (.B(_03489_),
    .C(_03491_),
    .Y(_03492_),
    .A_N(_03486_));
 sg13g2_mux4_1 _20079_ (.S0(net6224),
    .A0(\scanline[24][1] ),
    .A1(\scanline[25][1] ),
    .A2(\scanline[26][1] ),
    .A3(\scanline[27][1] ),
    .S1(net6169),
    .X(_03493_));
 sg13g2_a21oi_1 _20080_ (.A1(net6051),
    .A2(_03493_),
    .Y(_03494_),
    .B1(net6116));
 sg13g2_mux4_1 _20081_ (.S0(net6212),
    .A0(\scanline[20][1] ),
    .A1(\scanline[21][1] ),
    .A2(\scanline[22][1] ),
    .A3(\scanline[23][1] ),
    .S1(net6157),
    .X(_03495_));
 sg13g2_mux4_1 _20082_ (.S0(net6220),
    .A0(\scanline[28][1] ),
    .A1(\scanline[29][1] ),
    .A2(\scanline[30][1] ),
    .A3(\scanline[31][1] ),
    .S1(net6162),
    .X(_03496_));
 sg13g2_mux4_1 _20083_ (.S0(net6212),
    .A0(\scanline[16][1] ),
    .A1(\scanline[17][1] ),
    .A2(\scanline[18][1] ),
    .A3(\scanline[19][1] ),
    .S1(net6157),
    .X(_03497_));
 sg13g2_nand2_1 _20084_ (.Y(_03498_),
    .A(net6079),
    .B(_03497_));
 sg13g2_a22oi_1 _20085_ (.Y(_03499_),
    .B1(_03496_),
    .B2(net6095),
    .A2(_03495_),
    .A1(net6063));
 sg13g2_nand3_1 _20086_ (.B(_03498_),
    .C(_03499_),
    .A(_03494_),
    .Y(_03500_));
 sg13g2_and2_1 _20087_ (.A(_09226_),
    .B(_03500_),
    .X(_03501_));
 sg13g2_a221oi_1 _20088_ (.B2(_03501_),
    .C1(_03481_),
    .B1(_03492_),
    .A1(net6126),
    .Y(_03502_),
    .A2(_03466_));
 sg13g2_mux4_1 _20089_ (.S0(net6190),
    .A0(\scanline[132][1] ),
    .A1(\scanline[133][1] ),
    .A2(\scanline[134][1] ),
    .A3(\scanline[135][1] ),
    .S1(net6138),
    .X(_03503_));
 sg13g2_nor2_1 _20090_ (.A(net6056),
    .B(_03503_),
    .Y(_03504_));
 sg13g2_mux4_1 _20091_ (.S0(net6192),
    .A0(\scanline[128][1] ),
    .A1(\scanline[129][1] ),
    .A2(\scanline[130][1] ),
    .A3(\scanline[131][1] ),
    .S1(net6140),
    .X(_03505_));
 sg13g2_nor2_1 _20092_ (.A(net6074),
    .B(_03505_),
    .Y(_03506_));
 sg13g2_mux4_1 _20093_ (.S0(net6192),
    .A0(\scanline[136][1] ),
    .A1(\scanline[137][1] ),
    .A2(\scanline[138][1] ),
    .A3(\scanline[139][1] ),
    .S1(net6140),
    .X(_03507_));
 sg13g2_mux4_1 _20094_ (.S0(net6190),
    .A0(\scanline[140][1] ),
    .A1(\scanline[141][1] ),
    .A2(\scanline[142][1] ),
    .A3(\scanline[143][1] ),
    .S1(net6138),
    .X(_03508_));
 sg13g2_nor2_1 _20095_ (.A(net6091),
    .B(_03508_),
    .Y(_03509_));
 sg13g2_o21ai_1 _20096_ (.B1(net6117),
    .Y(_03510_),
    .A1(net6044),
    .A2(_03507_));
 sg13g2_nor4_2 _20097_ (.A(_03504_),
    .B(_03506_),
    .C(_03509_),
    .Y(_03511_),
    .D(_03510_));
 sg13g2_mux4_1 _20098_ (.S0(net6205),
    .A0(\scanline[152][1] ),
    .A1(\scanline[153][1] ),
    .A2(\scanline[154][1] ),
    .A3(\scanline[155][1] ),
    .S1(net6149),
    .X(_03512_));
 sg13g2_o21ai_1 _20099_ (.B1(net6128),
    .Y(_03513_),
    .A1(net6045),
    .A2(_03512_));
 sg13g2_mux4_1 _20100_ (.S0(net6204),
    .A0(\scanline[144][1] ),
    .A1(\scanline[145][1] ),
    .A2(\scanline[146][1] ),
    .A3(\scanline[147][1] ),
    .S1(net6149),
    .X(_03514_));
 sg13g2_nor2_1 _20101_ (.A(net6073),
    .B(_03514_),
    .Y(_03515_));
 sg13g2_mux4_1 _20102_ (.S0(net6207),
    .A0(\scanline[148][1] ),
    .A1(\scanline[149][1] ),
    .A2(\scanline[150][1] ),
    .A3(\scanline[151][1] ),
    .S1(net6152),
    .X(_03516_));
 sg13g2_nor2_1 _20103_ (.A(net6057),
    .B(_03516_),
    .Y(_03517_));
 sg13g2_mux2_1 _20104_ (.A0(\scanline[158][1] ),
    .A1(\scanline[159][1] ),
    .S(net6203),
    .X(_03518_));
 sg13g2_or2_1 _20105_ (.X(_03519_),
    .B(\scanline[156][1] ),
    .A(net6205));
 sg13g2_a21oi_1 _20106_ (.A1(net6205),
    .A2(_08671_),
    .Y(_03520_),
    .B1(net6148));
 sg13g2_a221oi_1 _20107_ (.B2(_03520_),
    .C1(net6090),
    .B1(_03519_),
    .A1(net6150),
    .Y(_03521_),
    .A2(_03518_));
 sg13g2_nor4_1 _20108_ (.A(_03513_),
    .B(_03515_),
    .C(_03517_),
    .D(_03521_),
    .Y(_03522_));
 sg13g2_o21ai_1 _20109_ (.B1(_09219_),
    .Y(_03523_),
    .A1(_03511_),
    .A2(_03522_));
 sg13g2_o21ai_1 _20110_ (.B1(_03523_),
    .Y(_03524_),
    .A1(net6125),
    .A2(_03502_));
 sg13g2_mux4_1 _20111_ (.S0(net6207),
    .A0(\scanline[148][2] ),
    .A1(\scanline[149][2] ),
    .A2(\scanline[150][2] ),
    .A3(\scanline[151][2] ),
    .S1(net6152),
    .X(_03525_));
 sg13g2_o21ai_1 _20112_ (.B1(net6128),
    .Y(_03526_),
    .A1(net6057),
    .A2(_03525_));
 sg13g2_mux4_1 _20113_ (.S0(net6205),
    .A0(\scanline[152][2] ),
    .A1(\scanline[153][2] ),
    .A2(\scanline[154][2] ),
    .A3(\scanline[155][2] ),
    .S1(net6150),
    .X(_03527_));
 sg13g2_nor2_1 _20114_ (.A(net6045),
    .B(_03527_),
    .Y(_03528_));
 sg13g2_mux4_1 _20115_ (.S0(net6203),
    .A0(\scanline[156][2] ),
    .A1(\scanline[157][2] ),
    .A2(\scanline[158][2] ),
    .A3(\scanline[159][2] ),
    .S1(net6148),
    .X(_03529_));
 sg13g2_nor2_1 _20116_ (.A(net6090),
    .B(_03529_),
    .Y(_03530_));
 sg13g2_mux4_1 _20117_ (.S0(net6204),
    .A0(\scanline[144][2] ),
    .A1(\scanline[145][2] ),
    .A2(\scanline[146][2] ),
    .A3(\scanline[147][2] ),
    .S1(net6149),
    .X(_03531_));
 sg13g2_nor2_1 _20118_ (.A(net6073),
    .B(_03531_),
    .Y(_03532_));
 sg13g2_nor4_1 _20119_ (.A(_03526_),
    .B(_03528_),
    .C(_03530_),
    .D(_03532_),
    .Y(_03533_));
 sg13g2_mux4_1 _20120_ (.S0(net6192),
    .A0(\scanline[128][2] ),
    .A1(\scanline[129][2] ),
    .A2(\scanline[130][2] ),
    .A3(\scanline[131][2] ),
    .S1(net6140),
    .X(_03534_));
 sg13g2_o21ai_1 _20121_ (.B1(net6117),
    .Y(_03535_),
    .A1(net6074),
    .A2(_03534_));
 sg13g2_mux4_1 _20122_ (.S0(net6191),
    .A0(\scanline[140][2] ),
    .A1(\scanline[141][2] ),
    .A2(\scanline[142][2] ),
    .A3(\scanline[143][2] ),
    .S1(net6139),
    .X(_03536_));
 sg13g2_nor2_1 _20123_ (.A(net6091),
    .B(_03536_),
    .Y(_03537_));
 sg13g2_mux4_1 _20124_ (.S0(net6191),
    .A0(\scanline[136][2] ),
    .A1(\scanline[137][2] ),
    .A2(\scanline[138][2] ),
    .A3(\scanline[139][2] ),
    .S1(net6139),
    .X(_03538_));
 sg13g2_nor2_1 _20125_ (.A(net6044),
    .B(_03538_),
    .Y(_03539_));
 sg13g2_mux4_1 _20126_ (.S0(net6190),
    .A0(\scanline[132][2] ),
    .A1(\scanline[133][2] ),
    .A2(\scanline[134][2] ),
    .A3(\scanline[135][2] ),
    .S1(net6138),
    .X(_03540_));
 sg13g2_nor2_1 _20127_ (.A(net6056),
    .B(_03540_),
    .Y(_03541_));
 sg13g2_nor4_2 _20128_ (.A(_03535_),
    .B(_03537_),
    .C(_03539_),
    .Y(_03542_),
    .D(_03541_));
 sg13g2_o21ai_1 _20129_ (.B1(_09219_),
    .Y(_03543_),
    .A1(_03533_),
    .A2(_03542_));
 sg13g2_mux4_1 _20130_ (.S0(net6215),
    .A0(\scanline[44][2] ),
    .A1(\scanline[45][2] ),
    .A2(\scanline[46][2] ),
    .A3(\scanline[47][2] ),
    .S1(net6160),
    .X(_03544_));
 sg13g2_mux4_1 _20131_ (.S0(net6211),
    .A0(\scanline[36][2] ),
    .A1(\scanline[37][2] ),
    .A2(\scanline[38][2] ),
    .A3(\scanline[39][2] ),
    .S1(net6156),
    .X(_03545_));
 sg13g2_mux4_1 _20132_ (.S0(net6215),
    .A0(\scanline[32][2] ),
    .A1(\scanline[33][2] ),
    .A2(\scanline[34][2] ),
    .A3(\scanline[35][2] ),
    .S1(net6160),
    .X(_03546_));
 sg13g2_mux4_1 _20133_ (.S0(net6195),
    .A0(\scanline[40][2] ),
    .A1(\scanline[41][2] ),
    .A2(\scanline[42][2] ),
    .A3(\scanline[43][2] ),
    .S1(net6142),
    .X(_03547_));
 sg13g2_a22oi_1 _20134_ (.Y(_03548_),
    .B1(_03547_),
    .B2(net6047),
    .A2(_03545_),
    .A1(net6060));
 sg13g2_a221oi_1 _20135_ (.B2(net6077),
    .C1(net6131),
    .B1(_03546_),
    .A1(net6093),
    .Y(_03549_),
    .A2(_03544_));
 sg13g2_nand2b_1 _20136_ (.Y(_03550_),
    .B(\scanline[48][2] ),
    .A_N(net6198));
 sg13g2_a21oi_1 _20137_ (.A1(net6198),
    .A2(\scanline[49][2] ),
    .Y(_03551_),
    .B1(net6144));
 sg13g2_nand2_1 _20138_ (.Y(_03552_),
    .A(net6198),
    .B(\scanline[51][2] ));
 sg13g2_nand2b_1 _20139_ (.Y(_03553_),
    .B(\scanline[50][2] ),
    .A_N(net6194));
 sg13g2_nand3_1 _20140_ (.B(_03552_),
    .C(_03553_),
    .A(net6144),
    .Y(_03554_));
 sg13g2_a21oi_1 _20141_ (.A1(_03550_),
    .A2(_03551_),
    .Y(_03555_),
    .B1(net6075));
 sg13g2_mux4_1 _20142_ (.S0(net6208),
    .A0(\scanline[52][2] ),
    .A1(\scanline[53][2] ),
    .A2(\scanline[54][2] ),
    .A3(\scanline[55][2] ),
    .S1(net6154),
    .X(_03556_));
 sg13g2_mux4_1 _20143_ (.S0(net6193),
    .A0(\scanline[60][2] ),
    .A1(\scanline[61][2] ),
    .A2(\scanline[62][2] ),
    .A3(\scanline[63][2] ),
    .S1(net6141),
    .X(_03557_));
 sg13g2_mux4_1 _20144_ (.S0(net6208),
    .A0(\scanline[56][2] ),
    .A1(\scanline[57][2] ),
    .A2(\scanline[58][2] ),
    .A3(\scanline[59][2] ),
    .S1(net6153),
    .X(_03558_));
 sg13g2_a22oi_1 _20145_ (.Y(_03559_),
    .B1(_03557_),
    .B2(net6093),
    .A2(_03555_),
    .A1(_03554_));
 sg13g2_a221oi_1 _20146_ (.B2(net6049),
    .C1(net6115),
    .B1(_03558_),
    .A1(net6061),
    .Y(_03560_),
    .A2(_03556_));
 sg13g2_a221oi_1 _20147_ (.B2(_03560_),
    .C1(net6113),
    .B1(_03559_),
    .A1(_03548_),
    .Y(_03561_),
    .A2(_03549_));
 sg13g2_mux4_1 _20148_ (.S0(net6212),
    .A0(\scanline[16][2] ),
    .A1(\scanline[17][2] ),
    .A2(\scanline[18][2] ),
    .A3(\scanline[19][2] ),
    .S1(net6157),
    .X(_03562_));
 sg13g2_mux4_1 _20149_ (.S0(net6213),
    .A0(\scanline[28][2] ),
    .A1(\scanline[29][2] ),
    .A2(\scanline[30][2] ),
    .A3(\scanline[31][2] ),
    .S1(net6158),
    .X(_03563_));
 sg13g2_a22oi_1 _20150_ (.Y(_03564_),
    .B1(_03563_),
    .B2(net6095),
    .A2(_03562_),
    .A1(net6079));
 sg13g2_mux4_1 _20151_ (.S0(net6221),
    .A0(\scanline[24][2] ),
    .A1(\scanline[25][2] ),
    .A2(\scanline[26][2] ),
    .A3(\scanline[27][2] ),
    .S1(net6164),
    .X(_03565_));
 sg13g2_mux4_1 _20152_ (.S0(net6221),
    .A0(\scanline[20][2] ),
    .A1(\scanline[21][2] ),
    .A2(\scanline[22][2] ),
    .A3(\scanline[23][2] ),
    .S1(net6164),
    .X(_03566_));
 sg13g2_a22oi_1 _20153_ (.Y(_03567_),
    .B1(_03566_),
    .B2(net6062),
    .A2(_03565_),
    .A1(net6050));
 sg13g2_a21oi_2 _20154_ (.B1(net6011),
    .Y(_03568_),
    .A2(_03567_),
    .A1(_03564_));
 sg13g2_mux4_1 _20155_ (.S0(net6193),
    .A0(\scanline[0][2] ),
    .A1(\scanline[1][2] ),
    .A2(\scanline[2][2] ),
    .A3(\scanline[3][2] ),
    .S1(net6141),
    .X(_03569_));
 sg13g2_mux4_1 _20156_ (.S0(net6188),
    .A0(\scanline[8][2] ),
    .A1(\scanline[9][2] ),
    .A2(\scanline[10][2] ),
    .A3(\scanline[11][2] ),
    .S1(net6136),
    .X(_03570_));
 sg13g2_mux4_1 _20157_ (.S0(net6187),
    .A0(\scanline[4][2] ),
    .A1(\scanline[5][2] ),
    .A2(\scanline[6][2] ),
    .A3(\scanline[7][2] ),
    .S1(net6136),
    .X(_03571_));
 sg13g2_mux4_1 _20158_ (.S0(net6189),
    .A0(\scanline[12][2] ),
    .A1(\scanline[13][2] ),
    .A2(\scanline[14][2] ),
    .A3(\scanline[15][2] ),
    .S1(net6137),
    .X(_03572_));
 sg13g2_a22oi_1 _20159_ (.Y(_03573_),
    .B1(_03572_),
    .B2(net6094),
    .A2(_03570_),
    .A1(net6048));
 sg13g2_a22oi_1 _20160_ (.Y(_03574_),
    .B1(_03571_),
    .B2(net6059),
    .A2(_03569_),
    .A1(net6076));
 sg13g2_a21oi_2 _20161_ (.B1(net6025),
    .Y(_03575_),
    .A2(_03574_),
    .A1(_03573_));
 sg13g2_nor4_2 _20162_ (.A(net6127),
    .B(_03561_),
    .C(_03568_),
    .Y(_03576_),
    .D(_03575_));
 sg13g2_nand2b_1 _20163_ (.Y(_03577_),
    .B(\scanline[124][2] ),
    .A_N(net6224));
 sg13g2_a21oi_1 _20164_ (.A1(net6224),
    .A2(\scanline[125][2] ),
    .Y(_03578_),
    .B1(net6162));
 sg13g2_nand2_1 _20165_ (.Y(_03579_),
    .A(net6217),
    .B(\scanline[127][2] ));
 sg13g2_nand2b_1 _20166_ (.Y(_03580_),
    .B(\scanline[126][2] ),
    .A_N(net6217));
 sg13g2_nand3_1 _20167_ (.B(_03579_),
    .C(_03580_),
    .A(net6162),
    .Y(_03581_));
 sg13g2_a21oi_1 _20168_ (.A1(_03577_),
    .A2(_03578_),
    .Y(_03582_),
    .B1(net6092));
 sg13g2_a21oi_2 _20169_ (.B1(net6116),
    .Y(_03583_),
    .A2(_03582_),
    .A1(_03581_));
 sg13g2_mux4_1 _20170_ (.S0(net6232),
    .A0(\scanline[120][2] ),
    .A1(\scanline[121][2] ),
    .A2(\scanline[122][2] ),
    .A3(\scanline[123][2] ),
    .S1(net6174),
    .X(_03584_));
 sg13g2_and2_1 _20171_ (.A(net6052),
    .B(_03584_),
    .X(_03585_));
 sg13g2_mux4_1 _20172_ (.S0(net6231),
    .A0(\scanline[112][2] ),
    .A1(\scanline[113][2] ),
    .A2(\scanline[114][2] ),
    .A3(\scanline[115][2] ),
    .S1(net6173),
    .X(_03586_));
 sg13g2_mux4_1 _20173_ (.S0(net6231),
    .A0(\scanline[116][2] ),
    .A1(\scanline[117][2] ),
    .A2(\scanline[118][2] ),
    .A3(\scanline[119][2] ),
    .S1(net6173),
    .X(_03587_));
 sg13g2_a221oi_1 _20174_ (.B2(net6064),
    .C1(_03585_),
    .B1(_03587_),
    .A1(net6083),
    .Y(_03588_),
    .A2(_03586_));
 sg13g2_nand2b_1 _20175_ (.Y(_03589_),
    .B(\scanline[100][2] ),
    .A_N(net6229));
 sg13g2_a21oi_1 _20176_ (.A1(net6229),
    .A2(\scanline[101][2] ),
    .Y(_03590_),
    .B1(net6172));
 sg13g2_nand2_1 _20177_ (.Y(_03591_),
    .A(net6229),
    .B(\scanline[103][2] ));
 sg13g2_nand2b_1 _20178_ (.Y(_03592_),
    .B(\scanline[102][2] ),
    .A_N(net6229));
 sg13g2_nand3_1 _20179_ (.B(_03591_),
    .C(_03592_),
    .A(net6172),
    .Y(_03593_));
 sg13g2_a21oi_1 _20180_ (.A1(_03589_),
    .A2(_03590_),
    .Y(_03594_),
    .B1(net6058));
 sg13g2_mux4_1 _20181_ (.S0(net6238),
    .A0(\scanline[96][2] ),
    .A1(\scanline[97][2] ),
    .A2(\scanline[98][2] ),
    .A3(\scanline[99][2] ),
    .S1(net6180),
    .X(_03595_));
 sg13g2_mux4_1 _20182_ (.S0(net6235),
    .A0(\scanline[104][2] ),
    .A1(\scanline[105][2] ),
    .A2(\scanline[106][2] ),
    .A3(\scanline[107][2] ),
    .S1(net6177),
    .X(_03596_));
 sg13g2_mux4_1 _20183_ (.S0(net6240),
    .A0(\scanline[108][2] ),
    .A1(\scanline[109][2] ),
    .A2(\scanline[110][2] ),
    .A3(\scanline[111][2] ),
    .S1(net6181),
    .X(_03597_));
 sg13g2_a22oi_1 _20184_ (.Y(_03598_),
    .B1(_03597_),
    .B2(net6098),
    .A2(_03595_),
    .A1(net6080));
 sg13g2_a221oi_1 _20185_ (.B2(net6052),
    .C1(net6132),
    .B1(_03596_),
    .A1(_03593_),
    .Y(_03599_),
    .A2(_03594_));
 sg13g2_a221oi_1 _20186_ (.B2(_03599_),
    .C1(net6114),
    .B1(_03598_),
    .A1(_03583_),
    .Y(_03600_),
    .A2(_03588_));
 sg13g2_mux4_1 _20187_ (.S0(net6222),
    .A0(\scanline[68][2] ),
    .A1(\scanline[69][2] ),
    .A2(\scanline[70][2] ),
    .A3(\scanline[71][2] ),
    .S1(net6165),
    .X(_03601_));
 sg13g2_mux4_1 _20188_ (.S0(net6225),
    .A0(\scanline[72][2] ),
    .A1(\scanline[73][2] ),
    .A2(\scanline[74][2] ),
    .A3(\scanline[75][2] ),
    .S1(net6167),
    .X(_03602_));
 sg13g2_mux4_1 _20189_ (.S0(net6225),
    .A0(\scanline[64][2] ),
    .A1(\scanline[65][2] ),
    .A2(\scanline[66][2] ),
    .A3(\scanline[67][2] ),
    .S1(net6167),
    .X(_03603_));
 sg13g2_mux4_1 _20190_ (.S0(net6225),
    .A0(\scanline[76][2] ),
    .A1(\scanline[77][2] ),
    .A2(\scanline[78][2] ),
    .A3(\scanline[79][2] ),
    .S1(net6167),
    .X(_03604_));
 sg13g2_a22oi_1 _20191_ (.Y(_03605_),
    .B1(_03604_),
    .B2(net6096),
    .A2(_03602_),
    .A1(net6051));
 sg13g2_a22oi_1 _20192_ (.Y(_03606_),
    .B1(_03603_),
    .B2(net6084),
    .A2(_03601_),
    .A1(net6062));
 sg13g2_a21oi_2 _20193_ (.B1(net6026),
    .Y(_03607_),
    .A2(_03606_),
    .A1(_03605_));
 sg13g2_mux4_1 _20194_ (.S0(net6241),
    .A0(\scanline[92][2] ),
    .A1(\scanline[93][2] ),
    .A2(\scanline[94][2] ),
    .A3(\scanline[95][2] ),
    .S1(net6182),
    .X(_03608_));
 sg13g2_mux4_1 _20195_ (.S0(net6239),
    .A0(\scanline[80][2] ),
    .A1(\scanline[81][2] ),
    .A2(\scanline[82][2] ),
    .A3(\scanline[83][2] ),
    .S1(net6179),
    .X(_03609_));
 sg13g2_a22oi_1 _20196_ (.Y(_03610_),
    .B1(_03609_),
    .B2(net6082),
    .A2(_03608_),
    .A1(net6098));
 sg13g2_mux4_1 _20197_ (.S0(net6242),
    .A0(\scanline[88][2] ),
    .A1(\scanline[89][2] ),
    .A2(\scanline[90][2] ),
    .A3(\scanline[91][2] ),
    .S1(net6183),
    .X(_03611_));
 sg13g2_mux4_1 _20198_ (.S0(net6241),
    .A0(\scanline[84][2] ),
    .A1(\scanline[85][2] ),
    .A2(\scanline[86][2] ),
    .A3(\scanline[87][2] ),
    .S1(net6182),
    .X(_03612_));
 sg13g2_a22oi_1 _20199_ (.Y(_03613_),
    .B1(_03612_),
    .B2(net6065),
    .A2(_03611_),
    .A1(net6053));
 sg13g2_a21oi_1 _20200_ (.A1(_03610_),
    .A2(_03613_),
    .Y(_03614_),
    .B1(net6012));
 sg13g2_or3_1 _20201_ (.A(_08656_),
    .B(_03607_),
    .C(_03614_),
    .X(_03615_));
 sg13g2_o21ai_1 _20202_ (.B1(_08655_),
    .Y(_03616_),
    .A1(_03600_),
    .A2(_03615_));
 sg13g2_o21ai_1 _20203_ (.B1(_03543_),
    .Y(_03617_),
    .A1(_03576_),
    .A2(_03616_));
 sg13g2_inv_2 _20204_ (.Y(_03618_),
    .A(net5920));
 sg13g2_mux4_1 _20205_ (.S0(net6206),
    .A0(\scanline[152][0] ),
    .A1(\scanline[153][0] ),
    .A2(\scanline[154][0] ),
    .A3(\scanline[155][0] ),
    .S1(net6151),
    .X(_03619_));
 sg13g2_nor2_1 _20206_ (.A(net6045),
    .B(_03619_),
    .Y(_03620_));
 sg13g2_mux4_1 _20207_ (.S0(net6205),
    .A0(\scanline[144][0] ),
    .A1(\scanline[145][0] ),
    .A2(\scanline[146][0] ),
    .A3(\scanline[147][0] ),
    .S1(net6150),
    .X(_03621_));
 sg13g2_nor2_1 _20208_ (.A(net6073),
    .B(_03621_),
    .Y(_03622_));
 sg13g2_mux4_1 _20209_ (.S0(net6206),
    .A0(\scanline[148][0] ),
    .A1(\scanline[149][0] ),
    .A2(\scanline[150][0] ),
    .A3(\scanline[151][0] ),
    .S1(net6151),
    .X(_03623_));
 sg13g2_nor2_1 _20210_ (.A(net6057),
    .B(_03623_),
    .Y(_03624_));
 sg13g2_nor3_1 _20211_ (.A(_03620_),
    .B(_03622_),
    .C(_03624_),
    .Y(_03625_));
 sg13g2_mux4_1 _20212_ (.S0(net6204),
    .A0(\scanline[156][0] ),
    .A1(\scanline[157][0] ),
    .A2(\scanline[158][0] ),
    .A3(\scanline[159][0] ),
    .S1(net6149),
    .X(_03626_));
 sg13g2_mux4_1 _20213_ (.S0(net6191),
    .A0(\scanline[140][0] ),
    .A1(\scanline[141][0] ),
    .A2(\scanline[142][0] ),
    .A3(\scanline[143][0] ),
    .S1(net6139),
    .X(_03627_));
 sg13g2_nor2_1 _20214_ (.A(net6091),
    .B(_03627_),
    .Y(_03628_));
 sg13g2_mux4_1 _20215_ (.S0(net6190),
    .A0(\scanline[136][0] ),
    .A1(\scanline[137][0] ),
    .A2(\scanline[138][0] ),
    .A3(\scanline[139][0] ),
    .S1(net6138),
    .X(_03629_));
 sg13g2_nor2_1 _20216_ (.A(net6044),
    .B(_03629_),
    .Y(_03630_));
 sg13g2_mux4_1 _20217_ (.S0(net6190),
    .A0(\scanline[132][0] ),
    .A1(\scanline[133][0] ),
    .A2(\scanline[134][0] ),
    .A3(\scanline[135][0] ),
    .S1(net6138),
    .X(_03631_));
 sg13g2_nor2_1 _20218_ (.A(net6056),
    .B(_03631_),
    .Y(_03632_));
 sg13g2_o21ai_1 _20219_ (.B1(_03625_),
    .Y(_03633_),
    .A1(net6091),
    .A2(_03626_));
 sg13g2_mux4_1 _20220_ (.S0(net6192),
    .A0(\scanline[128][0] ),
    .A1(\scanline[129][0] ),
    .A2(\scanline[130][0] ),
    .A3(\scanline[131][0] ),
    .S1(net6140),
    .X(_03634_));
 sg13g2_nor2_1 _20221_ (.A(net6074),
    .B(_03634_),
    .Y(_03635_));
 sg13g2_nor4_2 _20222_ (.A(_03628_),
    .B(_03630_),
    .C(_03632_),
    .Y(_03636_),
    .D(_03635_));
 sg13g2_nor2_1 _20223_ (.A(net6129),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_o21ai_1 _20224_ (.B1(_09219_),
    .Y(_03638_),
    .A1(net6129),
    .A2(_03636_));
 sg13g2_a21oi_1 _20225_ (.A1(net6129),
    .A2(_03633_),
    .Y(_03639_),
    .B1(_03637_));
 sg13g2_a21oi_1 _20226_ (.A1(net6129),
    .A2(_03633_),
    .Y(_03640_),
    .B1(_03638_));
 sg13g2_mux4_1 _20227_ (.S0(net6215),
    .A0(\scanline[44][0] ),
    .A1(\scanline[45][0] ),
    .A2(\scanline[46][0] ),
    .A3(\scanline[47][0] ),
    .S1(net6160),
    .X(_03641_));
 sg13g2_mux4_1 _20228_ (.S0(net6195),
    .A0(\scanline[40][0] ),
    .A1(\scanline[41][0] ),
    .A2(\scanline[42][0] ),
    .A3(\scanline[43][0] ),
    .S1(net6142),
    .X(_03642_));
 sg13g2_mux4_1 _20229_ (.S0(net6195),
    .A0(\scanline[36][0] ),
    .A1(\scanline[37][0] ),
    .A2(\scanline[38][0] ),
    .A3(\scanline[39][0] ),
    .S1(net6142),
    .X(_03643_));
 sg13g2_nand2b_1 _20230_ (.Y(_03644_),
    .B(\scanline[32][0] ),
    .A_N(net6216));
 sg13g2_a21oi_1 _20231_ (.A1(net6216),
    .A2(\scanline[33][0] ),
    .Y(_03645_),
    .B1(net6161));
 sg13g2_nand2_1 _20232_ (.Y(_03646_),
    .A(net6219),
    .B(\scanline[35][0] ));
 sg13g2_nand2b_1 _20233_ (.Y(_03647_),
    .B(\scanline[34][0] ),
    .A_N(net6219));
 sg13g2_nand3_1 _20234_ (.B(_03646_),
    .C(_03647_),
    .A(net6161),
    .Y(_03648_));
 sg13g2_a21oi_1 _20235_ (.A1(_03644_),
    .A2(_03645_),
    .Y(_03649_),
    .B1(net6075));
 sg13g2_a22oi_1 _20236_ (.Y(_03650_),
    .B1(_03643_),
    .B2(net6060),
    .A2(_03642_),
    .A1(net6047));
 sg13g2_a221oi_1 _20237_ (.B2(_03649_),
    .C1(net6131),
    .B1(_03648_),
    .A1(net6093),
    .Y(_03651_),
    .A2(_03641_));
 sg13g2_mux4_1 _20238_ (.S0(net6198),
    .A0(\scanline[48][0] ),
    .A1(\scanline[49][0] ),
    .A2(\scanline[50][0] ),
    .A3(\scanline[51][0] ),
    .S1(net6144),
    .X(_03652_));
 sg13g2_and2_1 _20239_ (.A(net6077),
    .B(_03652_),
    .X(_03653_));
 sg13g2_mux4_1 _20240_ (.S0(net6201),
    .A0(\scanline[56][0] ),
    .A1(\scanline[57][0] ),
    .A2(\scanline[58][0] ),
    .A3(\scanline[59][0] ),
    .S1(net6145),
    .X(_03654_));
 sg13g2_mux4_1 _20241_ (.S0(net6201),
    .A0(\scanline[52][0] ),
    .A1(\scanline[53][0] ),
    .A2(\scanline[54][0] ),
    .A3(\scanline[55][0] ),
    .S1(net6146),
    .X(_03655_));
 sg13g2_mux4_1 _20242_ (.S0(net6195),
    .A0(\scanline[60][0] ),
    .A1(\scanline[61][0] ),
    .A2(\scanline[62][0] ),
    .A3(\scanline[63][0] ),
    .S1(net6142),
    .X(_03656_));
 sg13g2_a21oi_1 _20243_ (.A1(net6047),
    .A2(_03654_),
    .Y(_03657_),
    .B1(net6115));
 sg13g2_a221oi_1 _20244_ (.B2(net6101),
    .C1(_03653_),
    .B1(_03656_),
    .A1(net6060),
    .Y(_03658_),
    .A2(_03655_));
 sg13g2_a221oi_1 _20245_ (.B2(_03658_),
    .C1(net6113),
    .B1(_03657_),
    .A1(_03650_),
    .Y(_03659_),
    .A2(_03651_));
 sg13g2_mux4_1 _20246_ (.S0(net6221),
    .A0(\scanline[20][0] ),
    .A1(\scanline[21][0] ),
    .A2(\scanline[22][0] ),
    .A3(\scanline[23][0] ),
    .S1(net6164),
    .X(_03660_));
 sg13g2_mux4_1 _20247_ (.S0(net6213),
    .A0(\scanline[16][0] ),
    .A1(\scanline[17][0] ),
    .A2(\scanline[18][0] ),
    .A3(\scanline[19][0] ),
    .S1(net6158),
    .X(_03661_));
 sg13g2_mux4_1 _20248_ (.S0(net6213),
    .A0(\scanline[28][0] ),
    .A1(\scanline[29][0] ),
    .A2(\scanline[30][0] ),
    .A3(\scanline[31][0] ),
    .S1(net6158),
    .X(_03662_));
 sg13g2_mux4_1 _20249_ (.S0(net6223),
    .A0(\scanline[24][0] ),
    .A1(\scanline[25][0] ),
    .A2(\scanline[26][0] ),
    .A3(\scanline[27][0] ),
    .S1(net6166),
    .X(_03663_));
 sg13g2_a22oi_1 _20250_ (.Y(_03664_),
    .B1(_03663_),
    .B2(net6051),
    .A2(_03661_),
    .A1(net6079));
 sg13g2_a22oi_1 _20251_ (.Y(_03665_),
    .B1(_03662_),
    .B2(net6096),
    .A2(_03660_),
    .A1(net6063));
 sg13g2_a21oi_2 _20252_ (.B1(net6011),
    .Y(_03666_),
    .A2(_03665_),
    .A1(_03664_));
 sg13g2_mux4_1 _20253_ (.S0(net6186),
    .A0(\scanline[4][0] ),
    .A1(\scanline[5][0] ),
    .A2(\scanline[6][0] ),
    .A3(\scanline[7][0] ),
    .S1(net6135),
    .X(_03667_));
 sg13g2_mux4_1 _20254_ (.S0(net6194),
    .A0(\scanline[0][0] ),
    .A1(\scanline[1][0] ),
    .A2(\scanline[2][0] ),
    .A3(\scanline[3][0] ),
    .S1(net6143),
    .X(_03668_));
 sg13g2_mux4_1 _20255_ (.S0(net6186),
    .A0(\scanline[12][0] ),
    .A1(\scanline[13][0] ),
    .A2(\scanline[14][0] ),
    .A3(\scanline[15][0] ),
    .S1(net6135),
    .X(_03669_));
 sg13g2_mux4_1 _20256_ (.S0(net6194),
    .A0(\scanline[8][0] ),
    .A1(\scanline[9][0] ),
    .A2(\scanline[10][0] ),
    .A3(\scanline[11][0] ),
    .S1(net6141),
    .X(_03670_));
 sg13g2_a22oi_1 _20257_ (.Y(_03671_),
    .B1(_03670_),
    .B2(net6048),
    .A2(_03668_),
    .A1(net6076));
 sg13g2_a22oi_1 _20258_ (.Y(_03672_),
    .B1(_03669_),
    .B2(net6094),
    .A2(_03667_),
    .A1(net6059));
 sg13g2_a21oi_1 _20259_ (.A1(_03671_),
    .A2(_03672_),
    .Y(_03673_),
    .B1(net6025));
 sg13g2_or4_2 _20260_ (.A(net6127),
    .B(_03659_),
    .C(_03666_),
    .D(_03673_),
    .X(_03674_));
 sg13g2_nand2b_1 _20261_ (.Y(_03675_),
    .B(\scanline[120][0] ),
    .A_N(net6231));
 sg13g2_a21oi_1 _20262_ (.A1(net6232),
    .A2(\scanline[121][0] ),
    .Y(_03676_),
    .B1(net6174));
 sg13g2_nand2_1 _20263_ (.Y(_03677_),
    .A(net6232),
    .B(\scanline[123][0] ));
 sg13g2_nand2b_1 _20264_ (.Y(_03678_),
    .B(\scanline[122][0] ),
    .A_N(net6232));
 sg13g2_nand3_1 _20265_ (.B(_03677_),
    .C(_03678_),
    .A(net6174),
    .Y(_03679_));
 sg13g2_a21oi_1 _20266_ (.A1(_03675_),
    .A2(_03676_),
    .Y(_03680_),
    .B1(net6046));
 sg13g2_mux4_1 _20267_ (.S0(net6231),
    .A0(\scanline[112][0] ),
    .A1(\scanline[113][0] ),
    .A2(\scanline[114][0] ),
    .A3(\scanline[115][0] ),
    .S1(net6173),
    .X(_03681_));
 sg13g2_mux4_1 _20268_ (.S0(net6219),
    .A0(\scanline[124][0] ),
    .A1(\scanline[125][0] ),
    .A2(\scanline[126][0] ),
    .A3(\scanline[127][0] ),
    .S1(net6162),
    .X(_03682_));
 sg13g2_and2_2 _20269_ (.A(net6099),
    .B(_03682_),
    .X(_03683_));
 sg13g2_mux4_1 _20270_ (.S0(net6232),
    .A0(\scanline[116][0] ),
    .A1(\scanline[117][0] ),
    .A2(\scanline[118][0] ),
    .A3(\scanline[119][0] ),
    .S1(net6174),
    .X(_03684_));
 sg13g2_a21oi_1 _20271_ (.A1(net6078),
    .A2(_03681_),
    .Y(_03685_),
    .B1(net6116));
 sg13g2_a221oi_1 _20272_ (.B2(net6064),
    .C1(_03683_),
    .B1(_03684_),
    .A1(_03679_),
    .Y(_03686_),
    .A2(_03680_));
 sg13g2_mux4_1 _20273_ (.S0(net6234),
    .A0(\scanline[108][0] ),
    .A1(\scanline[109][0] ),
    .A2(\scanline[110][0] ),
    .A3(\scanline[111][0] ),
    .S1(net6176),
    .X(_03687_));
 sg13g2_mux4_1 _20274_ (.S0(net6238),
    .A0(\scanline[96][0] ),
    .A1(\scanline[97][0] ),
    .A2(\scanline[98][0] ),
    .A3(\scanline[99][0] ),
    .S1(net6178),
    .X(_03688_));
 sg13g2_mux4_1 _20275_ (.S0(net6235),
    .A0(\scanline[104][0] ),
    .A1(\scanline[105][0] ),
    .A2(\scanline[106][0] ),
    .A3(\scanline[107][0] ),
    .S1(net6176),
    .X(_03689_));
 sg13g2_mux4_1 _20276_ (.S0(net6237),
    .A0(\scanline[100][0] ),
    .A1(\scanline[101][0] ),
    .A2(\scanline[102][0] ),
    .A3(\scanline[103][0] ),
    .S1(net6178),
    .X(_03690_));
 sg13g2_a22oi_1 _20277_ (.Y(_03691_),
    .B1(_03690_),
    .B2(net6066),
    .A2(_03688_),
    .A1(net6080));
 sg13g2_a221oi_1 _20278_ (.B2(net6053),
    .C1(net6132),
    .B1(_03689_),
    .A1(net6099),
    .Y(_03692_),
    .A2(_03687_));
 sg13g2_a21o_1 _20279_ (.A2(_03692_),
    .A1(_03691_),
    .B1(net6114),
    .X(_03693_));
 sg13g2_a21o_1 _20280_ (.A2(_03686_),
    .A1(_03685_),
    .B1(_03693_),
    .X(_03694_));
 sg13g2_mux4_1 _20281_ (.S0(net6241),
    .A0(\scanline[92][0] ),
    .A1(\scanline[93][0] ),
    .A2(\scanline[94][0] ),
    .A3(\scanline[95][0] ),
    .S1(net6182),
    .X(_03695_));
 sg13g2_mux4_1 _20282_ (.S0(net6242),
    .A0(\scanline[88][0] ),
    .A1(\scanline[89][0] ),
    .A2(\scanline[90][0] ),
    .A3(\scanline[91][0] ),
    .S1(net6183),
    .X(_03696_));
 sg13g2_a22oi_1 _20283_ (.Y(_03697_),
    .B1(_03696_),
    .B2(net6053),
    .A2(_03695_),
    .A1(net6097));
 sg13g2_mux4_1 _20284_ (.S0(net6241),
    .A0(\scanline[84][0] ),
    .A1(\scanline[85][0] ),
    .A2(\scanline[86][0] ),
    .A3(\scanline[87][0] ),
    .S1(net6182),
    .X(_03698_));
 sg13g2_mux4_1 _20285_ (.S0(net6239),
    .A0(\scanline[80][0] ),
    .A1(\scanline[81][0] ),
    .A2(\scanline[82][0] ),
    .A3(\scanline[83][0] ),
    .S1(net6179),
    .X(_03699_));
 sg13g2_a22oi_1 _20286_ (.Y(_03700_),
    .B1(_03699_),
    .B2(net6082),
    .A2(_03698_),
    .A1(net6065));
 sg13g2_a21oi_1 _20287_ (.A1(_03697_),
    .A2(_03700_),
    .Y(_03701_),
    .B1(net6012));
 sg13g2_mux4_1 _20288_ (.S0(net6225),
    .A0(\scanline[76][0] ),
    .A1(\scanline[77][0] ),
    .A2(\scanline[78][0] ),
    .A3(\scanline[79][0] ),
    .S1(net6167),
    .X(_03702_));
 sg13g2_mux4_1 _20289_ (.S0(net6225),
    .A0(\scanline[72][0] ),
    .A1(\scanline[73][0] ),
    .A2(\scanline[74][0] ),
    .A3(\scanline[75][0] ),
    .S1(net6167),
    .X(_03703_));
 sg13g2_mux4_1 _20290_ (.S0(net6222),
    .A0(\scanline[68][0] ),
    .A1(\scanline[69][0] ),
    .A2(\scanline[70][0] ),
    .A3(\scanline[71][0] ),
    .S1(net6165),
    .X(_03704_));
 sg13g2_mux4_1 _20291_ (.S0(net6225),
    .A0(\scanline[64][0] ),
    .A1(\scanline[65][0] ),
    .A2(\scanline[66][0] ),
    .A3(\scanline[67][0] ),
    .S1(net6167),
    .X(_03705_));
 sg13g2_a22oi_1 _20292_ (.Y(_03706_),
    .B1(_03705_),
    .B2(net6084),
    .A2(_03703_),
    .A1(net6051));
 sg13g2_a22oi_1 _20293_ (.Y(_03707_),
    .B1(_03704_),
    .B2(net6066),
    .A2(_03702_),
    .A1(net6096));
 sg13g2_a21oi_2 _20294_ (.B1(net6026),
    .Y(_03708_),
    .A2(_03707_),
    .A1(_03706_));
 sg13g2_nor3_2 _20295_ (.A(_08656_),
    .B(_03701_),
    .C(_03708_),
    .Y(_03709_));
 sg13g2_a21oi_2 _20296_ (.B1(net6125),
    .Y(_03710_),
    .A2(_03709_),
    .A1(_03694_));
 sg13g2_a22oi_1 _20297_ (.Y(_03711_),
    .B1(_03674_),
    .B2(_03710_),
    .A2(_03639_),
    .A1(_09219_));
 sg13g2_a21o_1 _20298_ (.A2(_03710_),
    .A1(_03674_),
    .B1(_03640_),
    .X(_03712_));
 sg13g2_nand2_2 _20299_ (.Y(_03713_),
    .A(net6085),
    .B(net5919));
 sg13g2_and2_1 _20300_ (.A(net6085),
    .B(net5923),
    .X(_03714_));
 sg13g2_nand2_1 _20301_ (.Y(_03715_),
    .A(net6085),
    .B(net5920));
 sg13g2_and3_2 _20302_ (.X(_03716_),
    .A(net6087),
    .B(net5921),
    .C(net5919));
 sg13g2_nand2_2 _20303_ (.Y(_03717_),
    .A(net6086),
    .B(net5926));
 sg13g2_and3_2 _20304_ (.X(_03718_),
    .A(net6086),
    .B(net5925),
    .C(net5922));
 sg13g2_nand3_1 _20305_ (.B(net5924),
    .C(net5921),
    .A(net6085),
    .Y(_03719_));
 sg13g2_and4_2 _20306_ (.A(net6086),
    .B(net5925),
    .C(net5922),
    .D(_03712_),
    .X(_03720_));
 sg13g2_nand3b_1 _20307_ (.B(net5924),
    .C(net6085),
    .Y(_03721_),
    .A_N(net5920));
 sg13g2_inv_1 _20308_ (.Y(_03722_),
    .A(net5893));
 sg13g2_and3_2 _20309_ (.X(_03723_),
    .A(net6086),
    .B(net5926),
    .C(_03711_));
 sg13g2_nor2_2 _20310_ (.A(net5919),
    .B(net5893),
    .Y(_03724_));
 sg13g2_a21oi_2 _20311_ (.B1(_03720_),
    .Y(_03725_),
    .A2(_03723_),
    .A1(_03618_));
 sg13g2_mux4_1 _20312_ (.S0(net6204),
    .A0(\scanline[152][4] ),
    .A1(\scanline[153][4] ),
    .A2(\scanline[154][4] ),
    .A3(\scanline[155][4] ),
    .S1(net6150),
    .X(_03726_));
 sg13g2_nor2_1 _20313_ (.A(net6045),
    .B(_03726_),
    .Y(_03727_));
 sg13g2_mux4_1 _20314_ (.S0(net6204),
    .A0(\scanline[156][4] ),
    .A1(\scanline[157][4] ),
    .A2(\scanline[158][4] ),
    .A3(\scanline[159][4] ),
    .S1(net6149),
    .X(_03728_));
 sg13g2_nor2_1 _20315_ (.A(net6090),
    .B(_03728_),
    .Y(_03729_));
 sg13g2_mux4_1 _20316_ (.S0(net6204),
    .A0(\scanline[144][4] ),
    .A1(\scanline[145][4] ),
    .A2(\scanline[146][4] ),
    .A3(\scanline[147][4] ),
    .S1(net6149),
    .X(_03730_));
 sg13g2_nor2_1 _20317_ (.A(net6073),
    .B(_03730_),
    .Y(_03731_));
 sg13g2_mux4_1 _20318_ (.S0(net6207),
    .A0(\scanline[148][4] ),
    .A1(\scanline[149][4] ),
    .A2(\scanline[150][4] ),
    .A3(\scanline[151][4] ),
    .S1(net6152),
    .X(_03732_));
 sg13g2_o21ai_1 _20319_ (.B1(net6128),
    .Y(_03733_),
    .A1(net6057),
    .A2(_03732_));
 sg13g2_nor4_1 _20320_ (.A(_03727_),
    .B(_03729_),
    .C(_03731_),
    .D(_03733_),
    .Y(_03734_));
 sg13g2_mux4_1 _20321_ (.S0(net6203),
    .A0(\scanline[140][4] ),
    .A1(\scanline[141][4] ),
    .A2(\scanline[142][4] ),
    .A3(\scanline[143][4] ),
    .S1(net6148),
    .X(_03735_));
 sg13g2_o21ai_1 _20322_ (.B1(net6117),
    .Y(_03736_),
    .A1(net6090),
    .A2(_03735_));
 sg13g2_mux4_1 _20323_ (.S0(net6190),
    .A0(\scanline[136][4] ),
    .A1(\scanline[137][4] ),
    .A2(\scanline[138][4] ),
    .A3(\scanline[139][4] ),
    .S1(net6138),
    .X(_03737_));
 sg13g2_nor2_1 _20324_ (.A(net6044),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_mux4_1 _20325_ (.S0(net6190),
    .A0(\scanline[132][4] ),
    .A1(\scanline[133][4] ),
    .A2(\scanline[134][4] ),
    .A3(\scanline[135][4] ),
    .S1(net6138),
    .X(_03739_));
 sg13g2_nor2_1 _20326_ (.A(net6056),
    .B(_03739_),
    .Y(_03740_));
 sg13g2_mux4_1 _20327_ (.S0(net6192),
    .A0(\scanline[128][4] ),
    .A1(\scanline[129][4] ),
    .A2(\scanline[130][4] ),
    .A3(\scanline[131][4] ),
    .S1(net6140),
    .X(_03741_));
 sg13g2_nor2_1 _20328_ (.A(net6074),
    .B(_03741_),
    .Y(_03742_));
 sg13g2_nor4_2 _20329_ (.A(_03736_),
    .B(_03738_),
    .C(_03740_),
    .Y(_03743_),
    .D(_03742_));
 sg13g2_o21ai_1 _20330_ (.B1(_09219_),
    .Y(_03744_),
    .A1(_03734_),
    .A2(_03743_));
 sg13g2_mux4_1 _20331_ (.S0(net6215),
    .A0(\scanline[44][4] ),
    .A1(\scanline[45][4] ),
    .A2(\scanline[46][4] ),
    .A3(\scanline[47][4] ),
    .S1(net6160),
    .X(_03745_));
 sg13g2_mux4_1 _20332_ (.S0(net6195),
    .A0(\scanline[40][4] ),
    .A1(\scanline[41][4] ),
    .A2(\scanline[42][4] ),
    .A3(\scanline[43][4] ),
    .S1(net6142),
    .X(_03746_));
 sg13g2_mux4_1 _20333_ (.S0(net6215),
    .A0(\scanline[32][4] ),
    .A1(\scanline[33][4] ),
    .A2(\scanline[34][4] ),
    .A3(\scanline[35][4] ),
    .S1(net6160),
    .X(_03747_));
 sg13g2_mux4_1 _20334_ (.S0(net6195),
    .A0(\scanline[36][4] ),
    .A1(\scanline[37][4] ),
    .A2(\scanline[38][4] ),
    .A3(\scanline[39][4] ),
    .S1(net6142),
    .X(_03748_));
 sg13g2_a22oi_1 _20335_ (.Y(_03749_),
    .B1(_03748_),
    .B2(net6060),
    .A2(_03746_),
    .A1(net6047));
 sg13g2_a221oi_1 _20336_ (.B2(net6077),
    .C1(net6131),
    .B1(_03747_),
    .A1(net6095),
    .Y(_03750_),
    .A2(_03745_));
 sg13g2_mux4_1 _20337_ (.S0(net6196),
    .A0(\scanline[60][4] ),
    .A1(\scanline[61][4] ),
    .A2(\scanline[62][4] ),
    .A3(\scanline[63][4] ),
    .S1(net6143),
    .X(_03751_));
 sg13g2_mux4_1 _20338_ (.S0(net6208),
    .A0(\scanline[56][4] ),
    .A1(\scanline[57][4] ),
    .A2(\scanline[58][4] ),
    .A3(\scanline[59][4] ),
    .S1(net6153),
    .X(_03752_));
 sg13g2_and2_1 _20339_ (.A(net6049),
    .B(_03752_),
    .X(_03753_));
 sg13g2_mux4_1 _20340_ (.S0(net6208),
    .A0(\scanline[52][4] ),
    .A1(\scanline[53][4] ),
    .A2(\scanline[54][4] ),
    .A3(\scanline[55][4] ),
    .S1(net6154),
    .X(_03754_));
 sg13g2_mux4_1 _20341_ (.S0(net6198),
    .A0(\scanline[48][4] ),
    .A1(\scanline[49][4] ),
    .A2(\scanline[50][4] ),
    .A3(\scanline[51][4] ),
    .S1(net6144),
    .X(_03755_));
 sg13g2_a21oi_2 _20342_ (.B1(_03753_),
    .Y(_03756_),
    .A2(_03754_),
    .A1(net6061));
 sg13g2_a221oi_1 _20343_ (.B2(net6077),
    .C1(net6117),
    .B1(_03755_),
    .A1(net6093),
    .Y(_03757_),
    .A2(_03751_));
 sg13g2_a221oi_1 _20344_ (.B2(_03757_),
    .C1(net6113),
    .B1(_03756_),
    .A1(_03749_),
    .Y(_03758_),
    .A2(_03750_));
 sg13g2_mux4_1 _20345_ (.S0(net6221),
    .A0(\scanline[20][4] ),
    .A1(\scanline[21][4] ),
    .A2(\scanline[22][4] ),
    .A3(\scanline[23][4] ),
    .S1(net6164),
    .X(_03759_));
 sg13g2_mux4_1 _20346_ (.S0(net6212),
    .A0(\scanline[16][4] ),
    .A1(\scanline[17][4] ),
    .A2(\scanline[18][4] ),
    .A3(\scanline[19][4] ),
    .S1(net6157),
    .X(_03760_));
 sg13g2_a22oi_1 _20347_ (.Y(_03761_),
    .B1(_03760_),
    .B2(net6079),
    .A2(_03759_),
    .A1(net6063));
 sg13g2_mux4_1 _20348_ (.S0(net6220),
    .A0(\scanline[28][4] ),
    .A1(\scanline[29][4] ),
    .A2(\scanline[30][4] ),
    .A3(\scanline[31][4] ),
    .S1(net6162),
    .X(_03762_));
 sg13g2_mux4_1 _20349_ (.S0(net6224),
    .A0(\scanline[24][4] ),
    .A1(\scanline[25][4] ),
    .A2(\scanline[26][4] ),
    .A3(\scanline[27][4] ),
    .S1(net6169),
    .X(_03763_));
 sg13g2_a22oi_1 _20350_ (.Y(_03764_),
    .B1(_03763_),
    .B2(net6051),
    .A2(_03762_),
    .A1(net6096));
 sg13g2_a21oi_2 _20351_ (.B1(net6011),
    .Y(_03765_),
    .A2(_03764_),
    .A1(_03761_));
 sg13g2_mux4_1 _20352_ (.S0(net6186),
    .A0(\scanline[12][4] ),
    .A1(\scanline[13][4] ),
    .A2(\scanline[14][4] ),
    .A3(\scanline[15][4] ),
    .S1(net6135),
    .X(_03766_));
 sg13g2_mux4_1 _20353_ (.S0(net6188),
    .A0(\scanline[4][4] ),
    .A1(\scanline[5][4] ),
    .A2(\scanline[6][4] ),
    .A3(\scanline[7][4] ),
    .S1(net6137),
    .X(_03767_));
 sg13g2_mux4_1 _20354_ (.S0(net6193),
    .A0(\scanline[0][4] ),
    .A1(\scanline[1][4] ),
    .A2(\scanline[2][4] ),
    .A3(\scanline[3][4] ),
    .S1(net6141),
    .X(_03768_));
 sg13g2_mux4_1 _20355_ (.S0(net6188),
    .A0(\scanline[8][4] ),
    .A1(\scanline[9][4] ),
    .A2(\scanline[10][4] ),
    .A3(\scanline[11][4] ),
    .S1(net6137),
    .X(_03769_));
 sg13g2_a22oi_1 _20356_ (.Y(_03770_),
    .B1(_03769_),
    .B2(net6048),
    .A2(_03767_),
    .A1(net6059));
 sg13g2_a22oi_1 _20357_ (.Y(_03771_),
    .B1(_03768_),
    .B2(net6076),
    .A2(_03766_),
    .A1(net6094));
 sg13g2_a21oi_2 _20358_ (.B1(net6025),
    .Y(_03772_),
    .A2(_03771_),
    .A1(_03770_));
 sg13g2_nor4_2 _20359_ (.A(net6127),
    .B(_03758_),
    .C(_03765_),
    .Y(_03773_),
    .D(_03772_));
 sg13g2_nand2b_1 _20360_ (.Y(_03774_),
    .B(\scanline[104][4] ),
    .A_N(net6235));
 sg13g2_a21oi_1 _20361_ (.A1(net6235),
    .A2(\scanline[105][4] ),
    .Y(_03775_),
    .B1(net6174));
 sg13g2_nand2_1 _20362_ (.Y(_03776_),
    .A(net6234),
    .B(\scanline[107][4] ));
 sg13g2_nand2b_1 _20363_ (.Y(_03777_),
    .B(\scanline[106][4] ),
    .A_N(net6234));
 sg13g2_nand3_1 _20364_ (.B(_03776_),
    .C(_03777_),
    .A(net6176),
    .Y(_03778_));
 sg13g2_a21oi_1 _20365_ (.A1(_03774_),
    .A2(_03775_),
    .Y(_03779_),
    .B1(net6046));
 sg13g2_a21oi_2 _20366_ (.B1(net6132),
    .Y(_03780_),
    .A2(_03779_),
    .A1(_03778_));
 sg13g2_mux4_1 _20367_ (.S0(net6243),
    .A0(\scanline[96][4] ),
    .A1(\scanline[97][4] ),
    .A2(\scanline[98][4] ),
    .A3(\scanline[99][4] ),
    .S1(net6180),
    .X(_03781_));
 sg13g2_mux4_1 _20368_ (.S0(net6240),
    .A0(\scanline[108][4] ),
    .A1(\scanline[109][4] ),
    .A2(\scanline[110][4] ),
    .A3(\scanline[111][4] ),
    .S1(net6181),
    .X(_03782_));
 sg13g2_and2_1 _20369_ (.A(net6098),
    .B(_03782_),
    .X(_03783_));
 sg13g2_mux4_1 _20370_ (.S0(net6238),
    .A0(\scanline[100][4] ),
    .A1(\scanline[101][4] ),
    .A2(\scanline[102][4] ),
    .A3(\scanline[103][4] ),
    .S1(net6180),
    .X(_03784_));
 sg13g2_a221oi_1 _20371_ (.B2(net6066),
    .C1(_03783_),
    .B1(_03784_),
    .A1(net6080),
    .Y(_03785_),
    .A2(_03781_));
 sg13g2_nand2b_1 _20372_ (.Y(_03786_),
    .B(\scanline[124][4] ),
    .A_N(net6218));
 sg13g2_a21oi_1 _20373_ (.A1(net6218),
    .A2(\scanline[125][4] ),
    .Y(_03787_),
    .B1(net6162));
 sg13g2_nand2_1 _20374_ (.Y(_03788_),
    .A(net6218),
    .B(\scanline[127][4] ));
 sg13g2_nand2b_1 _20375_ (.Y(_03789_),
    .B(\scanline[126][4] ),
    .A_N(net6219));
 sg13g2_nand3_1 _20376_ (.B(_03788_),
    .C(_03789_),
    .A(net6162),
    .Y(_03790_));
 sg13g2_a21oi_1 _20377_ (.A1(_03786_),
    .A2(_03787_),
    .Y(_03791_),
    .B1(net6092));
 sg13g2_mux4_1 _20378_ (.S0(net6232),
    .A0(\scanline[116][4] ),
    .A1(\scanline[117][4] ),
    .A2(\scanline[118][4] ),
    .A3(\scanline[119][4] ),
    .S1(net6174),
    .X(_03792_));
 sg13g2_mux4_1 _20379_ (.S0(net6232),
    .A0(\scanline[120][4] ),
    .A1(\scanline[121][4] ),
    .A2(\scanline[122][4] ),
    .A3(\scanline[123][4] ),
    .S1(net6175),
    .X(_03793_));
 sg13g2_mux4_1 _20380_ (.S0(net6230),
    .A0(\scanline[112][4] ),
    .A1(\scanline[113][4] ),
    .A2(\scanline[114][4] ),
    .A3(\scanline[115][4] ),
    .S1(net6171),
    .X(_03794_));
 sg13g2_a22oi_1 _20381_ (.Y(_03795_),
    .B1(_03793_),
    .B2(net6052),
    .A2(_03792_),
    .A1(net6064));
 sg13g2_a221oi_1 _20382_ (.B2(net6080),
    .C1(net6115),
    .B1(_03794_),
    .A1(_03790_),
    .Y(_03796_),
    .A2(_03791_));
 sg13g2_a221oi_1 _20383_ (.B2(_03796_),
    .C1(net6114),
    .B1(_03795_),
    .A1(_03780_),
    .Y(_03797_),
    .A2(_03785_));
 sg13g2_mux4_1 _20384_ (.S0(net6222),
    .A0(\scanline[68][4] ),
    .A1(\scanline[69][4] ),
    .A2(\scanline[70][4] ),
    .A3(\scanline[71][4] ),
    .S1(net6165),
    .X(_03798_));
 sg13g2_mux4_1 _20385_ (.S0(net6223),
    .A0(\scanline[72][4] ),
    .A1(\scanline[73][4] ),
    .A2(\scanline[74][4] ),
    .A3(\scanline[75][4] ),
    .S1(net6166),
    .X(_03799_));
 sg13g2_a22oi_1 _20386_ (.Y(_03800_),
    .B1(_03799_),
    .B2(net6050),
    .A2(_03798_),
    .A1(net6062));
 sg13g2_mux4_1 _20387_ (.S0(net6226),
    .A0(\scanline[64][4] ),
    .A1(\scanline[65][4] ),
    .A2(\scanline[66][4] ),
    .A3(\scanline[67][4] ),
    .S1(net6168),
    .X(_03801_));
 sg13g2_mux4_1 _20388_ (.S0(net6226),
    .A0(\scanline[76][4] ),
    .A1(\scanline[77][4] ),
    .A2(\scanline[78][4] ),
    .A3(\scanline[79][4] ),
    .S1(net6168),
    .X(_03802_));
 sg13g2_a22oi_1 _20389_ (.Y(_03803_),
    .B1(_03802_),
    .B2(net6095),
    .A2(_03801_),
    .A1(net6081));
 sg13g2_a21oi_1 _20390_ (.A1(_03800_),
    .A2(_03803_),
    .Y(_03804_),
    .B1(net6026));
 sg13g2_mux4_1 _20391_ (.S0(net6241),
    .A0(\scanline[84][4] ),
    .A1(\scanline[85][4] ),
    .A2(\scanline[86][4] ),
    .A3(\scanline[87][4] ),
    .S1(net6182),
    .X(_03805_));
 sg13g2_mux4_1 _20392_ (.S0(net6241),
    .A0(\scanline[92][4] ),
    .A1(\scanline[93][4] ),
    .A2(\scanline[94][4] ),
    .A3(\scanline[95][4] ),
    .S1(net6182),
    .X(_03806_));
 sg13g2_a22oi_1 _20393_ (.Y(_03807_),
    .B1(_03806_),
    .B2(net6097),
    .A2(_03805_),
    .A1(net6065));
 sg13g2_mux4_1 _20394_ (.S0(net6241),
    .A0(\scanline[88][4] ),
    .A1(\scanline[89][4] ),
    .A2(\scanline[90][4] ),
    .A3(\scanline[91][4] ),
    .S1(net6182),
    .X(_03808_));
 sg13g2_mux4_1 _20395_ (.S0(net6239),
    .A0(\scanline[80][4] ),
    .A1(\scanline[81][4] ),
    .A2(\scanline[82][4] ),
    .A3(\scanline[83][4] ),
    .S1(net6179),
    .X(_03809_));
 sg13g2_a22oi_1 _20396_ (.Y(_03810_),
    .B1(_03809_),
    .B2(net6081),
    .A2(_03808_),
    .A1(net6053));
 sg13g2_a21oi_1 _20397_ (.A1(_03807_),
    .A2(_03810_),
    .Y(_03811_),
    .B1(net6012));
 sg13g2_or3_1 _20398_ (.A(_08656_),
    .B(_03804_),
    .C(_03811_),
    .X(_03812_));
 sg13g2_o21ai_1 _20399_ (.B1(_08655_),
    .Y(_03813_),
    .A1(_03797_),
    .A2(_03812_));
 sg13g2_o21ai_1 _20400_ (.B1(_03744_),
    .Y(_03814_),
    .A1(_03773_),
    .A2(_03813_));
 sg13g2_and2_1 _20401_ (.A(net6089),
    .B(_03814_),
    .X(_03815_));
 sg13g2_nand2_1 _20402_ (.Y(_03816_),
    .A(net6089),
    .B(_03814_));
 sg13g2_nor2_1 _20403_ (.A(net5901),
    .B(net5891),
    .Y(_03817_));
 sg13g2_nand2_1 _20404_ (.Y(_03818_),
    .A(net5909),
    .B(net5880));
 sg13g2_and3_2 _20405_ (.X(_03819_),
    .A(net6088),
    .B(net5924),
    .C(net5919));
 sg13g2_nand3_1 _20406_ (.B(net5925),
    .C(_03712_),
    .A(net6087),
    .Y(_03820_));
 sg13g2_nand2_1 _20407_ (.Y(_03821_),
    .A(net5894),
    .B(_03820_));
 sg13g2_nand3_1 _20408_ (.B(net5922),
    .C(_03711_),
    .A(net6086),
    .Y(_03822_));
 sg13g2_nand2_2 _20409_ (.Y(_03823_),
    .A(_03719_),
    .B(_03821_));
 sg13g2_a21oi_1 _20410_ (.A1(net5895),
    .A2(_03820_),
    .Y(_03824_),
    .B1(_03720_));
 sg13g2_a21o_1 _20411_ (.A2(_03820_),
    .A1(net5895),
    .B1(_03720_),
    .X(_03825_));
 sg13g2_a21oi_2 _20412_ (.B1(net5890),
    .Y(_03826_),
    .A2(_03825_),
    .A1(net5901));
 sg13g2_o21ai_1 _20413_ (.B1(_03826_),
    .Y(_03827_),
    .A1(net5900),
    .A2(_03725_));
 sg13g2_nand2_1 _20414_ (.Y(_03828_),
    .A(net5904),
    .B(_03823_));
 sg13g2_nand2_1 _20415_ (.Y(_03829_),
    .A(net5907),
    .B(_03825_));
 sg13g2_a21oi_2 _20416_ (.B1(net5909),
    .Y(_03830_),
    .A2(_03723_),
    .A1(_03618_));
 sg13g2_nand2_1 _20417_ (.Y(_03831_),
    .A(net5900),
    .B(_03725_));
 sg13g2_mux2_1 _20418_ (.A0(_03725_),
    .A1(_03825_),
    .S(net5907),
    .X(_03832_));
 sg13g2_nor2_1 _20419_ (.A(\hvsync_gen.hpos[7] ),
    .B(_09220_),
    .Y(_03833_));
 sg13g2_mux4_1 _20420_ (.S0(net6209),
    .A0(\scanline[144][6] ),
    .A1(\scanline[145][6] ),
    .A2(\scanline[146][6] ),
    .A3(\scanline[147][6] ),
    .S1(net6153),
    .X(_03834_));
 sg13g2_o21ai_1 _20421_ (.B1(net6128),
    .Y(_03835_),
    .A1(net6074),
    .A2(_03834_));
 sg13g2_mux4_1 _20422_ (.S0(net6207),
    .A0(\scanline[156][6] ),
    .A1(\scanline[157][6] ),
    .A2(\scanline[158][6] ),
    .A3(\scanline[159][6] ),
    .S1(net6152),
    .X(_03836_));
 sg13g2_nor2_1 _20423_ (.A(net6090),
    .B(_03836_),
    .Y(_03837_));
 sg13g2_mux4_1 _20424_ (.S0(net6206),
    .A0(\scanline[148][6] ),
    .A1(\scanline[149][6] ),
    .A2(\scanline[150][6] ),
    .A3(\scanline[151][6] ),
    .S1(net6151),
    .X(_03838_));
 sg13g2_nor2_1 _20425_ (.A(net6057),
    .B(_03838_),
    .Y(_03839_));
 sg13g2_mux4_1 _20426_ (.S0(net6206),
    .A0(\scanline[152][6] ),
    .A1(\scanline[153][6] ),
    .A2(\scanline[154][6] ),
    .A3(\scanline[155][6] ),
    .S1(net6151),
    .X(_03840_));
 sg13g2_nor2_1 _20427_ (.A(net6045),
    .B(_03840_),
    .Y(_03841_));
 sg13g2_nor4_1 _20428_ (.A(_03835_),
    .B(_03837_),
    .C(_03839_),
    .D(_03841_),
    .Y(_03842_));
 sg13g2_mux4_1 _20429_ (.S0(net6204),
    .A0(\scanline[128][6] ),
    .A1(\scanline[129][6] ),
    .A2(\scanline[130][6] ),
    .A3(\scanline[131][6] ),
    .S1(net6149),
    .X(_03843_));
 sg13g2_o21ai_1 _20430_ (.B1(net6117),
    .Y(_03844_),
    .A1(net6073),
    .A2(_03843_));
 sg13g2_mux4_1 _20431_ (.S0(net6203),
    .A0(\scanline[140][6] ),
    .A1(\scanline[141][6] ),
    .A2(\scanline[142][6] ),
    .A3(\scanline[143][6] ),
    .S1(net6148),
    .X(_03845_));
 sg13g2_nor2_1 _20432_ (.A(net6090),
    .B(_03845_),
    .Y(_03846_));
 sg13g2_mux4_1 _20433_ (.S0(net6203),
    .A0(\scanline[136][6] ),
    .A1(\scanline[137][6] ),
    .A2(\scanline[138][6] ),
    .A3(\scanline[139][6] ),
    .S1(net6148),
    .X(_03847_));
 sg13g2_nor2_1 _20434_ (.A(net6044),
    .B(_03847_),
    .Y(_03848_));
 sg13g2_mux4_1 _20435_ (.S0(net6202),
    .A0(\scanline[132][6] ),
    .A1(\scanline[133][6] ),
    .A2(\scanline[134][6] ),
    .A3(\scanline[135][6] ),
    .S1(net6147),
    .X(_03849_));
 sg13g2_nor2_1 _20436_ (.A(net6056),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_nor4_2 _20437_ (.A(_03844_),
    .B(_03846_),
    .C(_03848_),
    .Y(_03851_),
    .D(_03850_));
 sg13g2_nor2_2 _20438_ (.A(_03842_),
    .B(_03851_),
    .Y(_03852_));
 sg13g2_nor2b_1 _20439_ (.A(_03852_),
    .B_N(_03833_),
    .Y(_03853_));
 sg13g2_nand2b_1 _20440_ (.Y(_03854_),
    .B(\scanline[100][6] ),
    .A_N(net6237));
 sg13g2_a21oi_1 _20441_ (.A1(net6237),
    .A2(\scanline[101][6] ),
    .Y(_03855_),
    .B1(net6178));
 sg13g2_nand2_1 _20442_ (.Y(_03856_),
    .A(net6237),
    .B(\scanline[103][6] ));
 sg13g2_nand2b_1 _20443_ (.Y(_03857_),
    .B(\scanline[102][6] ),
    .A_N(net6237));
 sg13g2_nand3_1 _20444_ (.B(_03856_),
    .C(_03857_),
    .A(net6171),
    .Y(_03858_));
 sg13g2_a21oi_1 _20445_ (.A1(_03854_),
    .A2(_03855_),
    .Y(_03859_),
    .B1(net6058));
 sg13g2_mux4_1 _20446_ (.S0(net6240),
    .A0(\scanline[108][6] ),
    .A1(\scanline[109][6] ),
    .A2(\scanline[110][6] ),
    .A3(\scanline[111][6] ),
    .S1(net6181),
    .X(_03860_));
 sg13g2_mux4_1 _20447_ (.S0(net6237),
    .A0(\scanline[96][6] ),
    .A1(\scanline[97][6] ),
    .A2(\scanline[98][6] ),
    .A3(\scanline[99][6] ),
    .S1(net6178),
    .X(_03861_));
 sg13g2_mux4_1 _20448_ (.S0(net6235),
    .A0(\scanline[104][6] ),
    .A1(\scanline[105][6] ),
    .A2(\scanline[106][6] ),
    .A3(\scanline[107][6] ),
    .S1(net6177),
    .X(_03862_));
 sg13g2_a22oi_1 _20449_ (.Y(_03863_),
    .B1(_03862_),
    .B2(net6052),
    .A2(_03860_),
    .A1(net6099));
 sg13g2_a221oi_1 _20450_ (.B2(net6080),
    .C1(net6131),
    .B1(_03861_),
    .A1(_03858_),
    .Y(_03864_),
    .A2(_03859_));
 sg13g2_mux4_1 _20451_ (.S0(net6231),
    .A0(\scanline[116][6] ),
    .A1(\scanline[117][6] ),
    .A2(\scanline[118][6] ),
    .A3(\scanline[119][6] ),
    .S1(net6173),
    .X(_03865_));
 sg13g2_and2_1 _20452_ (.A(net6064),
    .B(_03865_),
    .X(_03866_));
 sg13g2_mux4_1 _20453_ (.S0(net6230),
    .A0(\scanline[112][6] ),
    .A1(\scanline[113][6] ),
    .A2(\scanline[114][6] ),
    .A3(\scanline[115][6] ),
    .S1(net6171),
    .X(_03867_));
 sg13g2_mux4_1 _20454_ (.S0(net6232),
    .A0(\scanline[120][6] ),
    .A1(\scanline[121][6] ),
    .A2(\scanline[122][6] ),
    .A3(\scanline[123][6] ),
    .S1(net6174),
    .X(_03868_));
 sg13g2_mux4_1 _20455_ (.S0(net6227),
    .A0(\scanline[124][6] ),
    .A1(\scanline[125][6] ),
    .A2(\scanline[126][6] ),
    .A3(\scanline[127][6] ),
    .S1(net6169),
    .X(_03869_));
 sg13g2_a21oi_1 _20456_ (.A1(net6052),
    .A2(_03868_),
    .Y(_03870_),
    .B1(net6115));
 sg13g2_a221oi_1 _20457_ (.B2(net6099),
    .C1(_03866_),
    .B1(_03869_),
    .A1(net6083),
    .Y(_03871_),
    .A2(_03867_));
 sg13g2_a221oi_1 _20458_ (.B2(_03871_),
    .C1(net6113),
    .B1(_03870_),
    .A1(_03863_),
    .Y(_03872_),
    .A2(_03864_));
 sg13g2_mux4_1 _20459_ (.S0(net6239),
    .A0(\scanline[80][6] ),
    .A1(\scanline[81][6] ),
    .A2(\scanline[82][6] ),
    .A3(\scanline[83][6] ),
    .S1(net6179),
    .X(_03873_));
 sg13g2_mux4_1 _20460_ (.S0(net6241),
    .A0(\scanline[88][6] ),
    .A1(\scanline[89][6] ),
    .A2(\scanline[90][6] ),
    .A3(\scanline[91][6] ),
    .S1(net6182),
    .X(_03874_));
 sg13g2_a22oi_1 _20461_ (.Y(_03875_),
    .B1(_03874_),
    .B2(net6053),
    .A2(_03873_),
    .A1(net6081));
 sg13g2_mux4_1 _20462_ (.S0(net6240),
    .A0(\scanline[92][6] ),
    .A1(\scanline[93][6] ),
    .A2(\scanline[94][6] ),
    .A3(\scanline[95][6] ),
    .S1(net6181),
    .X(_03876_));
 sg13g2_mux4_1 _20463_ (.S0(net6242),
    .A0(\scanline[84][6] ),
    .A1(\scanline[85][6] ),
    .A2(\scanline[86][6] ),
    .A3(\scanline[87][6] ),
    .S1(net6181),
    .X(_03877_));
 sg13g2_a22oi_1 _20464_ (.Y(_03878_),
    .B1(_03877_),
    .B2(net6065),
    .A2(_03876_),
    .A1(net6097));
 sg13g2_a21oi_1 _20465_ (.A1(_03875_),
    .A2(_03878_),
    .Y(_03879_),
    .B1(net6011));
 sg13g2_mux4_1 _20466_ (.S0(net6226),
    .A0(\scanline[64][6] ),
    .A1(\scanline[65][6] ),
    .A2(\scanline[66][6] ),
    .A3(\scanline[67][6] ),
    .S1(net6168),
    .X(_03880_));
 sg13g2_mux4_1 _20467_ (.S0(net6225),
    .A0(\scanline[72][6] ),
    .A1(\scanline[73][6] ),
    .A2(\scanline[74][6] ),
    .A3(\scanline[75][6] ),
    .S1(net6167),
    .X(_03881_));
 sg13g2_a22oi_1 _20468_ (.Y(_03882_),
    .B1(_03881_),
    .B2(net6050),
    .A2(_03880_),
    .A1(net6079));
 sg13g2_mux4_1 _20469_ (.S0(net6222),
    .A0(\scanline[68][6] ),
    .A1(\scanline[69][6] ),
    .A2(\scanline[70][6] ),
    .A3(\scanline[71][6] ),
    .S1(net6165),
    .X(_03883_));
 sg13g2_mux4_1 _20470_ (.S0(net6224),
    .A0(\scanline[76][6] ),
    .A1(\scanline[77][6] ),
    .A2(\scanline[78][6] ),
    .A3(\scanline[79][6] ),
    .S1(net6169),
    .X(_03884_));
 sg13g2_a22oi_1 _20471_ (.Y(_03885_),
    .B1(_03884_),
    .B2(net6095),
    .A2(_03883_),
    .A1(net6066));
 sg13g2_a21oi_2 _20472_ (.B1(net6026),
    .Y(_03886_),
    .A2(_03885_),
    .A1(_03882_));
 sg13g2_or4_2 _20473_ (.A(_08656_),
    .B(_03872_),
    .C(_03879_),
    .D(_03886_),
    .X(_03887_));
 sg13g2_mux2_1 _20474_ (.A0(\scanline[40][6] ),
    .A1(\scanline[41][6] ),
    .S(net6196),
    .X(_03888_));
 sg13g2_nor2_1 _20475_ (.A(net6143),
    .B(_03888_),
    .Y(_03889_));
 sg13g2_mux2_1 _20476_ (.A0(\scanline[42][6] ),
    .A1(\scanline[43][6] ),
    .S(net6196),
    .X(_03890_));
 sg13g2_o21ai_1 _20477_ (.B1(net6047),
    .Y(_03891_),
    .A1(_08652_),
    .A2(_03890_));
 sg13g2_o21ai_1 _20478_ (.B1(net6115),
    .Y(_03892_),
    .A1(_03889_),
    .A2(_03891_));
 sg13g2_mux4_1 _20479_ (.S0(net6211),
    .A0(\scanline[36][6] ),
    .A1(\scanline[37][6] ),
    .A2(\scanline[38][6] ),
    .A3(\scanline[39][6] ),
    .S1(net6156),
    .X(_03893_));
 sg13g2_nand2_1 _20480_ (.Y(_03894_),
    .A(net6063),
    .B(_03893_));
 sg13g2_mux4_1 _20481_ (.S0(net6215),
    .A0(\scanline[32][6] ),
    .A1(\scanline[33][6] ),
    .A2(\scanline[34][6] ),
    .A3(\scanline[35][6] ),
    .S1(net6160),
    .X(_03895_));
 sg13g2_mux4_1 _20482_ (.S0(net6214),
    .A0(\scanline[44][6] ),
    .A1(\scanline[45][6] ),
    .A2(\scanline[46][6] ),
    .A3(\scanline[47][6] ),
    .S1(net6159),
    .X(_03896_));
 sg13g2_a22oi_1 _20483_ (.Y(_03897_),
    .B1(_03896_),
    .B2(net6095),
    .A2(_03895_),
    .A1(net6077));
 sg13g2_nand2_1 _20484_ (.Y(_03898_),
    .A(_03894_),
    .B(_03897_));
 sg13g2_mux4_1 _20485_ (.S0(net6198),
    .A0(\scanline[48][6] ),
    .A1(\scanline[49][6] ),
    .A2(\scanline[50][6] ),
    .A3(\scanline[51][6] ),
    .S1(net6144),
    .X(_03899_));
 sg13g2_mux4_1 _20486_ (.S0(net6199),
    .A0(\scanline[56][6] ),
    .A1(\scanline[57][6] ),
    .A2(\scanline[58][6] ),
    .A3(\scanline[59][6] ),
    .S1(net6146),
    .X(_03900_));
 sg13g2_mux4_1 _20487_ (.S0(net6231),
    .A0(\scanline[52][6] ),
    .A1(\scanline[53][6] ),
    .A2(\scanline[54][6] ),
    .A3(\scanline[55][6] ),
    .S1(net6173),
    .X(_03901_));
 sg13g2_mux4_1 _20488_ (.S0(net6200),
    .A0(\scanline[60][6] ),
    .A1(\scanline[61][6] ),
    .A2(\scanline[62][6] ),
    .A3(\scanline[63][6] ),
    .S1(net6145),
    .X(_03902_));
 sg13g2_a22oi_1 _20489_ (.Y(_03903_),
    .B1(_03900_),
    .B2(net6048),
    .A2(_03899_),
    .A1(net6076));
 sg13g2_a221oi_1 _20490_ (.B2(net6093),
    .C1(net6115),
    .B1(_03902_),
    .A1(net6060),
    .Y(_03904_),
    .A2(_03901_));
 sg13g2_a21oi_1 _20491_ (.A1(_03903_),
    .A2(_03904_),
    .Y(_03905_),
    .B1(net6113));
 sg13g2_o21ai_1 _20492_ (.B1(_03905_),
    .Y(_03906_),
    .A1(_03892_),
    .A2(_03898_));
 sg13g2_mux4_1 _20493_ (.S0(net6186),
    .A0(\scanline[12][6] ),
    .A1(\scanline[13][6] ),
    .A2(\scanline[14][6] ),
    .A3(\scanline[15][6] ),
    .S1(net6135),
    .X(_03907_));
 sg13g2_mux4_1 _20494_ (.S0(net6187),
    .A0(\scanline[4][6] ),
    .A1(\scanline[5][6] ),
    .A2(\scanline[6][6] ),
    .A3(\scanline[7][6] ),
    .S1(net6136),
    .X(_03908_));
 sg13g2_mux4_1 _20495_ (.S0(net6187),
    .A0(\scanline[0][6] ),
    .A1(\scanline[1][6] ),
    .A2(\scanline[2][6] ),
    .A3(\scanline[3][6] ),
    .S1(net6136),
    .X(_03909_));
 sg13g2_mux4_1 _20496_ (.S0(net6187),
    .A0(\scanline[8][6] ),
    .A1(\scanline[9][6] ),
    .A2(\scanline[10][6] ),
    .A3(\scanline[11][6] ),
    .S1(net6136),
    .X(_03910_));
 sg13g2_a22oi_1 _20497_ (.Y(_03911_),
    .B1(_03910_),
    .B2(net6048),
    .A2(_03908_),
    .A1(net6059));
 sg13g2_a22oi_1 _20498_ (.Y(_03912_),
    .B1(_03909_),
    .B2(net6076),
    .A2(_03907_),
    .A1(net6094));
 sg13g2_a21oi_2 _20499_ (.B1(net6025),
    .Y(_03913_),
    .A2(_03912_),
    .A1(_03911_));
 sg13g2_mux4_1 _20500_ (.S0(net6221),
    .A0(\scanline[24][6] ),
    .A1(\scanline[25][6] ),
    .A2(\scanline[26][6] ),
    .A3(\scanline[27][6] ),
    .S1(net6164),
    .X(_03914_));
 sg13g2_mux4_1 _20501_ (.S0(net6221),
    .A0(\scanline[20][6] ),
    .A1(\scanline[21][6] ),
    .A2(\scanline[22][6] ),
    .A3(\scanline[23][6] ),
    .S1(net6164),
    .X(_03915_));
 sg13g2_a22oi_1 _20502_ (.Y(_03916_),
    .B1(_03915_),
    .B2(net6062),
    .A2(_03914_),
    .A1(net6050));
 sg13g2_mux4_1 _20503_ (.S0(net6212),
    .A0(\scanline[16][6] ),
    .A1(\scanline[17][6] ),
    .A2(\scanline[18][6] ),
    .A3(\scanline[19][6] ),
    .S1(net6157),
    .X(_03917_));
 sg13g2_mux4_1 _20504_ (.S0(net6213),
    .A0(\scanline[28][6] ),
    .A1(\scanline[29][6] ),
    .A2(\scanline[30][6] ),
    .A3(\scanline[31][6] ),
    .S1(net6158),
    .X(_03918_));
 sg13g2_a22oi_1 _20505_ (.Y(_03919_),
    .B1(_03918_),
    .B2(net6095),
    .A2(_03917_),
    .A1(net6079));
 sg13g2_a21oi_2 _20506_ (.B1(net6011),
    .Y(_03920_),
    .A2(_03919_),
    .A1(_03916_));
 sg13g2_nor3_2 _20507_ (.A(net6127),
    .B(_03913_),
    .C(_03920_),
    .Y(_03921_));
 sg13g2_a21oi_2 _20508_ (.B1(\hvsync_gen.hpos[9] ),
    .Y(_03922_),
    .A2(_03921_),
    .A1(_03906_));
 sg13g2_a21oi_2 _20509_ (.B1(_03853_),
    .Y(_03923_),
    .A2(_03922_),
    .A1(_03887_));
 sg13g2_a21o_2 _20510_ (.A2(_03922_),
    .A1(_03887_),
    .B1(_03853_),
    .X(_03924_));
 sg13g2_mux4_1 _20511_ (.S0(net6207),
    .A0(\scanline[156][5] ),
    .A1(\scanline[157][5] ),
    .A2(\scanline[158][5] ),
    .A3(\scanline[159][5] ),
    .S1(net6152),
    .X(_03925_));
 sg13g2_o21ai_1 _20512_ (.B1(net6128),
    .Y(_03926_),
    .A1(net6091),
    .A2(_03925_));
 sg13g2_mux4_1 _20513_ (.S0(net6209),
    .A0(\scanline[144][5] ),
    .A1(\scanline[145][5] ),
    .A2(\scanline[146][5] ),
    .A3(\scanline[147][5] ),
    .S1(net6153),
    .X(_03927_));
 sg13g2_nor2_1 _20514_ (.A(net6073),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_mux4_1 _20515_ (.S0(net6206),
    .A0(\scanline[148][5] ),
    .A1(\scanline[149][5] ),
    .A2(\scanline[150][5] ),
    .A3(\scanline[151][5] ),
    .S1(net6151),
    .X(_03929_));
 sg13g2_nor2_1 _20516_ (.A(net6056),
    .B(_03929_),
    .Y(_03930_));
 sg13g2_mux4_1 _20517_ (.S0(net6206),
    .A0(\scanline[152][5] ),
    .A1(\scanline[153][5] ),
    .A2(\scanline[154][5] ),
    .A3(\scanline[155][5] ),
    .S1(net6151),
    .X(_03931_));
 sg13g2_nor2_1 _20518_ (.A(net6045),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_nor4_2 _20519_ (.A(_03926_),
    .B(_03928_),
    .C(_03930_),
    .Y(_03933_),
    .D(_03932_));
 sg13g2_mux4_1 _20520_ (.S0(net6186),
    .A0(\scanline[132][5] ),
    .A1(\scanline[133][5] ),
    .A2(\scanline[134][5] ),
    .A3(\scanline[135][5] ),
    .S1(net6135),
    .X(_03934_));
 sg13g2_o21ai_1 _20521_ (.B1(net6117),
    .Y(_03935_),
    .A1(net6056),
    .A2(_03934_));
 sg13g2_mux4_1 _20522_ (.S0(net6204),
    .A0(\scanline[128][5] ),
    .A1(\scanline[129][5] ),
    .A2(\scanline[130][5] ),
    .A3(\scanline[131][5] ),
    .S1(net6149),
    .X(_03936_));
 sg13g2_nor2_1 _20523_ (.A(net6073),
    .B(_03936_),
    .Y(_03937_));
 sg13g2_mux4_1 _20524_ (.S0(net6190),
    .A0(\scanline[136][5] ),
    .A1(\scanline[137][5] ),
    .A2(\scanline[138][5] ),
    .A3(\scanline[139][5] ),
    .S1(net6138),
    .X(_03938_));
 sg13g2_nor2_1 _20525_ (.A(net6044),
    .B(_03938_),
    .Y(_03939_));
 sg13g2_mux4_1 _20526_ (.S0(net6203),
    .A0(\scanline[140][5] ),
    .A1(\scanline[141][5] ),
    .A2(\scanline[142][5] ),
    .A3(\scanline[143][5] ),
    .S1(net6148),
    .X(_03940_));
 sg13g2_nor2_1 _20527_ (.A(net6091),
    .B(_03940_),
    .Y(_03941_));
 sg13g2_nor4_2 _20528_ (.A(_03935_),
    .B(_03937_),
    .C(_03939_),
    .Y(_03942_),
    .D(_03941_));
 sg13g2_o21ai_1 _20529_ (.B1(_03833_),
    .Y(_03943_),
    .A1(_03933_),
    .A2(_03942_));
 sg13g2_nand2b_1 _20530_ (.Y(_03944_),
    .B(\scanline[60][5] ),
    .A_N(net6200));
 sg13g2_a21oi_1 _20531_ (.A1(net6200),
    .A2(\scanline[61][5] ),
    .Y(_03945_),
    .B1(net6145));
 sg13g2_nand2_1 _20532_ (.Y(_03946_),
    .A(net6200),
    .B(\scanline[63][5] ));
 sg13g2_nand2b_1 _20533_ (.Y(_03947_),
    .B(\scanline[62][5] ),
    .A_N(net6200));
 sg13g2_nand3_1 _20534_ (.B(_03946_),
    .C(_03947_),
    .A(net6145),
    .Y(_03948_));
 sg13g2_a21oi_1 _20535_ (.A1(_03944_),
    .A2(_03945_),
    .Y(_03949_),
    .B1(net6092));
 sg13g2_mux4_1 _20536_ (.S0(net6200),
    .A0(\scanline[56][5] ),
    .A1(\scanline[57][5] ),
    .A2(\scanline[58][5] ),
    .A3(\scanline[59][5] ),
    .S1(net6145),
    .X(_03950_));
 sg13g2_mux4_1 _20537_ (.S0(net6216),
    .A0(\scanline[52][5] ),
    .A1(\scanline[53][5] ),
    .A2(\scanline[54][5] ),
    .A3(\scanline[55][5] ),
    .S1(net6161),
    .X(_03951_));
 sg13g2_mux4_1 _20538_ (.S0(net6198),
    .A0(\scanline[48][5] ),
    .A1(\scanline[49][5] ),
    .A2(\scanline[50][5] ),
    .A3(\scanline[51][5] ),
    .S1(net6144),
    .X(_03952_));
 sg13g2_a22oi_1 _20539_ (.Y(_03953_),
    .B1(_03950_),
    .B2(net6049),
    .A2(_03949_),
    .A1(_03948_));
 sg13g2_a221oi_1 _20540_ (.B2(net6077),
    .C1(net6115),
    .B1(_03952_),
    .A1(net6059),
    .Y(_03954_),
    .A2(_03951_));
 sg13g2_mux4_1 _20541_ (.S0(net6211),
    .A0(\scanline[44][5] ),
    .A1(\scanline[45][5] ),
    .A2(\scanline[46][5] ),
    .A3(\scanline[47][5] ),
    .S1(net6156),
    .X(_03955_));
 sg13g2_mux4_1 _20542_ (.S0(net6195),
    .A0(\scanline[40][5] ),
    .A1(\scanline[41][5] ),
    .A2(\scanline[42][5] ),
    .A3(\scanline[43][5] ),
    .S1(net6142),
    .X(_03956_));
 sg13g2_mux4_1 _20543_ (.S0(net6211),
    .A0(\scanline[36][5] ),
    .A1(\scanline[37][5] ),
    .A2(\scanline[38][5] ),
    .A3(\scanline[39][5] ),
    .S1(net6156),
    .X(_03957_));
 sg13g2_mux4_1 _20544_ (.S0(net6211),
    .A0(\scanline[32][5] ),
    .A1(\scanline[33][5] ),
    .A2(\scanline[34][5] ),
    .A3(\scanline[35][5] ),
    .S1(net6156),
    .X(_03958_));
 sg13g2_a22oi_1 _20545_ (.Y(_03959_),
    .B1(_03958_),
    .B2(net6077),
    .A2(_03957_),
    .A1(net6063));
 sg13g2_a221oi_1 _20546_ (.B2(net6047),
    .C1(net6131),
    .B1(_03956_),
    .A1(net6093),
    .Y(_03960_),
    .A2(_03955_));
 sg13g2_a221oi_1 _20547_ (.B2(_03960_),
    .C1(net6113),
    .B1(_03959_),
    .A1(_03953_),
    .Y(_03961_),
    .A2(_03954_));
 sg13g2_mux4_1 _20548_ (.S0(net6213),
    .A0(\scanline[28][5] ),
    .A1(\scanline[29][5] ),
    .A2(\scanline[30][5] ),
    .A3(\scanline[31][5] ),
    .S1(net6158),
    .X(_03962_));
 sg13g2_mux4_1 _20549_ (.S0(net6223),
    .A0(\scanline[24][5] ),
    .A1(\scanline[25][5] ),
    .A2(\scanline[26][5] ),
    .A3(\scanline[27][5] ),
    .S1(net6166),
    .X(_03963_));
 sg13g2_a22oi_1 _20550_ (.Y(_03964_),
    .B1(_03963_),
    .B2(net6051),
    .A2(_03962_),
    .A1(net6096));
 sg13g2_mux4_1 _20551_ (.S0(net6212),
    .A0(\scanline[20][5] ),
    .A1(\scanline[21][5] ),
    .A2(\scanline[22][5] ),
    .A3(\scanline[23][5] ),
    .S1(net6157),
    .X(_03965_));
 sg13g2_mux4_1 _20552_ (.S0(net6212),
    .A0(\scanline[16][5] ),
    .A1(\scanline[17][5] ),
    .A2(\scanline[18][5] ),
    .A3(\scanline[19][5] ),
    .S1(net6157),
    .X(_03966_));
 sg13g2_a22oi_1 _20553_ (.Y(_03967_),
    .B1(_03966_),
    .B2(net6079),
    .A2(_03965_),
    .A1(net6063));
 sg13g2_a21oi_2 _20554_ (.B1(net6011),
    .Y(_03968_),
    .A2(_03967_),
    .A1(_03964_));
 sg13g2_mux4_1 _20555_ (.S0(net6194),
    .A0(\scanline[8][5] ),
    .A1(\scanline[9][5] ),
    .A2(\scanline[10][5] ),
    .A3(\scanline[11][5] ),
    .S1(net6141),
    .X(_03969_));
 sg13g2_mux4_1 _20556_ (.S0(net6186),
    .A0(\scanline[12][5] ),
    .A1(\scanline[13][5] ),
    .A2(\scanline[14][5] ),
    .A3(\scanline[15][5] ),
    .S1(net6135),
    .X(_03970_));
 sg13g2_mux4_1 _20557_ (.S0(net6193),
    .A0(\scanline[0][5] ),
    .A1(\scanline[1][5] ),
    .A2(\scanline[2][5] ),
    .A3(\scanline[3][5] ),
    .S1(net6141),
    .X(_03971_));
 sg13g2_mux4_1 _20558_ (.S0(net6186),
    .A0(\scanline[4][5] ),
    .A1(\scanline[5][5] ),
    .A2(\scanline[6][5] ),
    .A3(\scanline[7][5] ),
    .S1(net6135),
    .X(_03972_));
 sg13g2_a22oi_1 _20559_ (.Y(_03973_),
    .B1(_03972_),
    .B2(net6059),
    .A2(_03970_),
    .A1(net6094));
 sg13g2_a22oi_1 _20560_ (.Y(_03974_),
    .B1(_03971_),
    .B2(net6076),
    .A2(_03969_),
    .A1(net6048));
 sg13g2_a21oi_2 _20561_ (.B1(net6025),
    .Y(_03975_),
    .A2(_03974_),
    .A1(_03973_));
 sg13g2_or4_2 _20562_ (.A(net6127),
    .B(_03961_),
    .C(_03968_),
    .D(_03975_),
    .X(_03976_));
 sg13g2_nor2b_1 _20563_ (.A(net6217),
    .B_N(\scanline[124][5] ),
    .Y(_03977_));
 sg13g2_a21oi_1 _20564_ (.A1(net6217),
    .A2(\scanline[125][5] ),
    .Y(_03978_),
    .B1(_03977_));
 sg13g2_nand2b_1 _20565_ (.Y(_03979_),
    .B(\scanline[126][5] ),
    .A_N(net6217));
 sg13g2_a21oi_1 _20566_ (.A1(net6217),
    .A2(\scanline[127][5] ),
    .Y(_03980_),
    .B1(_08652_));
 sg13g2_a221oi_1 _20567_ (.B2(_03980_),
    .C1(net6092),
    .B1(_03979_),
    .A1(_08652_),
    .Y(_03981_),
    .A2(_03978_));
 sg13g2_mux4_1 _20568_ (.S0(net6230),
    .A0(\scanline[112][5] ),
    .A1(\scanline[113][5] ),
    .A2(\scanline[114][5] ),
    .A3(\scanline[115][5] ),
    .S1(net6171),
    .X(_03982_));
 sg13g2_nand2_1 _20569_ (.Y(_03983_),
    .A(net6083),
    .B(_03982_));
 sg13g2_mux4_1 _20570_ (.S0(net6233),
    .A0(\scanline[120][5] ),
    .A1(\scanline[121][5] ),
    .A2(\scanline[122][5] ),
    .A3(\scanline[123][5] ),
    .S1(net6174),
    .X(_03984_));
 sg13g2_mux4_1 _20571_ (.S0(net6233),
    .A0(\scanline[116][5] ),
    .A1(\scanline[117][5] ),
    .A2(\scanline[118][5] ),
    .A3(\scanline[119][5] ),
    .S1(net6175),
    .X(_03985_));
 sg13g2_a22oi_1 _20572_ (.Y(_03986_),
    .B1(_03985_),
    .B2(net6064),
    .A2(_03984_),
    .A1(net6049));
 sg13g2_nand2_1 _20573_ (.Y(_03987_),
    .A(_03983_),
    .B(_03986_));
 sg13g2_nor3_1 _20574_ (.A(net6116),
    .B(_03981_),
    .C(_03987_),
    .Y(_03988_));
 sg13g2_mux4_1 _20575_ (.S0(net6229),
    .A0(\scanline[108][5] ),
    .A1(\scanline[109][5] ),
    .A2(\scanline[110][5] ),
    .A3(\scanline[111][5] ),
    .S1(net6171),
    .X(_03989_));
 sg13g2_mux4_1 _20576_ (.S0(net6237),
    .A0(\scanline[96][5] ),
    .A1(\scanline[97][5] ),
    .A2(\scanline[98][5] ),
    .A3(\scanline[99][5] ),
    .S1(net6178),
    .X(_03990_));
 sg13g2_mux4_1 _20577_ (.S0(net6234),
    .A0(\scanline[104][5] ),
    .A1(\scanline[105][5] ),
    .A2(\scanline[106][5] ),
    .A3(\scanline[107][5] ),
    .S1(net6176),
    .X(_03991_));
 sg13g2_nand2_1 _20578_ (.Y(_03992_),
    .A(net6052),
    .B(_03991_));
 sg13g2_mux2_1 _20579_ (.A0(\scanline[100][5] ),
    .A1(\scanline[101][5] ),
    .S(net6230),
    .X(_03993_));
 sg13g2_nor2_1 _20580_ (.A(net6171),
    .B(_03993_),
    .Y(_03994_));
 sg13g2_mux2_1 _20581_ (.A0(\scanline[102][5] ),
    .A1(\scanline[103][5] ),
    .S(net6217),
    .X(_03995_));
 sg13g2_o21ai_1 _20582_ (.B1(net6064),
    .Y(_03996_),
    .A1(_08652_),
    .A2(_03995_));
 sg13g2_o21ai_1 _20583_ (.B1(_03992_),
    .Y(_03997_),
    .A1(_03994_),
    .A2(_03996_));
 sg13g2_a221oi_1 _20584_ (.B2(net6080),
    .C1(net6131),
    .B1(_03990_),
    .A1(net6097),
    .Y(_03998_),
    .A2(_03989_));
 sg13g2_inv_1 _20585_ (.Y(_03999_),
    .A(_03998_));
 sg13g2_o21ai_1 _20586_ (.B1(\hvsync_gen.hpos[7] ),
    .Y(_04000_),
    .A1(_03997_),
    .A2(_03999_));
 sg13g2_mux4_1 _20587_ (.S0(net6242),
    .A0(\scanline[88][5] ),
    .A1(\scanline[89][5] ),
    .A2(\scanline[90][5] ),
    .A3(\scanline[91][5] ),
    .S1(net6183),
    .X(_04001_));
 sg13g2_mux4_1 _20588_ (.S0(net6239),
    .A0(\scanline[80][5] ),
    .A1(\scanline[81][5] ),
    .A2(\scanline[82][5] ),
    .A3(\scanline[83][5] ),
    .S1(net6179),
    .X(_04002_));
 sg13g2_mux4_1 _20589_ (.S0(net6240),
    .A0(\scanline[84][5] ),
    .A1(\scanline[85][5] ),
    .A2(\scanline[86][5] ),
    .A3(\scanline[87][5] ),
    .S1(net6181),
    .X(_04003_));
 sg13g2_mux4_1 _20590_ (.S0(net6239),
    .A0(\scanline[92][5] ),
    .A1(\scanline[93][5] ),
    .A2(\scanline[94][5] ),
    .A3(\scanline[95][5] ),
    .S1(net6179),
    .X(_04004_));
 sg13g2_a22oi_1 _20591_ (.Y(_04005_),
    .B1(_04004_),
    .B2(net6097),
    .A2(_04002_),
    .A1(net6081));
 sg13g2_a22oi_1 _20592_ (.Y(_04006_),
    .B1(_04003_),
    .B2(net6065),
    .A2(_04001_),
    .A1(net6053));
 sg13g2_a21oi_1 _20593_ (.A1(_04005_),
    .A2(_04006_),
    .Y(_04007_),
    .B1(net6011));
 sg13g2_mux4_1 _20594_ (.S0(net6223),
    .A0(\scanline[72][5] ),
    .A1(\scanline[73][5] ),
    .A2(\scanline[74][5] ),
    .A3(\scanline[75][5] ),
    .S1(net6166),
    .X(_04008_));
 sg13g2_mux4_1 _20595_ (.S0(net6222),
    .A0(\scanline[68][5] ),
    .A1(\scanline[69][5] ),
    .A2(\scanline[70][5] ),
    .A3(\scanline[71][5] ),
    .S1(net6165),
    .X(_04009_));
 sg13g2_a22oi_1 _20596_ (.Y(_04010_),
    .B1(_04009_),
    .B2(net6062),
    .A2(_04008_),
    .A1(net6050));
 sg13g2_mux4_1 _20597_ (.S0(net6226),
    .A0(\scanline[64][5] ),
    .A1(\scanline[65][5] ),
    .A2(\scanline[66][5] ),
    .A3(\scanline[67][5] ),
    .S1(net6168),
    .X(_04011_));
 sg13g2_mux4_1 _20598_ (.S0(net6226),
    .A0(\scanline[76][5] ),
    .A1(\scanline[77][5] ),
    .A2(\scanline[78][5] ),
    .A3(\scanline[79][5] ),
    .S1(net6167),
    .X(_04012_));
 sg13g2_a22oi_1 _20599_ (.Y(_04013_),
    .B1(_04012_),
    .B2(net6097),
    .A2(_04011_),
    .A1(net6081));
 sg13g2_a21oi_2 _20600_ (.B1(net6025),
    .Y(_04014_),
    .A2(_04013_),
    .A1(_04010_));
 sg13g2_nor3_2 _20601_ (.A(_08656_),
    .B(_04007_),
    .C(_04014_),
    .Y(_04015_));
 sg13g2_o21ai_1 _20602_ (.B1(_04015_),
    .Y(_04016_),
    .A1(_03988_),
    .A2(_04000_));
 sg13g2_nand3_1 _20603_ (.B(_03976_),
    .C(_04016_),
    .A(_08655_),
    .Y(_04017_));
 sg13g2_nand2_2 _20604_ (.Y(_04018_),
    .A(_03943_),
    .B(_04017_));
 sg13g2_inv_1 _20605_ (.Y(_04019_),
    .A(_04018_));
 sg13g2_nand2_2 _20606_ (.Y(_04020_),
    .A(net5918),
    .B(_04018_));
 sg13g2_inv_2 _20607_ (.Y(_04021_),
    .A(_04020_));
 sg13g2_a21oi_1 _20608_ (.A1(net5890),
    .A2(_03832_),
    .Y(_04022_),
    .B1(_04020_));
 sg13g2_nor2_2 _20609_ (.A(net5918),
    .B(net5849),
    .Y(_04023_));
 sg13g2_nand2_2 _20610_ (.Y(_04024_),
    .A(_03923_),
    .B(_04018_));
 sg13g2_nand4_1 _20611_ (.B(net5925),
    .C(net5921),
    .A(net6087),
    .Y(_04025_),
    .D(_03711_));
 sg13g2_nor3_2 _20612_ (.A(_09227_),
    .B(net5921),
    .C(_03711_),
    .Y(_04026_));
 sg13g2_or2_2 _20613_ (.X(_04027_),
    .B(_03713_),
    .A(net5920));
 sg13g2_nor2_1 _20614_ (.A(net5898),
    .B(_04026_),
    .Y(_04028_));
 sg13g2_and2_1 _20615_ (.A(net5907),
    .B(_04025_),
    .X(_04029_));
 sg13g2_nand2_1 _20616_ (.Y(_04030_),
    .A(_04027_),
    .B(_04029_));
 sg13g2_a21oi_1 _20617_ (.A1(_04027_),
    .A2(_04029_),
    .Y(_04031_),
    .B1(net5885));
 sg13g2_o21ai_1 _20618_ (.B1(net6088),
    .Y(_04032_),
    .A1(net5924),
    .A2(net5919));
 sg13g2_o21ai_1 _20619_ (.B1(net6085),
    .Y(_04033_),
    .A1(net5924),
    .A2(net5920));
 sg13g2_nand2_2 _20620_ (.Y(_04034_),
    .A(net5894),
    .B(_03717_));
 sg13g2_nor2_1 _20621_ (.A(_03716_),
    .B(_03819_),
    .Y(_04035_));
 sg13g2_nor2_2 _20622_ (.A(_03711_),
    .B(_04033_),
    .Y(_04036_));
 sg13g2_o21ai_1 _20623_ (.B1(net5900),
    .Y(_04037_),
    .A1(_03718_),
    .A2(_04036_));
 sg13g2_nor2_2 _20624_ (.A(_03718_),
    .B(net5890),
    .Y(_04038_));
 sg13g2_nor3_2 _20625_ (.A(_09227_),
    .B(net5925),
    .C(_03711_),
    .Y(_04039_));
 sg13g2_nor4_2 _20626_ (.A(_09227_),
    .B(net5925),
    .C(net5921),
    .Y(_04040_),
    .D(_03711_));
 sg13g2_nor3_1 _20627_ (.A(_03718_),
    .B(net5890),
    .C(_04040_),
    .Y(_04041_));
 sg13g2_a21o_1 _20628_ (.A2(_04037_),
    .A1(_04031_),
    .B1(_04041_),
    .X(_04042_));
 sg13g2_and3_1 _20629_ (.X(_04043_),
    .A(_03923_),
    .B(_03943_),
    .C(_04017_));
 sg13g2_nand2_2 _20630_ (.Y(_04044_),
    .A(_03923_),
    .B(_04019_));
 sg13g2_a22oi_1 _20631_ (.Y(_04045_),
    .B1(_03830_),
    .B2(_04038_),
    .A2(_03824_),
    .A1(_03817_));
 sg13g2_nand2b_1 _20632_ (.Y(_04046_),
    .B(net5878),
    .A_N(_04045_));
 sg13g2_nand2_1 _20633_ (.Y(_04047_),
    .A(net5897),
    .B(net5894));
 sg13g2_o21ai_1 _20634_ (.B1(net6086),
    .Y(_04048_),
    .A1(net5922),
    .A2(net5919));
 sg13g2_nand2_2 _20635_ (.Y(_04049_),
    .A(_03713_),
    .B(net5894));
 sg13g2_a221oi_1 _20636_ (.B2(net5921),
    .C1(_09227_),
    .B1(net5925),
    .A1(_03352_),
    .Y(_04050_),
    .A2(_03433_));
 sg13g2_nand2_2 _20637_ (.Y(_04051_),
    .A(net5904),
    .B(_03719_));
 sg13g2_mux2_1 _20638_ (.A0(net5876),
    .A1(net5900),
    .S(_04048_),
    .X(_04052_));
 sg13g2_nand2_2 _20639_ (.Y(_04053_),
    .A(net5888),
    .B(net5849));
 sg13g2_and2_1 _20640_ (.A(net5890),
    .B(net5878),
    .X(_04054_));
 sg13g2_nand2_1 _20641_ (.Y(_04055_),
    .A(net5890),
    .B(net5878));
 sg13g2_nor2_2 _20642_ (.A(_03923_),
    .B(_04018_),
    .Y(_04056_));
 sg13g2_inv_1 _20643_ (.Y(_04057_),
    .A(_04056_));
 sg13g2_nor2_1 _20644_ (.A(_03716_),
    .B(_04039_),
    .Y(_04058_));
 sg13g2_a22oi_1 _20645_ (.Y(_04059_),
    .B1(net5848),
    .B2(_04058_),
    .A2(_04054_),
    .A1(_04052_));
 sg13g2_o21ai_1 _20646_ (.B1(_04059_),
    .Y(_04060_),
    .A1(_04044_),
    .A2(_04045_));
 sg13g2_a221oi_1 _20647_ (.B2(_04042_),
    .C1(_04060_),
    .B1(_04023_),
    .A1(_03827_),
    .Y(_04061_),
    .A2(_04022_));
 sg13g2_nand2_1 _20648_ (.Y(_04062_),
    .A(net7563),
    .B(net6017));
 sg13g2_and3_1 _20649_ (.X(_04063_),
    .A(net7563),
    .B(net6016),
    .C(_04061_));
 sg13g2_inv_1 _20650_ (.Y(_04064_),
    .A(_04063_));
 sg13g2_nor2b_1 _20651_ (.A(_04061_),
    .B_N(_04062_),
    .Y(_04065_));
 sg13g2_nor3_1 _20652_ (.A(net5987),
    .B(_04063_),
    .C(_04065_),
    .Y(_00303_));
 sg13g2_nand2_1 _20653_ (.Y(_04066_),
    .A(\r_pwm_odd[4] ),
    .B(net6017));
 sg13g2_nor2_1 _20654_ (.A(net5904),
    .B(_04034_),
    .Y(_04067_));
 sg13g2_or2_1 _20655_ (.X(_04068_),
    .B(net5879),
    .A(net5896));
 sg13g2_nor2_2 _20656_ (.A(_03819_),
    .B(_04032_),
    .Y(_04069_));
 sg13g2_nor3_2 _20657_ (.A(net5896),
    .B(_03819_),
    .C(net5879),
    .Y(_04070_));
 sg13g2_or3_2 _20658_ (.A(net5896),
    .B(_03819_),
    .C(_04032_),
    .X(_04071_));
 sg13g2_a21oi_1 _20659_ (.A1(net5876),
    .A2(_04071_),
    .Y(_04072_),
    .B1(net5883));
 sg13g2_a221oi_1 _20660_ (.B2(_04071_),
    .C1(net5883),
    .B1(net5876),
    .A1(net5902),
    .Y(_04073_),
    .A2(_04033_));
 sg13g2_nand2_1 _20661_ (.Y(_04074_),
    .A(_03822_),
    .B(net5876));
 sg13g2_o21ai_1 _20662_ (.B1(net5898),
    .Y(_04075_),
    .A1(_04026_),
    .A2(net5879));
 sg13g2_and3_1 _20663_ (.X(_04076_),
    .A(net5883),
    .B(_04074_),
    .C(_04075_));
 sg13g2_nor3_1 _20664_ (.A(_04044_),
    .B(_04073_),
    .C(_04076_),
    .Y(_04077_));
 sg13g2_nor2_2 _20665_ (.A(net5905),
    .B(net5880),
    .Y(_04078_));
 sg13g2_nand2_2 _20666_ (.Y(_04079_),
    .A(net5897),
    .B(net5888));
 sg13g2_or2_1 _20667_ (.X(_04080_),
    .B(_04039_),
    .A(net5896));
 sg13g2_nor2_1 _20668_ (.A(net5899),
    .B(net5880),
    .Y(_04081_));
 sg13g2_and2_2 _20669_ (.A(_03717_),
    .B(_03822_),
    .X(_04082_));
 sg13g2_nand2_1 _20670_ (.Y(_04083_),
    .A(net5847),
    .B(_04082_));
 sg13g2_a22oi_1 _20671_ (.Y(_04084_),
    .B1(_04078_),
    .B2(_04080_),
    .A2(_04038_),
    .A1(_04034_));
 sg13g2_a21oi_1 _20672_ (.A1(_04083_),
    .A2(_04084_),
    .Y(_04085_),
    .B1(_04024_));
 sg13g2_o21ai_1 _20673_ (.B1(net5894),
    .Y(_04086_),
    .A1(_03819_),
    .A2(net5879));
 sg13g2_a21oi_1 _20674_ (.A1(_03719_),
    .A2(net5846),
    .Y(_04087_),
    .B1(_04057_));
 sg13g2_o21ai_1 _20675_ (.B1(net5902),
    .Y(_04088_),
    .A1(_03716_),
    .A2(_03819_));
 sg13g2_a21oi_1 _20676_ (.A1(_03822_),
    .A2(net5876),
    .Y(_04089_),
    .B1(net5884));
 sg13g2_a221oi_1 _20677_ (.B2(_04089_),
    .C1(_04020_),
    .B1(_04088_),
    .A1(net5884),
    .Y(_04090_),
    .A2(_04036_));
 sg13g2_or4_2 _20678_ (.A(_04077_),
    .B(_04085_),
    .C(_04087_),
    .D(_04090_),
    .X(_04091_));
 sg13g2_inv_1 _20679_ (.Y(_04092_),
    .A(_04091_));
 sg13g2_nor2_1 _20680_ (.A(_04061_),
    .B(_04091_),
    .Y(_04093_));
 sg13g2_xor2_1 _20681_ (.B(_04091_),
    .A(_04061_),
    .X(_04094_));
 sg13g2_xnor2_1 _20682_ (.Y(_04095_),
    .A(_04061_),
    .B(_04091_));
 sg13g2_nand2b_1 _20683_ (.Y(_04096_),
    .B(_04095_),
    .A_N(_04066_));
 sg13g2_xnor2_1 _20684_ (.Y(_04097_),
    .A(_04066_),
    .B(_04094_));
 sg13g2_xnor2_1 _20685_ (.Y(_04098_),
    .A(_04064_),
    .B(_04097_));
 sg13g2_nor2_1 _20686_ (.A(net5987),
    .B(_04098_),
    .Y(_00304_));
 sg13g2_o21ai_1 _20687_ (.B1(_04096_),
    .Y(_04099_),
    .A1(_04064_),
    .A2(_04097_));
 sg13g2_nand2_1 _20688_ (.Y(_04100_),
    .A(\r_pwm_odd[5] ),
    .B(net6016));
 sg13g2_nor2_2 _20689_ (.A(net5894),
    .B(net5879),
    .Y(_04101_));
 sg13g2_nand3b_1 _20690_ (.B(net5896),
    .C(_03820_),
    .Y(_04102_),
    .A_N(net5879));
 sg13g2_nand3_1 _20691_ (.B(net5846),
    .C(_04102_),
    .A(net5901),
    .Y(_04103_));
 sg13g2_o21ai_1 _20692_ (.B1(net5896),
    .Y(_04104_),
    .A1(_03819_),
    .A2(net5879));
 sg13g2_nand3_1 _20693_ (.B(_04071_),
    .C(net5845),
    .A(net5905),
    .Y(_04105_));
 sg13g2_nand3_1 _20694_ (.B(_04103_),
    .C(_04105_),
    .A(net5885),
    .Y(_04106_));
 sg13g2_and3_1 _20695_ (.X(_04107_),
    .A(net5906),
    .B(_03721_),
    .C(_04025_));
 sg13g2_nand3_1 _20696_ (.B(net5893),
    .C(_04025_),
    .A(net5908),
    .Y(_04108_));
 sg13g2_nor2_1 _20697_ (.A(_03716_),
    .B(_03724_),
    .Y(_04109_));
 sg13g2_nor2_1 _20698_ (.A(net5885),
    .B(_04107_),
    .Y(_04110_));
 sg13g2_o21ai_1 _20699_ (.B1(_04110_),
    .Y(_04111_),
    .A1(net5906),
    .A2(_04109_));
 sg13g2_a21o_1 _20700_ (.A2(_04111_),
    .A1(_04106_),
    .B1(_04024_),
    .X(_04112_));
 sg13g2_nor2b_1 _20701_ (.A(_03434_),
    .B_N(_03723_),
    .Y(_04113_));
 sg13g2_and3_1 _20702_ (.X(_04114_),
    .A(net5902),
    .B(_03717_),
    .C(_03822_));
 sg13g2_nor3_2 _20703_ (.A(net5892),
    .B(_04113_),
    .C(_04114_),
    .Y(_04115_));
 sg13g2_nor3_1 _20704_ (.A(net5900),
    .B(_03723_),
    .C(_04082_),
    .Y(_04116_));
 sg13g2_nand2b_1 _20705_ (.Y(_04117_),
    .B(_04115_),
    .A_N(_04116_));
 sg13g2_nand3b_1 _20706_ (.B(net5920),
    .C(net6085),
    .Y(_04118_),
    .A_N(net5924));
 sg13g2_nand3b_1 _20707_ (.B(_04118_),
    .C(net5907),
    .Y(_04119_),
    .A_N(_03716_));
 sg13g2_and2_1 _20708_ (.A(net5899),
    .B(_04118_),
    .X(_04120_));
 sg13g2_nand2_1 _20709_ (.Y(_04121_),
    .A(net5901),
    .B(_04118_));
 sg13g2_nand3_1 _20710_ (.B(_04119_),
    .C(_04121_),
    .A(net5891),
    .Y(_04122_));
 sg13g2_nand3_1 _20711_ (.B(_04117_),
    .C(_04122_),
    .A(_04021_),
    .Y(_04123_));
 sg13g2_nand3b_1 _20712_ (.B(net5845),
    .C(net5906),
    .Y(_04124_),
    .A_N(_04040_));
 sg13g2_o21ai_1 _20713_ (.B1(net5892),
    .Y(_04125_),
    .A1(_03434_),
    .A2(_03713_));
 sg13g2_nand2b_1 _20714_ (.Y(_04126_),
    .B(_04124_),
    .A_N(_04125_));
 sg13g2_a221oi_1 _20715_ (.B2(net5924),
    .C1(net5908),
    .B1(_04026_),
    .A1(_03711_),
    .Y(_04127_),
    .A2(_03714_));
 sg13g2_nor2_1 _20716_ (.A(net5891),
    .B(_04127_),
    .Y(_04128_));
 sg13g2_nand2_1 _20717_ (.Y(_04129_),
    .A(_04119_),
    .B(_04128_));
 sg13g2_nand3_1 _20718_ (.B(_04126_),
    .C(_04129_),
    .A(net5877),
    .Y(_04130_));
 sg13g2_nor2_1 _20719_ (.A(_03722_),
    .B(_04069_),
    .Y(_04131_));
 sg13g2_nand2_1 _20720_ (.Y(_04132_),
    .A(_04056_),
    .B(_04131_));
 sg13g2_and4_2 _20721_ (.A(_04112_),
    .B(_04123_),
    .C(_04130_),
    .D(_04132_),
    .X(_04133_));
 sg13g2_xnor2_1 _20722_ (.Y(_04134_),
    .A(_04093_),
    .B(_04133_));
 sg13g2_nor2_1 _20723_ (.A(_04100_),
    .B(_04134_),
    .Y(_04135_));
 sg13g2_nand2_1 _20724_ (.Y(_04136_),
    .A(_04100_),
    .B(_04134_));
 sg13g2_xnor2_1 _20725_ (.Y(_04137_),
    .A(_04100_),
    .B(_04134_));
 sg13g2_xnor2_1 _20726_ (.Y(_04138_),
    .A(_04099_),
    .B(_04137_));
 sg13g2_and2_1 _20727_ (.A(net5981),
    .B(_04138_),
    .X(_00305_));
 sg13g2_nand2_1 _20728_ (.Y(_04139_),
    .A(\r_pwm_odd[6] ),
    .B(net6015));
 sg13g2_o21ai_1 _20729_ (.B1(_04092_),
    .Y(_04140_),
    .A1(_04061_),
    .A2(_04133_));
 sg13g2_nand3_1 _20730_ (.B(_04109_),
    .C(_04118_),
    .A(net5848),
    .Y(_04141_));
 sg13g2_nand2_2 _20731_ (.Y(_04142_),
    .A(net5897),
    .B(_03719_));
 sg13g2_nor3_1 _20732_ (.A(net5906),
    .B(_03718_),
    .C(_04040_),
    .Y(_04143_));
 sg13g2_a21oi_1 _20733_ (.A1(_03822_),
    .A2(_04143_),
    .Y(_04144_),
    .B1(net5891));
 sg13g2_nand2_1 _20734_ (.Y(_04145_),
    .A(_04030_),
    .B(_04144_));
 sg13g2_nor2_2 _20735_ (.A(_03716_),
    .B(_04048_),
    .Y(_04146_));
 sg13g2_nor2_1 _20736_ (.A(_04051_),
    .B(_04146_),
    .Y(_04147_));
 sg13g2_nor2_1 _20737_ (.A(net5908),
    .B(_04048_),
    .Y(_04148_));
 sg13g2_nand2_1 _20738_ (.Y(_04149_),
    .A(net5898),
    .B(_04049_));
 sg13g2_nand2_1 _20739_ (.Y(_04150_),
    .A(net5899),
    .B(_04146_));
 sg13g2_nand3b_1 _20740_ (.B(_04150_),
    .C(net5889),
    .Y(_04151_),
    .A_N(_04147_));
 sg13g2_nand3_1 _20741_ (.B(_04145_),
    .C(_04151_),
    .A(_04021_),
    .Y(_04152_));
 sg13g2_nand2_1 _20742_ (.Y(_04153_),
    .A(_04071_),
    .B(_04120_));
 sg13g2_nand3b_1 _20743_ (.B(_04153_),
    .C(net5889),
    .Y(_04154_),
    .A_N(_04147_));
 sg13g2_nand3_1 _20744_ (.B(net5920),
    .C(_03820_),
    .A(net5908),
    .Y(_04155_));
 sg13g2_nand2_1 _20745_ (.Y(_04156_),
    .A(net5905),
    .B(_04040_));
 sg13g2_nand4_1 _20746_ (.B(_04075_),
    .C(_04155_),
    .A(net5882),
    .Y(_04157_),
    .D(_04156_));
 sg13g2_nand3_1 _20747_ (.B(_04154_),
    .C(_04157_),
    .A(net5816),
    .Y(_04158_));
 sg13g2_nand2_1 _20748_ (.Y(_04159_),
    .A(net5897),
    .B(_04069_));
 sg13g2_o21ai_1 _20749_ (.B1(net5905),
    .Y(_04160_),
    .A1(_04026_),
    .A2(net5879));
 sg13g2_and2_1 _20750_ (.A(net5888),
    .B(_04160_),
    .X(_04161_));
 sg13g2_nand2_1 _20751_ (.Y(_04162_),
    .A(_04159_),
    .B(_04161_));
 sg13g2_nand2_1 _20752_ (.Y(_04163_),
    .A(_03830_),
    .B(net5845));
 sg13g2_o21ai_1 _20753_ (.B1(net5880),
    .Y(_04164_),
    .A1(_04051_),
    .A2(_04146_));
 sg13g2_nand2b_1 _20754_ (.Y(_04165_),
    .B(_04163_),
    .A_N(_04164_));
 sg13g2_nand3_1 _20755_ (.B(_04162_),
    .C(_04165_),
    .A(net5877),
    .Y(_04166_));
 sg13g2_nand4_1 _20756_ (.B(_04152_),
    .C(_04158_),
    .A(_04141_),
    .Y(_04167_),
    .D(_04166_));
 sg13g2_inv_1 _20757_ (.Y(_04168_),
    .A(_04167_));
 sg13g2_nand2_1 _20758_ (.Y(_04169_),
    .A(_04133_),
    .B(_04168_));
 sg13g2_nor2_1 _20759_ (.A(_04133_),
    .B(_04168_),
    .Y(_04170_));
 sg13g2_xnor2_1 _20760_ (.Y(_04171_),
    .A(_04133_),
    .B(_04167_));
 sg13g2_xnor2_1 _20761_ (.Y(_04172_),
    .A(_04140_),
    .B(_04171_));
 sg13g2_nand2b_1 _20762_ (.Y(_04173_),
    .B(_04172_),
    .A_N(_04139_));
 sg13g2_xnor2_1 _20763_ (.Y(_04174_),
    .A(_04139_),
    .B(_04172_));
 sg13g2_a21oi_1 _20764_ (.A1(_04099_),
    .A2(_04136_),
    .Y(_04175_),
    .B1(_04135_));
 sg13g2_nand2b_1 _20765_ (.Y(_04176_),
    .B(_04174_),
    .A_N(_04175_));
 sg13g2_xnor2_1 _20766_ (.Y(_04177_),
    .A(_04174_),
    .B(_04175_));
 sg13g2_and2_1 _20767_ (.A(net5982),
    .B(_04177_),
    .X(_00306_));
 sg13g2_and2_1 _20768_ (.A(_04173_),
    .B(_04176_),
    .X(_04178_));
 sg13g2_nand2_1 _20769_ (.Y(_04179_),
    .A(\r_pwm_odd[7] ),
    .B(net6015));
 sg13g2_or2_2 _20770_ (.X(_04180_),
    .B(_03822_),
    .A(net5925));
 sg13g2_a21o_1 _20771_ (.A2(_04180_),
    .A1(net5893),
    .B1(net5899),
    .X(_04181_));
 sg13g2_a21oi_1 _20772_ (.A1(net5903),
    .A2(_03823_),
    .Y(_04182_),
    .B1(net5880));
 sg13g2_nand2_1 _20773_ (.Y(_04183_),
    .A(_04181_),
    .B(_04182_));
 sg13g2_a21oi_2 _20774_ (.B1(net5905),
    .Y(_04184_),
    .A2(_03820_),
    .A1(net5894));
 sg13g2_nand2_1 _20775_ (.Y(_04185_),
    .A(net5897),
    .B(_03821_));
 sg13g2_a21oi_1 _20776_ (.A1(net5904),
    .A2(_04068_),
    .Y(_04186_),
    .B1(_04184_));
 sg13g2_nand2_1 _20777_ (.Y(_04187_),
    .A(net5899),
    .B(net5880));
 sg13g2_inv_1 _20778_ (.Y(_04188_),
    .A(_04187_));
 sg13g2_nand2_1 _20779_ (.Y(_04189_),
    .A(net5882),
    .B(_04186_));
 sg13g2_nand2_1 _20780_ (.Y(_04190_),
    .A(_04183_),
    .B(_04189_));
 sg13g2_a22oi_1 _20781_ (.Y(_04191_),
    .B1(_04190_),
    .B2(net5816),
    .A2(net5848),
    .A1(_03823_));
 sg13g2_nor2_1 _20782_ (.A(net5889),
    .B(_04181_),
    .Y(_04192_));
 sg13g2_nor2_1 _20783_ (.A(_04069_),
    .B(_04101_),
    .Y(_04193_));
 sg13g2_a21o_1 _20784_ (.A2(_04193_),
    .A1(_04188_),
    .B1(_04192_),
    .X(_04194_));
 sg13g2_nand3_1 _20785_ (.B(_03820_),
    .C(net5847),
    .A(_03618_),
    .Y(_04195_));
 sg13g2_nand2_2 _20786_ (.Y(_04196_),
    .A(_03713_),
    .B(_04033_));
 sg13g2_nand2_1 _20787_ (.Y(_04197_),
    .A(_04078_),
    .B(_04196_));
 sg13g2_o21ai_1 _20788_ (.B1(_04195_),
    .Y(_04198_),
    .A1(_04101_),
    .A2(_04197_));
 sg13g2_o21ai_1 _20789_ (.B1(net5877),
    .Y(_04199_),
    .A1(_04194_),
    .A2(_04198_));
 sg13g2_nor2_1 _20790_ (.A(_04070_),
    .B(_04142_),
    .Y(_04200_));
 sg13g2_nand2b_1 _20791_ (.Y(_04201_),
    .B(_04071_),
    .A_N(_04142_));
 sg13g2_nand3b_1 _20792_ (.B(net5893),
    .C(net5904),
    .Y(_04202_),
    .A_N(_03720_));
 sg13g2_and2_1 _20793_ (.A(net5897),
    .B(net5893),
    .X(_04203_));
 sg13g2_nand2_1 _20794_ (.Y(_04204_),
    .A(_04180_),
    .B(_04203_));
 sg13g2_a21oi_1 _20795_ (.A1(_04180_),
    .A2(_04203_),
    .Y(_04205_),
    .B1(net5888));
 sg13g2_a21oi_1 _20796_ (.A1(_04202_),
    .A2(_04204_),
    .Y(_04206_),
    .B1(net5889));
 sg13g2_a21oi_1 _20797_ (.A1(_04181_),
    .A2(_04201_),
    .Y(_04207_),
    .B1(net5880));
 sg13g2_o21ai_1 _20798_ (.B1(_04021_),
    .Y(_04208_),
    .A1(_04206_),
    .A2(_04207_));
 sg13g2_nand3_1 _20799_ (.B(_04199_),
    .C(_04208_),
    .A(_04191_),
    .Y(_04209_));
 sg13g2_xnor2_1 _20800_ (.Y(_04210_),
    .A(_04168_),
    .B(_04209_));
 sg13g2_o21ai_1 _20801_ (.B1(_04169_),
    .Y(_04211_),
    .A1(_04140_),
    .A2(_04170_));
 sg13g2_nand2_1 _20802_ (.Y(_04212_),
    .A(_04210_),
    .B(_04211_));
 sg13g2_xnor2_1 _20803_ (.Y(_04213_),
    .A(_04210_),
    .B(_04211_));
 sg13g2_nor2_1 _20804_ (.A(_04179_),
    .B(_04213_),
    .Y(_04214_));
 sg13g2_xor2_1 _20805_ (.B(_04213_),
    .A(_04179_),
    .X(_04215_));
 sg13g2_nor2b_1 _20806_ (.A(_04178_),
    .B_N(_04215_),
    .Y(_04216_));
 sg13g2_xnor2_1 _20807_ (.Y(_04217_),
    .A(_04178_),
    .B(_04215_));
 sg13g2_and2_1 _20808_ (.A(net5983),
    .B(_04217_),
    .X(_00307_));
 sg13g2_nor2_2 _20809_ (.A(_04214_),
    .B(_04216_),
    .Y(_04218_));
 sg13g2_nor2_1 _20810_ (.A(_03818_),
    .B(_04196_),
    .Y(_04219_));
 sg13g2_nor3_1 _20811_ (.A(net5882),
    .B(_04101_),
    .C(_04184_),
    .Y(_04220_));
 sg13g2_o21ai_1 _20812_ (.B1(net5816),
    .Y(_04221_),
    .A1(_04219_),
    .A2(_04220_));
 sg13g2_o21ai_1 _20813_ (.B1(net6085),
    .Y(_04222_),
    .A1(_03434_),
    .A2(net5924));
 sg13g2_a21oi_1 _20814_ (.A1(_03713_),
    .A2(_04222_),
    .Y(_04223_),
    .B1(_03618_));
 sg13g2_nand2_1 _20815_ (.Y(_04224_),
    .A(net5882),
    .B(_04223_));
 sg13g2_o21ai_1 _20816_ (.B1(_04185_),
    .Y(_04225_),
    .A1(net5897),
    .A2(_04033_));
 sg13g2_a21oi_1 _20817_ (.A1(net5888),
    .A2(_04225_),
    .Y(_04226_),
    .B1(_04020_));
 sg13g2_nor2_1 _20818_ (.A(_04079_),
    .B(_04196_),
    .Y(_04227_));
 sg13g2_nor2_1 _20819_ (.A(net5888),
    .B(_04225_),
    .Y(_04228_));
 sg13g2_o21ai_1 _20820_ (.B1(net5877),
    .Y(_04229_),
    .A1(_04227_),
    .A2(_04228_));
 sg13g2_a22oi_1 _20821_ (.Y(_04230_),
    .B1(_04224_),
    .B2(_04226_),
    .A2(net5848),
    .A1(_03719_));
 sg13g2_nand3_1 _20822_ (.B(_04229_),
    .C(_04230_),
    .A(_04221_),
    .Y(_04231_));
 sg13g2_xor2_1 _20823_ (.B(_04231_),
    .A(_04209_),
    .X(_04232_));
 sg13g2_o21ai_1 _20824_ (.B1(_04212_),
    .Y(_04233_),
    .A1(_04167_),
    .A2(_04209_));
 sg13g2_nand2_1 _20825_ (.Y(_04234_),
    .A(_04232_),
    .B(_04233_));
 sg13g2_xor2_1 _20826_ (.B(_04233_),
    .A(_04232_),
    .X(_04235_));
 sg13g2_nand2b_1 _20827_ (.Y(_04236_),
    .B(_04218_),
    .A_N(_04235_));
 sg13g2_o21ai_1 _20828_ (.B1(_04235_),
    .Y(_04237_),
    .A1(_04214_),
    .A2(_04216_));
 sg13g2_and3_1 _20829_ (.X(_00308_),
    .A(net5983),
    .B(_04236_),
    .C(_04237_));
 sg13g2_a21oi_2 _20830_ (.B1(_04231_),
    .Y(_04238_),
    .A2(_04212_),
    .A1(_04209_));
 sg13g2_a21o_1 _20831_ (.A2(_04234_),
    .A1(_04231_),
    .B1(_04238_),
    .X(_04239_));
 sg13g2_and2_1 _20832_ (.A(_04237_),
    .B(_04239_),
    .X(_04240_));
 sg13g2_nor2_1 _20833_ (.A(_04237_),
    .B(_04239_),
    .Y(_04241_));
 sg13g2_nor3_2 _20834_ (.A(net5986),
    .B(_04240_),
    .C(_04241_),
    .Y(_00309_));
 sg13g2_nor2_1 _20835_ (.A(_04238_),
    .B(_04241_),
    .Y(_04242_));
 sg13g2_nor2_2 _20836_ (.A(net5986),
    .B(_04242_),
    .Y(_00310_));
 sg13g2_and3_1 _20837_ (.X(_00311_),
    .A(net2991),
    .B(net5982),
    .C(net6019));
 sg13g2_nor2_1 _20838_ (.A(_03714_),
    .B(_03723_),
    .Y(_04243_));
 sg13g2_or2_1 _20839_ (.X(_04244_),
    .B(_03723_),
    .A(net5896));
 sg13g2_a21o_1 _20840_ (.A2(_04244_),
    .A1(_04104_),
    .B1(net5900),
    .X(_04245_));
 sg13g2_nand2_2 _20841_ (.Y(_04246_),
    .A(net5896),
    .B(_04039_));
 sg13g2_o21ai_1 _20842_ (.B1(net5908),
    .Y(_04247_),
    .A1(_03713_),
    .A2(_04118_));
 sg13g2_a21oi_1 _20843_ (.A1(_03831_),
    .A2(_04247_),
    .Y(_04248_),
    .B1(net5886));
 sg13g2_a21oi_1 _20844_ (.A1(_03826_),
    .A2(_04245_),
    .Y(_04249_),
    .B1(_04057_));
 sg13g2_nand2b_1 _20845_ (.Y(_04250_),
    .B(_04249_),
    .A_N(_04248_));
 sg13g2_a21o_1 _20846_ (.A2(_04196_),
    .A1(_04035_),
    .B1(net5906),
    .X(_04251_));
 sg13g2_nand2_1 _20847_ (.Y(_04252_),
    .A(net5907),
    .B(_04058_));
 sg13g2_a21oi_1 _20848_ (.A1(_04251_),
    .A2(_04252_),
    .Y(_04253_),
    .B1(_04055_));
 sg13g2_xnor2_1 _20849_ (.Y(_04254_),
    .A(net5901),
    .B(net5891));
 sg13g2_nand3_1 _20850_ (.B(_04244_),
    .C(_04254_),
    .A(net5845),
    .Y(_04255_));
 sg13g2_nor2_1 _20851_ (.A(_03725_),
    .B(_04254_),
    .Y(_04256_));
 sg13g2_nor2_1 _20852_ (.A(_04024_),
    .B(_04256_),
    .Y(_04257_));
 sg13g2_a21oi_1 _20853_ (.A1(_04255_),
    .A2(_04257_),
    .Y(_04258_),
    .B1(_04253_));
 sg13g2_mux2_1 _20854_ (.A0(net5921),
    .A1(net5894),
    .S(net5902),
    .X(_04259_));
 sg13g2_a21o_1 _20855_ (.A2(_04246_),
    .A1(_04086_),
    .B1(_04259_),
    .X(_04260_));
 sg13g2_o21ai_1 _20856_ (.B1(net5902),
    .Y(_04261_),
    .A1(_03717_),
    .A2(_04048_));
 sg13g2_nand2_1 _20857_ (.Y(_04262_),
    .A(_03829_),
    .B(_04261_));
 sg13g2_a21oi_1 _20858_ (.A1(net5884),
    .A2(_04260_),
    .Y(_04263_),
    .B1(_04020_));
 sg13g2_o21ai_1 _20859_ (.B1(_04263_),
    .Y(_04264_),
    .A1(net5885),
    .A2(_04262_));
 sg13g2_nand4_1 _20860_ (.B(_04250_),
    .C(_04258_),
    .A(_04046_),
    .Y(_04265_),
    .D(_04264_));
 sg13g2_nand2b_1 _20861_ (.Y(_04266_),
    .B(net6019),
    .A_N(net7512));
 sg13g2_nand2_1 _20862_ (.Y(_04267_),
    .A(_04265_),
    .B(_04266_));
 sg13g2_inv_1 _20863_ (.Y(_04268_),
    .A(_04267_));
 sg13g2_nor2_2 _20864_ (.A(_04265_),
    .B(_04266_),
    .Y(_04269_));
 sg13g2_nor3_1 _20865_ (.A(net5987),
    .B(_04268_),
    .C(_04269_),
    .Y(_00312_));
 sg13g2_nand2_1 _20866_ (.Y(_04270_),
    .A(\g_pwm_odd[4] ),
    .B(net6019));
 sg13g2_a21o_1 _20867_ (.A2(_04155_),
    .A1(_04088_),
    .B1(net5883),
    .X(_04271_));
 sg13g2_nand3_1 _20868_ (.B(_04088_),
    .C(_04108_),
    .A(net5883),
    .Y(_04272_));
 sg13g2_nand3_1 _20869_ (.B(_04271_),
    .C(_04272_),
    .A(_04019_),
    .Y(_04273_));
 sg13g2_o21ai_1 _20870_ (.B1(net5892),
    .Y(_04274_),
    .A1(_04113_),
    .A2(_04114_));
 sg13g2_nor2_1 _20871_ (.A(net5895),
    .B(net5892),
    .Y(_04275_));
 sg13g2_o21ai_1 _20872_ (.B1(_04275_),
    .Y(_04276_),
    .A1(_03713_),
    .A2(_04222_));
 sg13g2_a21oi_1 _20873_ (.A1(_04036_),
    .A2(net5847),
    .Y(_04277_),
    .B1(net5849));
 sg13g2_nand3_1 _20874_ (.B(_04276_),
    .C(_04277_),
    .A(_04274_),
    .Y(_04278_));
 sg13g2_nand3_1 _20875_ (.B(_04273_),
    .C(_04278_),
    .A(_03924_),
    .Y(_04279_));
 sg13g2_a21oi_1 _20876_ (.A1(_04203_),
    .A2(_04246_),
    .Y(_04280_),
    .B1(net5892));
 sg13g2_nand2b_1 _20877_ (.Y(_04281_),
    .B(net5893),
    .A_N(_04247_));
 sg13g2_a21oi_1 _20878_ (.A1(_04025_),
    .A2(_04203_),
    .Y(_04282_),
    .B1(net5884));
 sg13g2_a22oi_1 _20879_ (.Y(_04283_),
    .B1(_04281_),
    .B2(_04282_),
    .A2(_04280_),
    .A1(_04108_));
 sg13g2_a221oi_1 _20880_ (.B2(_04069_),
    .C1(net5883),
    .B1(_04148_),
    .A1(_04050_),
    .Y(_04284_),
    .A2(net5846));
 sg13g2_nor3_1 _20881_ (.A(_04044_),
    .B(_04076_),
    .C(_04284_),
    .Y(_04285_));
 sg13g2_a21oi_2 _20882_ (.B1(_04285_),
    .Y(_04286_),
    .A2(_04283_),
    .A1(net5816));
 sg13g2_and2_1 _20883_ (.A(_04279_),
    .B(_04286_),
    .X(_04287_));
 sg13g2_nand2_1 _20884_ (.Y(_04288_),
    .A(_04279_),
    .B(_04286_));
 sg13g2_nand2_2 _20885_ (.Y(_04289_),
    .A(_04265_),
    .B(_04287_));
 sg13g2_nand2b_1 _20886_ (.Y(_04290_),
    .B(_04288_),
    .A_N(_04265_));
 sg13g2_nand2_1 _20887_ (.Y(_04291_),
    .A(_04289_),
    .B(_04290_));
 sg13g2_a21oi_1 _20888_ (.A1(_04289_),
    .A2(_04290_),
    .Y(_04292_),
    .B1(_04270_));
 sg13g2_nand3_1 _20889_ (.B(_04289_),
    .C(_04290_),
    .A(_04270_),
    .Y(_04293_));
 sg13g2_nand2b_1 _20890_ (.Y(_04294_),
    .B(_04293_),
    .A_N(_04292_));
 sg13g2_xnor2_1 _20891_ (.Y(_04295_),
    .A(_04269_),
    .B(_04294_));
 sg13g2_and2_1 _20892_ (.A(net5982),
    .B(_04295_),
    .X(_00313_));
 sg13g2_nand2_2 _20893_ (.Y(_04296_),
    .A(\g_pwm_odd[5] ),
    .B(net6018));
 sg13g2_o21ai_1 _20894_ (.B1(_04115_),
    .Y(_04297_),
    .A1(net5900),
    .A2(_04104_));
 sg13g2_nand3_1 _20895_ (.B(_04025_),
    .C(_04121_),
    .A(net5891),
    .Y(_04298_));
 sg13g2_a21oi_1 _20896_ (.A1(_04297_),
    .A2(_04298_),
    .Y(_04299_),
    .B1(_04057_));
 sg13g2_a221oi_1 _20897_ (.B2(_03820_),
    .C1(net5902),
    .B1(net5895),
    .A1(net5921),
    .Y(_04300_),
    .A2(net5919));
 sg13g2_nand2b_1 _20898_ (.Y(_04301_),
    .B(_04282_),
    .A_N(_04300_));
 sg13g2_a21oi_1 _20899_ (.A1(_04129_),
    .A2(_04301_),
    .Y(_04302_),
    .B1(_04044_));
 sg13g2_a22oi_1 _20900_ (.Y(_04303_),
    .B1(_04184_),
    .B2(_04025_),
    .A2(_04118_),
    .A1(net5908));
 sg13g2_nor3_1 _20901_ (.A(net5892),
    .B(_04102_),
    .C(_04222_),
    .Y(_04304_));
 sg13g2_o21ai_1 _20902_ (.B1(_04021_),
    .Y(_04305_),
    .A1(net5883),
    .A2(_04303_));
 sg13g2_nor2_1 _20903_ (.A(_04304_),
    .B(_04305_),
    .Y(_04306_));
 sg13g2_and2_1 _20904_ (.A(_04034_),
    .B(_04102_),
    .X(_04307_));
 sg13g2_o21ai_1 _20905_ (.B1(net5816),
    .Y(_04308_),
    .A1(_04254_),
    .A2(_04307_));
 sg13g2_a21oi_1 _20906_ (.A1(_04082_),
    .A2(_04254_),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_nor4_2 _20907_ (.A(_04299_),
    .B(_04302_),
    .C(_04306_),
    .Y(_04310_),
    .D(_04309_));
 sg13g2_xnor2_1 _20908_ (.Y(_04311_),
    .A(_04289_),
    .B(_04310_));
 sg13g2_xnor2_1 _20909_ (.Y(_04312_),
    .A(_04296_),
    .B(_04311_));
 sg13g2_a21o_1 _20910_ (.A2(_04293_),
    .A1(_04269_),
    .B1(_04292_),
    .X(_04313_));
 sg13g2_nand2b_1 _20911_ (.Y(_04314_),
    .B(_04313_),
    .A_N(_04312_));
 sg13g2_xor2_1 _20912_ (.B(_04313_),
    .A(_04312_),
    .X(_04315_));
 sg13g2_nor2_1 _20913_ (.A(net5987),
    .B(_04315_),
    .Y(_00314_));
 sg13g2_nand2_2 _20914_ (.Y(_04316_),
    .A(\g_pwm_odd[6] ),
    .B(net6018));
 sg13g2_a21o_1 _20915_ (.A2(_04246_),
    .A1(net5846),
    .B1(net5906),
    .X(_04317_));
 sg13g2_nand3_1 _20916_ (.B(_04105_),
    .C(_04317_),
    .A(net5881),
    .Y(_04318_));
 sg13g2_nand2b_1 _20917_ (.Y(_04319_),
    .B(net5846),
    .A_N(_04247_));
 sg13g2_a21oi_1 _20918_ (.A1(_04103_),
    .A2(_04319_),
    .Y(_04320_),
    .B1(net5881));
 sg13g2_nand3b_1 _20919_ (.B(net5816),
    .C(_04318_),
    .Y(_04321_),
    .A_N(_04320_));
 sg13g2_or2_1 _20920_ (.X(_04322_),
    .B(_04039_),
    .A(_04026_));
 sg13g2_nand2_1 _20921_ (.Y(_04323_),
    .A(net5905),
    .B(_04322_));
 sg13g2_nand3_1 _20922_ (.B(_04150_),
    .C(_04323_),
    .A(net5889),
    .Y(_04324_));
 sg13g2_nand3_1 _20923_ (.B(_04145_),
    .C(_04324_),
    .A(net5848),
    .Y(_04325_));
 sg13g2_nand3_1 _20924_ (.B(_04078_),
    .C(net5845),
    .A(_04049_),
    .Y(_04326_));
 sg13g2_a22oi_1 _20925_ (.Y(_04327_),
    .B1(_04322_),
    .B2(net5881),
    .A2(_04146_),
    .A1(net5847));
 sg13g2_a21o_1 _20926_ (.A2(_04327_),
    .A1(_04326_),
    .B1(_04020_),
    .X(_04328_));
 sg13g2_a21oi_1 _20927_ (.A1(_03719_),
    .A2(_04028_),
    .Y(_04329_),
    .B1(net5882));
 sg13g2_nand2_1 _20928_ (.Y(_04330_),
    .A(_04103_),
    .B(_04329_));
 sg13g2_nand3_1 _20929_ (.B(_04165_),
    .C(_04330_),
    .A(net5877),
    .Y(_04331_));
 sg13g2_nand4_1 _20930_ (.B(_04325_),
    .C(_04328_),
    .A(_04321_),
    .Y(_04332_),
    .D(_04331_));
 sg13g2_nand2b_1 _20931_ (.Y(_04333_),
    .B(_04287_),
    .A_N(_04310_));
 sg13g2_o21ai_1 _20932_ (.B1(_04310_),
    .Y(_04334_),
    .A1(_04265_),
    .A2(_04288_));
 sg13g2_inv_1 _20933_ (.Y(_04335_),
    .A(_04334_));
 sg13g2_nand2_1 _20934_ (.Y(_04336_),
    .A(_04333_),
    .B(_04334_));
 sg13g2_xor2_1 _20935_ (.B(_04336_),
    .A(_04332_),
    .X(_04337_));
 sg13g2_inv_1 _20936_ (.Y(_04338_),
    .A(_04337_));
 sg13g2_nor2_1 _20937_ (.A(_04316_),
    .B(_04338_),
    .Y(_04339_));
 sg13g2_xnor2_1 _20938_ (.Y(_04340_),
    .A(_04316_),
    .B(_04337_));
 sg13g2_o21ai_1 _20939_ (.B1(_04314_),
    .Y(_04341_),
    .A1(_04296_),
    .A2(_04311_));
 sg13g2_xnor2_1 _20940_ (.Y(_04342_),
    .A(_04340_),
    .B(_04341_));
 sg13g2_nor2_1 _20941_ (.A(net5988),
    .B(_04342_),
    .Y(_00315_));
 sg13g2_nand2_2 _20942_ (.Y(_04343_),
    .A(\g_pwm_odd[7] ),
    .B(net6014));
 sg13g2_nand2_2 _20943_ (.Y(_04344_),
    .A(net5882),
    .B(net5849));
 sg13g2_inv_1 _20944_ (.Y(_04345_),
    .A(_04344_));
 sg13g2_o21ai_1 _20945_ (.B1(_03721_),
    .Y(_04346_),
    .A1(_03434_),
    .A2(_03713_));
 sg13g2_a21oi_2 _20946_ (.B1(net5882),
    .Y(_04347_),
    .A2(_04346_),
    .A1(_04118_));
 sg13g2_nor3_1 _20947_ (.A(_04018_),
    .B(_04194_),
    .C(_04347_),
    .Y(_04348_));
 sg13g2_or2_1 _20948_ (.X(_04349_),
    .B(_03823_),
    .A(_03716_));
 sg13g2_nor2_1 _20949_ (.A(net5918),
    .B(_04348_),
    .Y(_04350_));
 sg13g2_o21ai_1 _20950_ (.B1(_04350_),
    .Y(_04351_),
    .A1(net5849),
    .A2(_04349_));
 sg13g2_nor3_1 _20951_ (.A(_04069_),
    .B(net5847),
    .C(_04101_),
    .Y(_04352_));
 sg13g2_nor3_1 _20952_ (.A(net5880),
    .B(_04051_),
    .C(_04070_),
    .Y(_04353_));
 sg13g2_o21ai_1 _20953_ (.B1(_04021_),
    .Y(_04354_),
    .A1(_04352_),
    .A2(_04353_));
 sg13g2_a221oi_1 _20954_ (.B2(net5889),
    .C1(_04206_),
    .B1(_04200_),
    .A1(net5847),
    .Y(_04355_),
    .A2(_04193_));
 sg13g2_nand2b_1 _20955_ (.Y(_04356_),
    .B(net5848),
    .A_N(_04355_));
 sg13g2_nand3_1 _20956_ (.B(_04354_),
    .C(_04356_),
    .A(_04351_),
    .Y(_04357_));
 sg13g2_xor2_1 _20957_ (.B(_04357_),
    .A(_04332_),
    .X(_04358_));
 sg13g2_o21ai_1 _20958_ (.B1(_04333_),
    .Y(_04359_),
    .A1(_04332_),
    .A2(_04335_));
 sg13g2_nand2_1 _20959_ (.Y(_04360_),
    .A(_04358_),
    .B(_04359_));
 sg13g2_xnor2_1 _20960_ (.Y(_04361_),
    .A(_04358_),
    .B(_04359_));
 sg13g2_xor2_1 _20961_ (.B(_04361_),
    .A(_04343_),
    .X(_04362_));
 sg13g2_a21oi_2 _20962_ (.B1(_04339_),
    .Y(_04363_),
    .A2(_04341_),
    .A1(_04340_));
 sg13g2_nand2b_1 _20963_ (.Y(_04364_),
    .B(_04362_),
    .A_N(_04363_));
 sg13g2_xor2_1 _20964_ (.B(_04363_),
    .A(_04362_),
    .X(_04365_));
 sg13g2_nor2_1 _20965_ (.A(net5988),
    .B(_04365_),
    .Y(_00316_));
 sg13g2_o21ai_1 _20966_ (.B1(_04364_),
    .Y(_04366_),
    .A1(_04343_),
    .A2(_04361_));
 sg13g2_o21ai_1 _20967_ (.B1(_04360_),
    .Y(_04367_),
    .A1(_04332_),
    .A2(_04357_));
 sg13g2_nor2_1 _20968_ (.A(_04223_),
    .B(_04344_),
    .Y(_04368_));
 sg13g2_o21ai_1 _20969_ (.B1(net5918),
    .Y(_04369_),
    .A1(_03821_),
    .A2(_04345_));
 sg13g2_nor2_1 _20970_ (.A(_04368_),
    .B(_04369_),
    .Y(_04370_));
 sg13g2_o21ai_1 _20971_ (.B1(net5877),
    .Y(_04371_),
    .A1(net5920),
    .A2(net5882));
 sg13g2_a21oi_1 _20972_ (.A1(net5816),
    .A2(_04101_),
    .Y(_04372_),
    .B1(_04370_));
 sg13g2_o21ai_1 _20973_ (.B1(_04372_),
    .Y(_04373_),
    .A1(_04228_),
    .A2(_04371_));
 sg13g2_nand2b_1 _20974_ (.Y(_04374_),
    .B(_04373_),
    .A_N(_04357_));
 sg13g2_xor2_1 _20975_ (.B(_04373_),
    .A(_04357_),
    .X(_04375_));
 sg13g2_nand2b_1 _20976_ (.Y(_04376_),
    .B(_04367_),
    .A_N(_04375_));
 sg13g2_xnor2_1 _20977_ (.Y(_04377_),
    .A(_04367_),
    .B(_04375_));
 sg13g2_o21ai_1 _20978_ (.B1(net5983),
    .Y(_04378_),
    .A1(_04366_),
    .A2(_04377_));
 sg13g2_a21oi_1 _20979_ (.A1(_04366_),
    .A2(_04377_),
    .Y(_00317_),
    .B1(_04378_));
 sg13g2_nand2_1 _20980_ (.Y(_04379_),
    .A(_04374_),
    .B(_04376_));
 sg13g2_nand2_1 _20981_ (.Y(_04380_),
    .A(_04373_),
    .B(_04379_));
 sg13g2_xor2_1 _20982_ (.B(_04379_),
    .A(_04373_),
    .X(_04381_));
 sg13g2_a21o_1 _20983_ (.A2(_04377_),
    .A1(_04366_),
    .B1(_04381_),
    .X(_04382_));
 sg13g2_nand3_1 _20984_ (.B(_04377_),
    .C(_04381_),
    .A(_04366_),
    .Y(_04383_));
 sg13g2_and3_2 _20985_ (.X(_00318_),
    .A(net5980),
    .B(_04382_),
    .C(_04383_));
 sg13g2_a21oi_2 _20986_ (.B1(net5984),
    .Y(_00319_),
    .A2(_04383_),
    .A1(_04380_));
 sg13g2_and2_1 _20987_ (.A(net7576),
    .B(net6014),
    .X(_04384_));
 sg13g2_nor3_2 _20988_ (.A(net5906),
    .B(_04055_),
    .C(_04180_),
    .Y(_04385_));
 sg13g2_nand2_1 _20989_ (.Y(_04386_),
    .A(\b_pwm_odd[1] ),
    .B(net6018));
 sg13g2_nand2_1 _20990_ (.Y(_04387_),
    .A(_04385_),
    .B(_04386_));
 sg13g2_xor2_1 _20991_ (.B(_04387_),
    .A(_04384_),
    .X(_04388_));
 sg13g2_nor2_1 _20992_ (.A(net5987),
    .B(_04388_),
    .Y(_00320_));
 sg13g2_a22oi_1 _20993_ (.Y(_04389_),
    .B1(_04120_),
    .B2(_04027_),
    .A2(net5845),
    .A1(net5905));
 sg13g2_a22oi_1 _20994_ (.Y(_04390_),
    .B1(_04107_),
    .B2(net5885),
    .A2(_04038_),
    .A1(_03830_));
 sg13g2_o21ai_1 _20995_ (.B1(_04390_),
    .Y(_04391_),
    .A1(net5885),
    .A2(_04389_));
 sg13g2_nand2_1 _20996_ (.Y(_04392_),
    .A(_03826_),
    .B(_04252_));
 sg13g2_nand3_1 _20997_ (.B(_04102_),
    .C(_04196_),
    .A(_04078_),
    .Y(_04393_));
 sg13g2_o21ai_1 _20998_ (.B1(net5847),
    .Y(_04394_),
    .A1(_03718_),
    .A2(_04036_));
 sg13g2_nand4_1 _20999_ (.B(_04392_),
    .C(_04393_),
    .A(_04021_),
    .Y(_04395_),
    .D(_04394_));
 sg13g2_a21oi_1 _21000_ (.A1(net5907),
    .A2(_04244_),
    .Y(_04396_),
    .B1(net5890));
 sg13g2_a22oi_1 _21001_ (.Y(_04397_),
    .B1(_04243_),
    .B2(net5900),
    .A2(net5876),
    .A1(_04049_));
 sg13g2_a221oi_1 _21002_ (.B2(net5890),
    .C1(_04024_),
    .B1(_04397_),
    .A1(_03831_),
    .Y(_04398_),
    .A2(_04396_));
 sg13g2_nor4_1 _21003_ (.A(net5906),
    .B(_03718_),
    .C(net5891),
    .D(_04040_),
    .Y(_04399_));
 sg13g2_a21o_1 _21004_ (.A2(_04070_),
    .A1(_03817_),
    .B1(_04399_),
    .X(_04400_));
 sg13g2_a21o_1 _21005_ (.A2(_04251_),
    .A1(_04031_),
    .B1(_04400_),
    .X(_04401_));
 sg13g2_a221oi_1 _21006_ (.B2(net5848),
    .C1(_04398_),
    .B1(_04401_),
    .A1(net5878),
    .Y(_04402_),
    .A2(_04391_));
 sg13g2_nand2_2 _21007_ (.Y(_04403_),
    .A(_04395_),
    .B(_04402_));
 sg13g2_and2_1 _21008_ (.A(\b_pwm_odd[3] ),
    .B(net6014),
    .X(_04404_));
 sg13g2_nor2b_1 _21009_ (.A(_04403_),
    .B_N(_04404_),
    .Y(_04405_));
 sg13g2_a21o_1 _21010_ (.A2(_04402_),
    .A1(_04395_),
    .B1(_04404_),
    .X(_04406_));
 sg13g2_xnor2_1 _21011_ (.Y(_04407_),
    .A(_04403_),
    .B(_04404_));
 sg13g2_o21ai_1 _21012_ (.B1(net6014),
    .Y(_04408_),
    .A1(\b_pwm_odd[2] ),
    .A2(\b_pwm_odd[1] ));
 sg13g2_nand2b_1 _21013_ (.Y(_04409_),
    .B(_04385_),
    .A_N(_04408_));
 sg13g2_inv_1 _21014_ (.Y(_04410_),
    .A(_04409_));
 sg13g2_xnor2_1 _21015_ (.Y(_04411_),
    .A(_04407_),
    .B(_04410_));
 sg13g2_nor2_1 _21016_ (.A(net5985),
    .B(_04411_),
    .Y(_00321_));
 sg13g2_nand2_1 _21017_ (.Y(_04412_),
    .A(\b_pwm_odd[4] ),
    .B(net6013));
 sg13g2_a221oi_1 _21018_ (.B2(net5846),
    .C1(net5892),
    .B1(net5876),
    .A1(net5902),
    .Y(_04413_),
    .A2(_04036_));
 sg13g2_nand2_1 _21019_ (.Y(_04414_),
    .A(net5908),
    .B(_04080_));
 sg13g2_a221oi_1 _21020_ (.B2(_04180_),
    .C1(net5883),
    .B1(_04148_),
    .A1(net5908),
    .Y(_04415_),
    .A2(_04080_));
 sg13g2_o21ai_1 _21021_ (.B1(_04018_),
    .Y(_04416_),
    .A1(_04413_),
    .A2(_04415_));
 sg13g2_nand2b_1 _21022_ (.Y(_04417_),
    .B(_04120_),
    .A_N(_03724_));
 sg13g2_a21oi_1 _21023_ (.A1(net5847),
    .A2(_04082_),
    .Y(_04418_),
    .B1(_04053_));
 sg13g2_o21ai_1 _21024_ (.B1(_04156_),
    .Y(_04419_),
    .A1(_04033_),
    .A2(_04142_));
 sg13g2_a221oi_1 _21025_ (.B2(_04345_),
    .C1(_03923_),
    .B1(_04419_),
    .A1(_04417_),
    .Y(_04420_),
    .A2(_04418_));
 sg13g2_nand2_1 _21026_ (.Y(_04421_),
    .A(net5902),
    .B(_04070_));
 sg13g2_a221oi_1 _21027_ (.B2(_04072_),
    .C1(net5849),
    .B1(_04421_),
    .A1(_04280_),
    .Y(_04422_),
    .A2(_04414_));
 sg13g2_a21oi_1 _21028_ (.A1(_04051_),
    .A2(_04075_),
    .Y(_04423_),
    .B1(_04344_));
 sg13g2_o21ai_1 _21029_ (.B1(_04180_),
    .Y(_04424_),
    .A1(_04028_),
    .A2(_04067_));
 sg13g2_nor2_1 _21030_ (.A(_04053_),
    .B(_04424_),
    .Y(_04425_));
 sg13g2_nor4_1 _21031_ (.A(net5918),
    .B(_04422_),
    .C(_04423_),
    .D(_04425_),
    .Y(_04426_));
 sg13g2_a21oi_2 _21032_ (.B1(_04426_),
    .Y(_04427_),
    .A2(_04420_),
    .A1(_04416_));
 sg13g2_a21oi_1 _21033_ (.A1(_04395_),
    .A2(_04402_),
    .Y(_04428_),
    .B1(_04427_));
 sg13g2_xnor2_1 _21034_ (.Y(_04429_),
    .A(_04403_),
    .B(_04427_));
 sg13g2_xor2_1 _21035_ (.B(_04427_),
    .A(_04403_),
    .X(_04430_));
 sg13g2_nor2_1 _21036_ (.A(_04412_),
    .B(_04429_),
    .Y(_04431_));
 sg13g2_nand2_1 _21037_ (.Y(_04432_),
    .A(_04412_),
    .B(_04429_));
 sg13g2_nand2b_1 _21038_ (.Y(_04433_),
    .B(_04432_),
    .A_N(_04431_));
 sg13g2_a21o_1 _21039_ (.A2(_04410_),
    .A1(_04406_),
    .B1(_04405_),
    .X(_04434_));
 sg13g2_xnor2_1 _21040_ (.Y(_04435_),
    .A(_04433_),
    .B(_04434_));
 sg13g2_and2_1 _21041_ (.A(net5980),
    .B(_04435_),
    .X(_00322_));
 sg13g2_nand2_2 _21042_ (.Y(_04436_),
    .A(\b_pwm_odd[5] ),
    .B(net6013));
 sg13g2_nand2_1 _21043_ (.Y(_04437_),
    .A(net5907),
    .B(_04131_));
 sg13g2_nand3_1 _21044_ (.B(_04081_),
    .C(_04196_),
    .A(_04035_),
    .Y(_04438_));
 sg13g2_and2_1 _21045_ (.A(_03822_),
    .B(net5846),
    .X(_04439_));
 sg13g2_a22oi_1 _21046_ (.Y(_04440_),
    .B1(_04439_),
    .B2(_04078_),
    .A2(_04437_),
    .A1(_04115_));
 sg13g2_a21oi_1 _21047_ (.A1(_04438_),
    .A2(_04440_),
    .Y(_04441_),
    .B1(_04020_));
 sg13g2_a21oi_1 _21048_ (.A1(_04049_),
    .A2(net5845),
    .Y(_04442_),
    .B1(_03818_));
 sg13g2_a21oi_1 _21049_ (.A1(_04029_),
    .A2(net5846),
    .Y(_04443_),
    .B1(_04125_));
 sg13g2_and2_1 _21050_ (.A(net5885),
    .B(_04127_),
    .X(_04444_));
 sg13g2_nor4_2 _21051_ (.A(_04044_),
    .B(_04442_),
    .C(_04443_),
    .Y(_04445_),
    .D(_04444_));
 sg13g2_nor2_1 _21052_ (.A(net5919),
    .B(_04033_),
    .Y(_04446_));
 sg13g2_a21o_1 _21053_ (.A2(_04446_),
    .A1(net5881),
    .B1(_04188_),
    .X(_04447_));
 sg13g2_o21ai_1 _21054_ (.B1(net5889),
    .Y(_04448_),
    .A1(net5899),
    .A2(net5845));
 sg13g2_o21ai_1 _21055_ (.B1(_04056_),
    .Y(_04449_),
    .A1(_04127_),
    .A2(_04448_));
 sg13g2_a21oi_1 _21056_ (.A1(_04103_),
    .A2(_04447_),
    .Y(_04450_),
    .B1(_04449_));
 sg13g2_a21oi_1 _21057_ (.A1(net5901),
    .A2(_04446_),
    .Y(_04451_),
    .B1(net5885));
 sg13g2_nand2_1 _21058_ (.Y(_04452_),
    .A(_04124_),
    .B(_04451_));
 sg13g2_a22oi_1 _21059_ (.Y(_04453_),
    .B1(_04188_),
    .B2(_04307_),
    .A2(_04109_),
    .A1(_03817_));
 sg13g2_a21oi_1 _21060_ (.A1(_04452_),
    .A2(_04453_),
    .Y(_04454_),
    .B1(_04024_));
 sg13g2_nor4_2 _21061_ (.A(_04441_),
    .B(_04445_),
    .C(_04450_),
    .Y(_04455_),
    .D(_04454_));
 sg13g2_xnor2_1 _21062_ (.Y(_04456_),
    .A(_04428_),
    .B(_04455_));
 sg13g2_nand2b_1 _21063_ (.Y(_04457_),
    .B(_04456_),
    .A_N(_04436_));
 sg13g2_xor2_1 _21064_ (.B(_04456_),
    .A(_04436_),
    .X(_04458_));
 sg13g2_a21oi_2 _21065_ (.B1(_04431_),
    .Y(_04459_),
    .A2(_04434_),
    .A1(_04432_));
 sg13g2_xnor2_1 _21066_ (.Y(_04460_),
    .A(_04458_),
    .B(_04459_));
 sg13g2_nor2_1 _21067_ (.A(net5984),
    .B(_04460_),
    .Y(_00323_));
 sg13g2_nand2_2 _21068_ (.Y(_04461_),
    .A(\b_pwm_odd[6] ),
    .B(net6013));
 sg13g2_a21oi_2 _21069_ (.B1(_04427_),
    .Y(_04462_),
    .A2(_04455_),
    .A1(_04403_));
 sg13g2_nand3_1 _21070_ (.B(_04124_),
    .C(_04317_),
    .A(net5881),
    .Y(_04463_));
 sg13g2_o21ai_1 _21071_ (.B1(_04161_),
    .Y(_04464_),
    .A1(net5926),
    .A2(_04149_));
 sg13g2_nand3_1 _21072_ (.B(_04463_),
    .C(_04464_),
    .A(_04018_),
    .Y(_04465_));
 sg13g2_nor2_1 _21073_ (.A(_03724_),
    .B(_04247_),
    .Y(_04466_));
 sg13g2_nor2_1 _21074_ (.A(_04222_),
    .B(_04466_),
    .Y(_04467_));
 sg13g2_nor2_1 _21075_ (.A(_04053_),
    .B(_04467_),
    .Y(_04468_));
 sg13g2_a21oi_1 _21076_ (.A1(_04163_),
    .A2(_04202_),
    .Y(_04469_),
    .B1(_04344_));
 sg13g2_nor3_1 _21077_ (.A(_03924_),
    .B(_04468_),
    .C(_04469_),
    .Y(_04470_));
 sg13g2_o21ai_1 _21078_ (.B1(_04144_),
    .Y(_04471_),
    .A1(_03724_),
    .A2(_04119_));
 sg13g2_nand3_1 _21079_ (.B(_04245_),
    .C(_04417_),
    .A(net5889),
    .Y(_04472_));
 sg13g2_nand3_1 _21080_ (.B(_04471_),
    .C(_04472_),
    .A(_04018_),
    .Y(_04473_));
 sg13g2_a21oi_1 _21081_ (.A1(_03719_),
    .A2(_04027_),
    .Y(_04474_),
    .B1(net5904));
 sg13g2_nor3_1 _21082_ (.A(_04053_),
    .B(_04147_),
    .C(_04474_),
    .Y(_04475_));
 sg13g2_or3_1 _21083_ (.A(net5898),
    .B(net5926),
    .C(_04048_),
    .X(_04476_));
 sg13g2_a21oi_1 _21084_ (.A1(_04075_),
    .A2(_04476_),
    .Y(_04477_),
    .B1(_04344_));
 sg13g2_nor2_1 _21085_ (.A(_04475_),
    .B(_04477_),
    .Y(_04478_));
 sg13g2_and2_1 _21086_ (.A(_04473_),
    .B(_04478_),
    .X(_04479_));
 sg13g2_a22oi_1 _21087_ (.Y(_04480_),
    .B1(_04479_),
    .B2(net5918),
    .A2(_04470_),
    .A1(_04465_));
 sg13g2_nor2_1 _21088_ (.A(_04455_),
    .B(_04480_),
    .Y(_04481_));
 sg13g2_nand2_1 _21089_ (.Y(_04482_),
    .A(_04455_),
    .B(_04480_));
 sg13g2_nand2b_1 _21090_ (.Y(_04483_),
    .B(_04482_),
    .A_N(_04481_));
 sg13g2_xor2_1 _21091_ (.B(_04483_),
    .A(_04462_),
    .X(_04484_));
 sg13g2_nor2_1 _21092_ (.A(_04461_),
    .B(_04484_),
    .Y(_04485_));
 sg13g2_xor2_1 _21093_ (.B(_04484_),
    .A(_04461_),
    .X(_04486_));
 sg13g2_o21ai_1 _21094_ (.B1(_04457_),
    .Y(_04487_),
    .A1(_04458_),
    .A2(_04459_));
 sg13g2_xnor2_1 _21095_ (.Y(_04488_),
    .A(_04486_),
    .B(_04487_));
 sg13g2_nor2_1 _21096_ (.A(net5984),
    .B(_04488_),
    .Y(_00324_));
 sg13g2_nand2_2 _21097_ (.Y(_04489_),
    .A(\b_pwm_odd[7] ),
    .B(net6013));
 sg13g2_and2_1 _21098_ (.A(_04188_),
    .B(_04349_),
    .X(_04490_));
 sg13g2_o21ai_1 _21099_ (.B1(_04195_),
    .Y(_04491_),
    .A1(_04068_),
    .A2(_04079_));
 sg13g2_nor4_1 _21100_ (.A(net5918),
    .B(_04192_),
    .C(_04490_),
    .D(_04491_),
    .Y(_04492_));
 sg13g2_a21oi_1 _21101_ (.A1(_03828_),
    .A2(_04047_),
    .Y(_04493_),
    .B1(_04053_));
 sg13g2_a21oi_1 _21102_ (.A1(_04159_),
    .A2(_04368_),
    .Y(_04494_),
    .B1(_04493_));
 sg13g2_o21ai_1 _21103_ (.B1(_04494_),
    .Y(_04495_),
    .A1(net5877),
    .A2(_04492_));
 sg13g2_o21ai_1 _21104_ (.B1(_04189_),
    .Y(_04496_),
    .A1(net5893),
    .A2(_04079_));
 sg13g2_o21ai_1 _21105_ (.B1(net5849),
    .Y(_04497_),
    .A1(_04353_),
    .A2(_04496_));
 sg13g2_a221oi_1 _21106_ (.B2(_03828_),
    .C1(net5849),
    .B1(_04205_),
    .A1(_03829_),
    .Y(_04498_),
    .A2(_04182_));
 sg13g2_nand2_1 _21107_ (.Y(_04499_),
    .A(net5918),
    .B(_04497_));
 sg13g2_o21ai_1 _21108_ (.B1(_04495_),
    .Y(_04500_),
    .A1(_04498_),
    .A2(_04499_));
 sg13g2_inv_1 _21109_ (.Y(_04501_),
    .A(_04500_));
 sg13g2_nand2b_1 _21110_ (.Y(_04502_),
    .B(_04500_),
    .A_N(_04480_));
 sg13g2_xor2_1 _21111_ (.B(_04500_),
    .A(_04480_),
    .X(_04503_));
 sg13g2_a21oi_2 _21112_ (.B1(_04481_),
    .Y(_04504_),
    .A2(_04482_),
    .A1(_04462_));
 sg13g2_or2_1 _21113_ (.X(_04505_),
    .B(_04504_),
    .A(_04503_));
 sg13g2_xor2_1 _21114_ (.B(_04504_),
    .A(_04503_),
    .X(_04506_));
 sg13g2_xnor2_1 _21115_ (.Y(_04507_),
    .A(_04503_),
    .B(_04504_));
 sg13g2_nand2b_1 _21116_ (.Y(_04508_),
    .B(_04506_),
    .A_N(_04489_));
 sg13g2_xnor2_1 _21117_ (.Y(_04509_),
    .A(_04489_),
    .B(_04506_));
 sg13g2_a21oi_2 _21118_ (.B1(_04485_),
    .Y(_04510_),
    .A2(_04487_),
    .A1(_04486_));
 sg13g2_nand2b_1 _21119_ (.Y(_04511_),
    .B(_04509_),
    .A_N(_04510_));
 sg13g2_xor2_1 _21120_ (.B(_04510_),
    .A(_04509_),
    .X(_04512_));
 sg13g2_nor2_1 _21121_ (.A(net5984),
    .B(_04512_),
    .Y(_00325_));
 sg13g2_nand2_2 _21122_ (.Y(_04513_),
    .A(_04508_),
    .B(_04511_));
 sg13g2_o21ai_1 _21123_ (.B1(net5888),
    .Y(_04514_),
    .A1(net5897),
    .A2(_03720_));
 sg13g2_nand2b_1 _21124_ (.Y(_04515_),
    .B(_04142_),
    .A_N(_04514_));
 sg13g2_nor2_1 _21125_ (.A(net5888),
    .B(net5876),
    .Y(_04516_));
 sg13g2_o21ai_1 _21126_ (.B1(_04516_),
    .Y(_04517_),
    .A1(net5904),
    .A2(_04101_));
 sg13g2_nand3_1 _21127_ (.B(_04515_),
    .C(_04517_),
    .A(_04021_),
    .Y(_04518_));
 sg13g2_a21oi_1 _21128_ (.A1(_03718_),
    .A2(_03814_),
    .Y(_04519_),
    .B1(_04184_));
 sg13g2_o21ai_1 _21129_ (.B1(net5877),
    .Y(_04520_),
    .A1(_04078_),
    .A2(_04519_));
 sg13g2_o21ai_1 _21130_ (.B1(_04195_),
    .Y(_04521_),
    .A1(_04034_),
    .A2(_04079_));
 sg13g2_o21ai_1 _21131_ (.B1(net5848),
    .Y(_04522_),
    .A1(_04219_),
    .A2(_04521_));
 sg13g2_a221oi_1 _21132_ (.B2(net5904),
    .C1(_04101_),
    .B1(_04034_),
    .A1(net6089),
    .Y(_04523_),
    .A2(_03814_));
 sg13g2_o21ai_1 _21133_ (.B1(net5816),
    .Y(_04524_),
    .A1(_04227_),
    .A2(_04523_));
 sg13g2_nand4_1 _21134_ (.B(_04520_),
    .C(_04522_),
    .A(_04518_),
    .Y(_04525_),
    .D(_04524_));
 sg13g2_xor2_1 _21135_ (.B(_04525_),
    .A(_04500_),
    .X(_04526_));
 sg13g2_a21o_1 _21136_ (.A2(_04505_),
    .A1(_04502_),
    .B1(_04526_),
    .X(_04527_));
 sg13g2_nand3_1 _21137_ (.B(_04505_),
    .C(_04526_),
    .A(_04502_),
    .Y(_04528_));
 sg13g2_nand2_1 _21138_ (.Y(_04529_),
    .A(_04527_),
    .B(_04528_));
 sg13g2_nand3_1 _21139_ (.B(_04511_),
    .C(_04529_),
    .A(_04508_),
    .Y(_04530_));
 sg13g2_nand2b_1 _21140_ (.Y(_04531_),
    .B(_04513_),
    .A_N(_04529_));
 sg13g2_and3_1 _21141_ (.X(_00326_),
    .A(net5980),
    .B(_04530_),
    .C(_04531_));
 sg13g2_a21oi_2 _21142_ (.B1(_04525_),
    .Y(_04532_),
    .A2(_04505_),
    .A1(_04501_));
 sg13g2_a21o_1 _21143_ (.A2(_04527_),
    .A1(_04525_),
    .B1(_04532_),
    .X(_04533_));
 sg13g2_and2_1 _21144_ (.A(_04531_),
    .B(_04533_),
    .X(_04534_));
 sg13g2_nor2_1 _21145_ (.A(_04531_),
    .B(_04533_),
    .Y(_04535_));
 sg13g2_nor3_2 _21146_ (.A(net5985),
    .B(_04534_),
    .C(_04535_),
    .Y(_00327_));
 sg13g2_nor2_1 _21147_ (.A(_04532_),
    .B(_04535_),
    .Y(_04536_));
 sg13g2_nor2_2 _21148_ (.A(net5984),
    .B(_04536_),
    .Y(_00328_));
 sg13g2_nor2_1 _21149_ (.A(net2988),
    .B(\r_pwm_even[2] ),
    .Y(_04537_));
 sg13g2_nand3_1 _21150_ (.B(\r_pwm_even[2] ),
    .C(net6016),
    .A(net2988),
    .Y(_04538_));
 sg13g2_nand2_1 _21151_ (.Y(_04539_),
    .A(net6016),
    .B(_04538_));
 sg13g2_nor2_1 _21152_ (.A(_04537_),
    .B(_04539_),
    .Y(_04540_));
 sg13g2_nand3_1 _21153_ (.B(net7450),
    .C(net6016),
    .A(net7357),
    .Y(_04541_));
 sg13g2_o21ai_1 _21154_ (.B1(_04541_),
    .Y(_04542_),
    .A1(_04537_),
    .A2(_04539_));
 sg13g2_nand3_1 _21155_ (.B(net7450),
    .C(_04540_),
    .A(net7357),
    .Y(_04543_));
 sg13g2_and3_1 _21156_ (.X(_00329_),
    .A(net5981),
    .B(net7451),
    .C(net7358));
 sg13g2_xor2_1 _21157_ (.B(\r_pwm_even[3] ),
    .A(\r_pwm_odd[3] ),
    .X(_04544_));
 sg13g2_nand2b_1 _21158_ (.Y(_04545_),
    .B(_04544_),
    .A_N(_04538_));
 sg13g2_mux2_1 _21159_ (.A0(_04538_),
    .A1(_04539_),
    .S(_04544_),
    .X(_04546_));
 sg13g2_o21ai_1 _21160_ (.B1(net5981),
    .Y(_04547_),
    .A1(net7358),
    .A2(_04546_));
 sg13g2_a21oi_1 _21161_ (.A1(net7358),
    .A2(_04546_),
    .Y(_00330_),
    .B1(_04547_));
 sg13g2_o21ai_1 _21162_ (.B1(_04545_),
    .Y(_04548_),
    .A1(_04543_),
    .A2(_04546_));
 sg13g2_inv_1 _21163_ (.Y(_04549_),
    .A(_04548_));
 sg13g2_nand2_1 _21164_ (.Y(_04550_),
    .A(\r_pwm_even[4] ),
    .B(net6017));
 sg13g2_nor2_1 _21165_ (.A(_04098_),
    .B(_04550_),
    .Y(_04551_));
 sg13g2_xor2_1 _21166_ (.B(_04550_),
    .A(_04098_),
    .X(_04552_));
 sg13g2_xnor2_1 _21167_ (.Y(_04553_),
    .A(_04094_),
    .B(_04552_));
 sg13g2_nor2_1 _21168_ (.A(\r_pwm_even[3] ),
    .B(_04062_),
    .Y(_04554_));
 sg13g2_nor2_1 _21169_ (.A(_04065_),
    .B(_04554_),
    .Y(_04555_));
 sg13g2_nand2_1 _21170_ (.Y(_04556_),
    .A(_04553_),
    .B(_04555_));
 sg13g2_xnor2_1 _21171_ (.Y(_04557_),
    .A(_04553_),
    .B(_04555_));
 sg13g2_o21ai_1 _21172_ (.B1(net5981),
    .Y(_04558_),
    .A1(_04549_),
    .A2(_04557_));
 sg13g2_a21oi_1 _21173_ (.A1(_04549_),
    .A2(_04557_),
    .Y(_00331_),
    .B1(_04558_));
 sg13g2_o21ai_1 _21174_ (.B1(_04556_),
    .Y(_04559_),
    .A1(_04549_),
    .A2(_04557_));
 sg13g2_and2_1 _21175_ (.A(\r_pwm_even[5] ),
    .B(net6016),
    .X(_04560_));
 sg13g2_xnor2_1 _21176_ (.Y(_04561_),
    .A(_04138_),
    .B(_04560_));
 sg13g2_nor2_1 _21177_ (.A(_04134_),
    .B(_04561_),
    .Y(_04562_));
 sg13g2_xor2_1 _21178_ (.B(_04561_),
    .A(_04134_),
    .X(_04563_));
 sg13g2_a21oi_1 _21179_ (.A1(_04095_),
    .A2(_04552_),
    .Y(_04564_),
    .B1(_04551_));
 sg13g2_nor2b_1 _21180_ (.A(_04564_),
    .B_N(_04563_),
    .Y(_04565_));
 sg13g2_xnor2_1 _21181_ (.Y(_04566_),
    .A(_04563_),
    .B(_04564_));
 sg13g2_a21oi_1 _21182_ (.A1(_04559_),
    .A2(_04566_),
    .Y(_04567_),
    .B1(net5987));
 sg13g2_o21ai_1 _21183_ (.B1(_04567_),
    .Y(_04568_),
    .A1(_04559_),
    .A2(_04566_));
 sg13g2_inv_1 _21184_ (.Y(_00332_),
    .A(_04568_));
 sg13g2_a21oi_1 _21185_ (.A1(_04559_),
    .A2(_04566_),
    .Y(_04569_),
    .B1(_04565_));
 sg13g2_nand2_1 _21186_ (.Y(_04570_),
    .A(\r_pwm_even[6] ),
    .B(net6016));
 sg13g2_and3_1 _21187_ (.X(_04571_),
    .A(\r_pwm_even[6] ),
    .B(net6016),
    .C(_04177_));
 sg13g2_xor2_1 _21188_ (.B(_04570_),
    .A(_04177_),
    .X(_04572_));
 sg13g2_inv_1 _21189_ (.Y(_04573_),
    .A(_04572_));
 sg13g2_xor2_1 _21190_ (.B(_04572_),
    .A(_04172_),
    .X(_04574_));
 sg13g2_a21oi_1 _21191_ (.A1(_04138_),
    .A2(_04560_),
    .Y(_04575_),
    .B1(_04562_));
 sg13g2_nor2_1 _21192_ (.A(_04574_),
    .B(_04575_),
    .Y(_04576_));
 sg13g2_xnor2_1 _21193_ (.Y(_04577_),
    .A(_04574_),
    .B(_04575_));
 sg13g2_nor2_1 _21194_ (.A(_04569_),
    .B(_04577_),
    .Y(_04578_));
 sg13g2_a21oi_1 _21195_ (.A1(_04569_),
    .A2(_04577_),
    .Y(_04579_),
    .B1(net5987));
 sg13g2_nor2b_1 _21196_ (.A(_04578_),
    .B_N(_04579_),
    .Y(_00333_));
 sg13g2_or2_1 _21197_ (.X(_04580_),
    .B(_04578_),
    .A(_04576_));
 sg13g2_and2_1 _21198_ (.A(\r_pwm_even[7] ),
    .B(net6015),
    .X(_04581_));
 sg13g2_xnor2_1 _21199_ (.Y(_04582_),
    .A(_04217_),
    .B(_04581_));
 sg13g2_nor2_1 _21200_ (.A(_04213_),
    .B(_04582_),
    .Y(_04583_));
 sg13g2_xor2_1 _21201_ (.B(_04582_),
    .A(_04213_),
    .X(_04584_));
 sg13g2_a21oi_1 _21202_ (.A1(_04172_),
    .A2(_04573_),
    .Y(_04585_),
    .B1(_04571_));
 sg13g2_nor2b_1 _21203_ (.A(_04585_),
    .B_N(_04584_),
    .Y(_04586_));
 sg13g2_xnor2_1 _21204_ (.Y(_04587_),
    .A(_04584_),
    .B(_04585_));
 sg13g2_nor2_1 _21205_ (.A(_04580_),
    .B(_04587_),
    .Y(_04588_));
 sg13g2_and2_1 _21206_ (.A(_04580_),
    .B(_04587_),
    .X(_04589_));
 sg13g2_nor3_1 _21207_ (.A(net5987),
    .B(_04588_),
    .C(_04589_),
    .Y(_00334_));
 sg13g2_nor2_1 _21208_ (.A(_04586_),
    .B(_04589_),
    .Y(_04590_));
 sg13g2_a21oi_1 _21209_ (.A1(_04217_),
    .A2(_04581_),
    .Y(_04591_),
    .B1(_04583_));
 sg13g2_nor2_1 _21210_ (.A(_04218_),
    .B(_04591_),
    .Y(_04592_));
 sg13g2_xnor2_1 _21211_ (.Y(_04593_),
    .A(_04218_),
    .B(_04591_));
 sg13g2_nor2_1 _21212_ (.A(_04590_),
    .B(_04593_),
    .Y(_04594_));
 sg13g2_a21oi_1 _21213_ (.A1(_04590_),
    .A2(_04593_),
    .Y(_04595_),
    .B1(net5986));
 sg13g2_nor2b_1 _21214_ (.A(_04594_),
    .B_N(_04595_),
    .Y(_00335_));
 sg13g2_nor2_1 _21215_ (.A(_04592_),
    .B(_04594_),
    .Y(_04596_));
 sg13g2_nand2_1 _21216_ (.Y(_04597_),
    .A(_04218_),
    .B(_04235_));
 sg13g2_nor2_1 _21217_ (.A(_04239_),
    .B(_04597_),
    .Y(_04598_));
 sg13g2_xnor2_1 _21218_ (.Y(_04599_),
    .A(_04239_),
    .B(_04597_));
 sg13g2_and2_1 _21219_ (.A(_04596_),
    .B(_04599_),
    .X(_04600_));
 sg13g2_nor2_1 _21220_ (.A(_04596_),
    .B(_04599_),
    .Y(_04601_));
 sg13g2_nor3_2 _21221_ (.A(net5986),
    .B(_04600_),
    .C(_04601_),
    .Y(_00336_));
 sg13g2_nor3_1 _21222_ (.A(_04238_),
    .B(_04598_),
    .C(_04601_),
    .Y(_04602_));
 sg13g2_a21oi_1 _21223_ (.A1(_04238_),
    .A2(_04601_),
    .Y(_04603_),
    .B1(net5986));
 sg13g2_nor2b_2 _21224_ (.A(_04602_),
    .B_N(_04603_),
    .Y(_00337_));
 sg13g2_nand3_1 _21225_ (.B(\g_pwm_even[2] ),
    .C(net6019),
    .A(net2991),
    .Y(_04604_));
 sg13g2_or2_1 _21226_ (.X(_04605_),
    .B(\g_pwm_even[2] ),
    .A(net2991));
 sg13g2_nand3_1 _21227_ (.B(_04604_),
    .C(_04605_),
    .A(net6018),
    .Y(_04606_));
 sg13g2_nand3_1 _21228_ (.B(\g_pwm_odd[1] ),
    .C(net6019),
    .A(net4275),
    .Y(_04607_));
 sg13g2_or2_1 _21229_ (.X(_04608_),
    .B(net4276),
    .A(_04606_));
 sg13g2_nand2_1 _21230_ (.Y(_04609_),
    .A(net5981),
    .B(_04608_));
 sg13g2_a21oi_1 _21231_ (.A1(_04606_),
    .A2(net4276),
    .Y(_00338_),
    .B1(_04609_));
 sg13g2_nand2_1 _21232_ (.Y(_04610_),
    .A(_04604_),
    .B(_04608_));
 sg13g2_or2_1 _21233_ (.X(_04611_),
    .B(_04266_),
    .A(\g_pwm_even[3] ));
 sg13g2_nand3_1 _21234_ (.B(\g_pwm_even[3] ),
    .C(net6019),
    .A(net7512),
    .Y(_04612_));
 sg13g2_nand2_1 _21235_ (.Y(_04613_),
    .A(_04611_),
    .B(net7513));
 sg13g2_and2_1 _21236_ (.A(_04610_),
    .B(_04613_),
    .X(_04614_));
 sg13g2_o21ai_1 _21237_ (.B1(net5981),
    .Y(_04615_),
    .A1(_04610_),
    .A2(_04613_));
 sg13g2_nor2_1 _21238_ (.A(_04614_),
    .B(net7514),
    .Y(_00339_));
 sg13g2_nand2_1 _21239_ (.Y(_04616_),
    .A(\g_pwm_even[4] ),
    .B(net6019));
 sg13g2_xnor2_1 _21240_ (.Y(_04617_),
    .A(_04269_),
    .B(_04270_));
 sg13g2_nor2b_1 _21241_ (.A(_04616_),
    .B_N(_04617_),
    .Y(_04618_));
 sg13g2_xnor2_1 _21242_ (.Y(_04619_),
    .A(_04616_),
    .B(_04617_));
 sg13g2_and2_1 _21243_ (.A(_04267_),
    .B(_04611_),
    .X(_04620_));
 sg13g2_nand2_1 _21244_ (.Y(_04621_),
    .A(_04619_),
    .B(_04620_));
 sg13g2_xor2_1 _21245_ (.B(_04620_),
    .A(_04619_),
    .X(_04622_));
 sg13g2_nand2_1 _21246_ (.Y(_04623_),
    .A(_04614_),
    .B(_04622_));
 sg13g2_o21ai_1 _21247_ (.B1(net5981),
    .Y(_04624_),
    .A1(_04614_),
    .A2(_04622_));
 sg13g2_nor2b_1 _21248_ (.A(_04624_),
    .B_N(_04623_),
    .Y(_00340_));
 sg13g2_nand2_1 _21249_ (.Y(_04625_),
    .A(_04621_),
    .B(_04623_));
 sg13g2_nand2_1 _21250_ (.Y(_04626_),
    .A(\g_pwm_even[5] ),
    .B(net6018));
 sg13g2_nor2_1 _21251_ (.A(_04311_),
    .B(_04315_),
    .Y(_04627_));
 sg13g2_xnor2_1 _21252_ (.Y(_04628_),
    .A(_04296_),
    .B(_04313_));
 sg13g2_nor2b_1 _21253_ (.A(_04626_),
    .B_N(_04628_),
    .Y(_04629_));
 sg13g2_xor2_1 _21254_ (.B(_04628_),
    .A(_04626_),
    .X(_04630_));
 sg13g2_a21oi_1 _21255_ (.A1(_04291_),
    .A2(_04295_),
    .Y(_04631_),
    .B1(_04618_));
 sg13g2_nor2_1 _21256_ (.A(_04630_),
    .B(_04631_),
    .Y(_04632_));
 sg13g2_xor2_1 _21257_ (.B(_04631_),
    .A(_04630_),
    .X(_04633_));
 sg13g2_nor2_1 _21258_ (.A(_04625_),
    .B(_04633_),
    .Y(_04634_));
 sg13g2_and2_1 _21259_ (.A(_04625_),
    .B(_04633_),
    .X(_04635_));
 sg13g2_nor3_1 _21260_ (.A(net5988),
    .B(_04634_),
    .C(_04635_),
    .Y(_00341_));
 sg13g2_nor2_1 _21261_ (.A(_04632_),
    .B(_04635_),
    .Y(_04636_));
 sg13g2_nand2_1 _21262_ (.Y(_04637_),
    .A(\g_pwm_even[6] ),
    .B(net6018));
 sg13g2_nor2_1 _21263_ (.A(_04338_),
    .B(_04342_),
    .Y(_04638_));
 sg13g2_xor2_1 _21264_ (.B(_04341_),
    .A(_04316_),
    .X(_04639_));
 sg13g2_nor2_1 _21265_ (.A(_04637_),
    .B(_04639_),
    .Y(_04640_));
 sg13g2_xor2_1 _21266_ (.B(_04639_),
    .A(_04637_),
    .X(_04641_));
 sg13g2_nor2_1 _21267_ (.A(_04627_),
    .B(_04629_),
    .Y(_04642_));
 sg13g2_nor2b_1 _21268_ (.A(_04642_),
    .B_N(_04641_),
    .Y(_04643_));
 sg13g2_xor2_1 _21269_ (.B(_04642_),
    .A(_04641_),
    .X(_04644_));
 sg13g2_nor2_1 _21270_ (.A(_04636_),
    .B(_04644_),
    .Y(_04645_));
 sg13g2_a21oi_1 _21271_ (.A1(_04636_),
    .A2(_04644_),
    .Y(_04646_),
    .B1(net5988));
 sg13g2_nor2b_1 _21272_ (.A(_04645_),
    .B_N(_04646_),
    .Y(_00342_));
 sg13g2_nand2_1 _21273_ (.Y(_04647_),
    .A(\g_pwm_even[7] ),
    .B(net6018));
 sg13g2_nor2_1 _21274_ (.A(_04361_),
    .B(_04365_),
    .Y(_04648_));
 sg13g2_xnor2_1 _21275_ (.Y(_04649_),
    .A(_04343_),
    .B(_04363_));
 sg13g2_nor2_1 _21276_ (.A(_04647_),
    .B(_04649_),
    .Y(_04650_));
 sg13g2_xor2_1 _21277_ (.B(_04649_),
    .A(_04647_),
    .X(_04651_));
 sg13g2_nor2_1 _21278_ (.A(_04638_),
    .B(_04640_),
    .Y(_04652_));
 sg13g2_nand2b_1 _21279_ (.Y(_04653_),
    .B(_04651_),
    .A_N(_04652_));
 sg13g2_xnor2_1 _21280_ (.Y(_04654_),
    .A(_04651_),
    .B(_04652_));
 sg13g2_nor3_1 _21281_ (.A(_04643_),
    .B(_04645_),
    .C(_04654_),
    .Y(_04655_));
 sg13g2_o21ai_1 _21282_ (.B1(_04654_),
    .Y(_04656_),
    .A1(_04643_),
    .A2(_04645_));
 sg13g2_nand2_1 _21283_ (.Y(_04657_),
    .A(net5982),
    .B(_04656_));
 sg13g2_nor2_1 _21284_ (.A(_04655_),
    .B(_04657_),
    .Y(_00343_));
 sg13g2_nand2_1 _21285_ (.Y(_04658_),
    .A(_04653_),
    .B(_04656_));
 sg13g2_o21ai_1 _21286_ (.B1(_04366_),
    .Y(_04659_),
    .A1(_04648_),
    .A2(_04650_));
 sg13g2_or3_1 _21287_ (.A(_04366_),
    .B(_04648_),
    .C(_04650_),
    .X(_04660_));
 sg13g2_and2_1 _21288_ (.A(_04659_),
    .B(_04660_),
    .X(_04661_));
 sg13g2_nand2_1 _21289_ (.Y(_04662_),
    .A(_04658_),
    .B(_04661_));
 sg13g2_o21ai_1 _21290_ (.B1(net5982),
    .Y(_04663_),
    .A1(_04658_),
    .A2(_04661_));
 sg13g2_nor2b_1 _21291_ (.A(_04663_),
    .B_N(_04662_),
    .Y(_00344_));
 sg13g2_nand2b_1 _21292_ (.Y(_04664_),
    .B(_04377_),
    .A_N(_04366_));
 sg13g2_nand3b_1 _21293_ (.B(_04377_),
    .C(_04381_),
    .Y(_04665_),
    .A_N(_04366_));
 sg13g2_xor2_1 _21294_ (.B(_04664_),
    .A(_04381_),
    .X(_04666_));
 sg13g2_and2_1 _21295_ (.A(_04659_),
    .B(_04662_),
    .X(_04667_));
 sg13g2_and2_1 _21296_ (.A(_04666_),
    .B(_04667_),
    .X(_04668_));
 sg13g2_nor2_1 _21297_ (.A(_04666_),
    .B(_04667_),
    .Y(_04669_));
 sg13g2_nor3_2 _21298_ (.A(net5984),
    .B(_04668_),
    .C(_04669_),
    .Y(_00345_));
 sg13g2_xor2_1 _21299_ (.B(_04669_),
    .A(_04380_),
    .X(_04670_));
 sg13g2_a21oi_2 _21300_ (.B1(net5984),
    .Y(_00346_),
    .A2(_04670_),
    .A1(_04665_));
 sg13g2_nor2b_2 _21301_ (.A(tia_vsync_last),
    .B_N(\atari2600.tia.vid_vsync ),
    .Y(_04671_));
 sg13g2_o21ai_1 _21302_ (.B1(net6570),
    .Y(_04672_),
    .A1(\frame_counter[0] ),
    .A2(_04671_));
 sg13g2_a21oi_1 _21303_ (.A1(_08569_),
    .A2(_04671_),
    .Y(_00347_),
    .B1(_04672_));
 sg13g2_o21ai_1 _21304_ (.B1(net6582),
    .Y(_04673_),
    .A1(\frame_counter[1] ),
    .A2(_04671_));
 sg13g2_a21oi_1 _21305_ (.A1(net4244),
    .A2(_04671_),
    .Y(_00348_),
    .B1(_04673_));
 sg13g2_o21ai_1 _21306_ (.B1(net6582),
    .Y(_04674_),
    .A1(net4244),
    .A2(_04671_));
 sg13g2_a21oi_1 _21307_ (.A1(_08568_),
    .A2(_04671_),
    .Y(_00349_),
    .B1(_04674_));
 sg13g2_nor4_2 _21308_ (.A(net2),
    .B(net1),
    .C(net3),
    .Y(_04675_),
    .D(_11079_));
 sg13g2_or4_2 _21309_ (.A(net2),
    .B(net1),
    .C(net3),
    .D(_11079_),
    .X(_04676_));
 sg13g2_nor2_1 _21310_ (.A(_08649_),
    .B(_08651_),
    .Y(_04677_));
 sg13g2_nand4_1 _21311_ (.B(\gamepad_pmod.decoder.data_reg[6] ),
    .C(\gamepad_pmod.decoder.data_reg[7] ),
    .A(\gamepad_pmod.decoder.data_reg[5] ),
    .Y(_04678_),
    .D(\gamepad_pmod.decoder.data_reg[8] ));
 sg13g2_nand4_1 _21312_ (.B(\gamepad_pmod.decoder.data_reg[4] ),
    .C(\gamepad_pmod.decoder.data_reg[10] ),
    .A(\gamepad_pmod.decoder.data_reg[0] ),
    .Y(_04679_),
    .D(_04677_));
 sg13g2_nor4_2 _21313_ (.A(_08642_),
    .B(_08643_),
    .C(_04678_),
    .Y(_04680_),
    .D(_04679_));
 sg13g2_nand2_2 _21314_ (.Y(_04681_),
    .A(\gamepad_pmod.decoder.data_reg[1] ),
    .B(_04680_));
 sg13g2_a21oi_1 _21315_ (.A1(net4350),
    .A2(_04681_),
    .Y(_04682_),
    .B1(_04676_));
 sg13g2_nor2_1 _21316_ (.A(net1),
    .B(_04682_),
    .Y(_04683_));
 sg13g2_nor3_1 _21317_ (.A(_08641_),
    .B(_04676_),
    .C(_04680_),
    .Y(_04684_));
 sg13g2_a21oi_2 _21318_ (.B1(_04684_),
    .Y(_04685_),
    .A2(_04676_),
    .A1(_08657_));
 sg13g2_a21oi_1 _21319_ (.A1(net7285),
    .A2(_04685_),
    .Y(_04686_),
    .B1(net6527));
 sg13g2_o21ai_1 _21320_ (.B1(_04686_),
    .Y(_00350_),
    .A1(_04683_),
    .A2(_04685_));
 sg13g2_a21oi_1 _21321_ (.A1(net4103),
    .A2(_04681_),
    .Y(_04687_),
    .B1(_04676_));
 sg13g2_nor2_2 _21322_ (.A(net2),
    .B(_04687_),
    .Y(_04688_));
 sg13g2_a21oi_1 _21323_ (.A1(net7234),
    .A2(_04685_),
    .Y(_04689_),
    .B1(net6527));
 sg13g2_o21ai_1 _21324_ (.B1(_04689_),
    .Y(_00351_),
    .A1(_04685_),
    .A2(_04688_));
 sg13g2_a21oi_1 _21325_ (.A1(net4450),
    .A2(_04681_),
    .Y(_04690_),
    .B1(_04676_));
 sg13g2_nor2_2 _21326_ (.A(net3),
    .B(_04690_),
    .Y(_04691_));
 sg13g2_a21oi_1 _21327_ (.A1(net7200),
    .A2(_04685_),
    .Y(_04692_),
    .B1(net6527));
 sg13g2_o21ai_1 _21328_ (.B1(_04692_),
    .Y(_00352_),
    .A1(_04685_),
    .A2(_04691_));
 sg13g2_a21oi_1 _21329_ (.A1(net3786),
    .A2(_04681_),
    .Y(_04693_),
    .B1(_04676_));
 sg13g2_nor2_1 _21330_ (.A(net4),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_a21oi_1 _21331_ (.A1(net7345),
    .A2(_04685_),
    .Y(_04695_),
    .B1(net6523));
 sg13g2_o21ai_1 _21332_ (.B1(_04695_),
    .Y(_00353_),
    .A1(_04685_),
    .A2(_04694_));
 sg13g2_o21ai_1 _21333_ (.B1(_04387_),
    .Y(_04696_),
    .A1(_08674_),
    .A2(_04386_));
 sg13g2_nor2b_1 _21334_ (.A(_04388_),
    .B_N(_04385_),
    .Y(_04697_));
 sg13g2_nand2b_1 _21335_ (.Y(_04698_),
    .B(_04385_),
    .A_N(_04388_));
 sg13g2_nor2_1 _21336_ (.A(_04384_),
    .B(_04385_),
    .Y(_04699_));
 sg13g2_nor2_1 _21337_ (.A(_04697_),
    .B(_04699_),
    .Y(_04700_));
 sg13g2_nand2_1 _21338_ (.Y(_04701_),
    .A(\b_pwm_even[2] ),
    .B(net6018));
 sg13g2_xnor2_1 _21339_ (.Y(_04702_),
    .A(_04700_),
    .B(_04701_));
 sg13g2_or2_1 _21340_ (.X(_04703_),
    .B(_04702_),
    .A(_04696_));
 sg13g2_nand2_2 _21341_ (.Y(_04704_),
    .A(net7557),
    .B(_04702_));
 sg13g2_and3_1 _21342_ (.X(_00354_),
    .A(net5982),
    .B(_04703_),
    .C(_04704_));
 sg13g2_and2_1 _21343_ (.A(\b_pwm_even[3] ),
    .B(net6014),
    .X(_04705_));
 sg13g2_or2_1 _21344_ (.X(_04706_),
    .B(_04411_),
    .A(_04403_));
 sg13g2_o21ai_1 _21345_ (.B1(_04406_),
    .Y(_04707_),
    .A1(_04403_),
    .A2(_04411_));
 sg13g2_nand3_1 _21346_ (.B(_04705_),
    .C(_04706_),
    .A(_04406_),
    .Y(_04708_));
 sg13g2_xnor2_1 _21347_ (.Y(_04709_),
    .A(_04705_),
    .B(_04707_));
 sg13g2_o21ai_1 _21348_ (.B1(_04698_),
    .Y(_04710_),
    .A1(_04699_),
    .A2(_04701_));
 sg13g2_nand2_1 _21349_ (.Y(_04711_),
    .A(_04709_),
    .B(_04710_));
 sg13g2_xnor2_1 _21350_ (.Y(_04712_),
    .A(_04709_),
    .B(_04710_));
 sg13g2_o21ai_1 _21351_ (.B1(net5982),
    .Y(_04713_),
    .A1(_04704_),
    .A2(_04712_));
 sg13g2_a21oi_1 _21352_ (.A1(net7558),
    .A2(_04712_),
    .Y(_00355_),
    .B1(_04713_));
 sg13g2_o21ai_1 _21353_ (.B1(_04711_),
    .Y(_04714_),
    .A1(_04704_),
    .A2(_04712_));
 sg13g2_nand2_1 _21354_ (.Y(_04715_),
    .A(\b_pwm_even[4] ),
    .B(net6013));
 sg13g2_xor2_1 _21355_ (.B(_04434_),
    .A(_04412_),
    .X(_04716_));
 sg13g2_nor2_1 _21356_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_xor2_1 _21357_ (.B(_04716_),
    .A(_04715_),
    .X(_04718_));
 sg13g2_nand2_1 _21358_ (.Y(_04719_),
    .A(_04706_),
    .B(_04708_));
 sg13g2_and2_1 _21359_ (.A(_04718_),
    .B(_04719_),
    .X(_04720_));
 sg13g2_xor2_1 _21360_ (.B(_04719_),
    .A(_04718_),
    .X(_04721_));
 sg13g2_o21ai_1 _21361_ (.B1(net5980),
    .Y(_04722_),
    .A1(_04714_),
    .A2(_04721_));
 sg13g2_a21oi_1 _21362_ (.A1(_04714_),
    .A2(_04721_),
    .Y(_00356_),
    .B1(_04722_));
 sg13g2_a21oi_2 _21363_ (.B1(_04720_),
    .Y(_04723_),
    .A2(_04721_),
    .A1(_04714_));
 sg13g2_nand2_1 _21364_ (.Y(_04724_),
    .A(\b_pwm_even[5] ),
    .B(net6013));
 sg13g2_nor2b_1 _21365_ (.A(_04460_),
    .B_N(_04456_),
    .Y(_04725_));
 sg13g2_xnor2_1 _21366_ (.Y(_04726_),
    .A(_04436_),
    .B(_04459_));
 sg13g2_nor2_1 _21367_ (.A(_04724_),
    .B(_04726_),
    .Y(_04727_));
 sg13g2_xor2_1 _21368_ (.B(_04726_),
    .A(_04724_),
    .X(_04728_));
 sg13g2_a21oi_1 _21369_ (.A1(_04430_),
    .A2(_04435_),
    .Y(_04729_),
    .B1(_04717_));
 sg13g2_nand2b_1 _21370_ (.Y(_04730_),
    .B(_04728_),
    .A_N(_04729_));
 sg13g2_xor2_1 _21371_ (.B(_04729_),
    .A(_04728_),
    .X(_04731_));
 sg13g2_o21ai_1 _21372_ (.B1(net5980),
    .Y(_04732_),
    .A1(_04723_),
    .A2(_04731_));
 sg13g2_a21oi_1 _21373_ (.A1(_04723_),
    .A2(_04731_),
    .Y(_00357_),
    .B1(_04732_));
 sg13g2_o21ai_1 _21374_ (.B1(_04730_),
    .Y(_04733_),
    .A1(_04723_),
    .A2(_04731_));
 sg13g2_nand2_1 _21375_ (.Y(_04734_),
    .A(\b_pwm_even[6] ),
    .B(net6013));
 sg13g2_nor2_1 _21376_ (.A(_04484_),
    .B(_04488_),
    .Y(_04735_));
 sg13g2_xor2_1 _21377_ (.B(_04487_),
    .A(_04461_),
    .X(_04736_));
 sg13g2_nor2_1 _21378_ (.A(_04734_),
    .B(_04736_),
    .Y(_04737_));
 sg13g2_xor2_1 _21379_ (.B(_04736_),
    .A(_04734_),
    .X(_04738_));
 sg13g2_nor2_1 _21380_ (.A(_04725_),
    .B(_04727_),
    .Y(_04739_));
 sg13g2_nand2b_1 _21381_ (.Y(_04740_),
    .B(_04738_),
    .A_N(_04739_));
 sg13g2_xnor2_1 _21382_ (.Y(_04741_),
    .A(_04738_),
    .B(_04739_));
 sg13g2_nand2_1 _21383_ (.Y(_04742_),
    .A(_04733_),
    .B(_04741_));
 sg13g2_o21ai_1 _21384_ (.B1(net5980),
    .Y(_04743_),
    .A1(_04733_),
    .A2(_04741_));
 sg13g2_nor2b_1 _21385_ (.A(_04743_),
    .B_N(_04742_),
    .Y(_00358_));
 sg13g2_nand2_1 _21386_ (.Y(_04744_),
    .A(\b_pwm_even[7] ),
    .B(net6013));
 sg13g2_xor2_1 _21387_ (.B(_04510_),
    .A(_04489_),
    .X(_04745_));
 sg13g2_nand2b_1 _21388_ (.Y(_04746_),
    .B(_04745_),
    .A_N(_04744_));
 sg13g2_xnor2_1 _21389_ (.Y(_04747_),
    .A(_04744_),
    .B(_04745_));
 sg13g2_nor2_1 _21390_ (.A(_04735_),
    .B(_04737_),
    .Y(_04748_));
 sg13g2_nand2b_1 _21391_ (.Y(_04749_),
    .B(_04747_),
    .A_N(_04748_));
 sg13g2_xor2_1 _21392_ (.B(_04748_),
    .A(_04747_),
    .X(_04750_));
 sg13g2_nand3_1 _21393_ (.B(_04742_),
    .C(_04750_),
    .A(_04740_),
    .Y(_04751_));
 sg13g2_a21o_1 _21394_ (.A2(_04742_),
    .A1(_04740_),
    .B1(_04750_),
    .X(_04752_));
 sg13g2_and3_1 _21395_ (.X(_00359_),
    .A(net5980),
    .B(_04751_),
    .C(_04752_));
 sg13g2_and2_1 _21396_ (.A(_04749_),
    .B(_04752_),
    .X(_04753_));
 sg13g2_o21ai_1 _21397_ (.B1(_04746_),
    .Y(_04754_),
    .A1(_04507_),
    .A2(_04512_));
 sg13g2_nand2_1 _21398_ (.Y(_04755_),
    .A(_04513_),
    .B(_04754_));
 sg13g2_xnor2_1 _21399_ (.Y(_04756_),
    .A(_04513_),
    .B(_04754_));
 sg13g2_or2_1 _21400_ (.X(_04757_),
    .B(_04756_),
    .A(_04753_));
 sg13g2_nand2_1 _21401_ (.Y(_04758_),
    .A(net5980),
    .B(_04757_));
 sg13g2_a21oi_1 _21402_ (.A1(_04753_),
    .A2(_04756_),
    .Y(_00360_),
    .B1(_04758_));
 sg13g2_and2_1 _21403_ (.A(_04755_),
    .B(_04757_),
    .X(_04759_));
 sg13g2_nor2_1 _21404_ (.A(_04513_),
    .B(_04529_),
    .Y(_04760_));
 sg13g2_nor3_1 _21405_ (.A(_04513_),
    .B(_04529_),
    .C(_04533_),
    .Y(_04761_));
 sg13g2_xor2_1 _21406_ (.B(_04760_),
    .A(_04533_),
    .X(_04762_));
 sg13g2_and2_1 _21407_ (.A(_04759_),
    .B(_04762_),
    .X(_04763_));
 sg13g2_nor2_1 _21408_ (.A(_04759_),
    .B(_04762_),
    .Y(_04764_));
 sg13g2_nor3_2 _21409_ (.A(net5985),
    .B(_04763_),
    .C(_04764_),
    .Y(_00361_));
 sg13g2_nor3_1 _21410_ (.A(_04532_),
    .B(_04761_),
    .C(_04764_),
    .Y(_04765_));
 sg13g2_a21oi_1 _21411_ (.A1(_04532_),
    .A2(_04764_),
    .Y(_04766_),
    .B1(net5984));
 sg13g2_nor2b_2 _21412_ (.A(_04765_),
    .B_N(_04766_),
    .Y(_00362_));
 sg13g2_nand3_1 _21413_ (.B(net5527),
    .C(_03092_),
    .A(net5557),
    .Y(_04767_));
 sg13g2_nor2_1 _21414_ (.A(_03091_),
    .B(net5236),
    .Y(_04768_));
 sg13g2_nor2_1 _21415_ (.A(net4472),
    .B(net5191),
    .Y(_04769_));
 sg13g2_a21oi_1 _21416_ (.A1(net5773),
    .A2(net5191),
    .Y(_00363_),
    .B1(_04769_));
 sg13g2_nor2_1 _21417_ (.A(net3714),
    .B(net5192),
    .Y(_04770_));
 sg13g2_a21oi_1 _21418_ (.A1(net5793),
    .A2(net5192),
    .Y(_00364_),
    .B1(_04770_));
 sg13g2_nor2_1 _21419_ (.A(net3333),
    .B(net5192),
    .Y(_04771_));
 sg13g2_a21oi_1 _21420_ (.A1(net5723),
    .A2(net5192),
    .Y(_00365_),
    .B1(_04771_));
 sg13g2_nor2_1 _21421_ (.A(net3322),
    .B(net5192),
    .Y(_04772_));
 sg13g2_a21oi_1 _21422_ (.A1(net5699),
    .A2(net5192),
    .Y(_00366_),
    .B1(_04772_));
 sg13g2_nor2_1 _21423_ (.A(net3854),
    .B(net5192),
    .Y(_04773_));
 sg13g2_a21oi_1 _21424_ (.A1(net5679),
    .A2(_04768_),
    .Y(_00367_),
    .B1(_04773_));
 sg13g2_nor2_1 _21425_ (.A(net3231),
    .B(net5191),
    .Y(_04774_));
 sg13g2_a21oi_1 _21426_ (.A1(net5599),
    .A2(net5191),
    .Y(_00368_),
    .B1(_04774_));
 sg13g2_nor2_1 _21427_ (.A(net3834),
    .B(net5191),
    .Y(_04775_));
 sg13g2_a21oi_1 _21428_ (.A1(net5661),
    .A2(net5191),
    .Y(_00369_),
    .B1(_04775_));
 sg13g2_nor2_1 _21429_ (.A(net3280),
    .B(net5191),
    .Y(_04776_));
 sg13g2_a21oi_1 _21430_ (.A1(net5633),
    .A2(net5191),
    .Y(_00370_),
    .B1(_04776_));
 sg13g2_nand2_2 _21431_ (.Y(_04777_),
    .A(_09264_),
    .B(net5252));
 sg13g2_mux2_1 _21432_ (.A0(net5741),
    .A1(net6674),
    .S(_04777_),
    .X(_00371_));
 sg13g2_mux2_1 _21433_ (.A0(net5744),
    .A1(net6681),
    .S(_04777_),
    .X(_00372_));
 sg13g2_mux2_1 _21434_ (.A0(net5617),
    .A1(net4496),
    .S(_04777_),
    .X(_00373_));
 sg13g2_mux2_1 _21435_ (.A0(net5614),
    .A1(net4893),
    .S(_04777_),
    .X(_00374_));
 sg13g2_mux2_1 _21436_ (.A0(net5608),
    .A1(net6802),
    .S(_04777_),
    .X(_00375_));
 sg13g2_mux2_1 _21437_ (.A0(net5581),
    .A1(net4817),
    .S(_04777_),
    .X(_00376_));
 sg13g2_mux2_1 _21438_ (.A0(net5578),
    .A1(net6669),
    .S(_04777_),
    .X(_00377_));
 sg13g2_mux2_1 _21439_ (.A0(net5644),
    .A1(net4885),
    .S(_04777_),
    .X(_00378_));
 sg13g2_nor2_2 _21440_ (.A(net5266),
    .B(_03123_),
    .Y(_04778_));
 sg13g2_nand2_2 _21441_ (.Y(_04779_),
    .A(_09319_),
    .B(_03122_));
 sg13g2_nand2_2 _21442_ (.Y(_04780_),
    .A(net5253),
    .B(_04778_));
 sg13g2_mux2_1 _21443_ (.A0(net5742),
    .A1(net4788),
    .S(_04780_),
    .X(_00379_));
 sg13g2_mux2_1 _21444_ (.A0(net5747),
    .A1(net4701),
    .S(_04780_),
    .X(_00380_));
 sg13g2_mux2_1 _21445_ (.A0(net5619),
    .A1(net4625),
    .S(_04780_),
    .X(_00381_));
 sg13g2_mux2_1 _21446_ (.A0(net5613),
    .A1(net4944),
    .S(_04780_),
    .X(_00382_));
 sg13g2_mux2_1 _21447_ (.A0(net5609),
    .A1(net4899),
    .S(_04780_),
    .X(_00383_));
 sg13g2_mux2_1 _21448_ (.A0(net5584),
    .A1(net7121),
    .S(_04780_),
    .X(_00384_));
 sg13g2_mux2_1 _21449_ (.A0(net5577),
    .A1(net6656),
    .S(_04780_),
    .X(_00385_));
 sg13g2_mux2_1 _21450_ (.A0(net5643),
    .A1(net4839),
    .S(_04780_),
    .X(_00386_));
 sg13g2_nor2b_1 _21451_ (.A(_09437_),
    .B_N(_03026_),
    .Y(_04781_));
 sg13g2_nand2_2 _21452_ (.Y(_04782_),
    .A(_04778_),
    .B(net5251));
 sg13g2_mux2_1 _21453_ (.A0(net5742),
    .A1(net4764),
    .S(_04782_),
    .X(_00387_));
 sg13g2_mux2_1 _21454_ (.A0(net5747),
    .A1(net6913),
    .S(_04782_),
    .X(_00388_));
 sg13g2_mux2_1 _21455_ (.A0(net5618),
    .A1(net6889),
    .S(_04782_),
    .X(_00389_));
 sg13g2_mux2_1 _21456_ (.A0(net5613),
    .A1(net4915),
    .S(_04782_),
    .X(_00390_));
 sg13g2_mux2_1 _21457_ (.A0(net5609),
    .A1(net4878),
    .S(_04782_),
    .X(_00391_));
 sg13g2_mux2_1 _21458_ (.A0(net5583),
    .A1(net4681),
    .S(_04782_),
    .X(_00392_));
 sg13g2_mux2_1 _21459_ (.A0(net5578),
    .A1(net7015),
    .S(_04782_),
    .X(_00393_));
 sg13g2_mux2_1 _21460_ (.A0(net5644),
    .A1(net6739),
    .S(_04782_),
    .X(_00394_));
 sg13g2_nor2_1 _21461_ (.A(net5239),
    .B(_04779_),
    .Y(_04783_));
 sg13g2_nor2_1 _21462_ (.A(net3549),
    .B(net5189),
    .Y(_04784_));
 sg13g2_a21oi_1 _21463_ (.A1(net5774),
    .A2(net5189),
    .Y(_00395_),
    .B1(_04784_));
 sg13g2_nor2_1 _21464_ (.A(net3811),
    .B(net5189),
    .Y(_04785_));
 sg13g2_a21oi_1 _21465_ (.A1(net5795),
    .A2(net5189),
    .Y(_00396_),
    .B1(_04785_));
 sg13g2_nor2_1 _21466_ (.A(net4114),
    .B(net5189),
    .Y(_04786_));
 sg13g2_a21oi_1 _21467_ (.A1(net5725),
    .A2(net5189),
    .Y(_00397_),
    .B1(_04786_));
 sg13g2_nor2_1 _21468_ (.A(net3965),
    .B(net5189),
    .Y(_04787_));
 sg13g2_a21oi_1 _21469_ (.A1(net5700),
    .A2(net5189),
    .Y(_00398_),
    .B1(_04787_));
 sg13g2_nor2_1 _21470_ (.A(net4220),
    .B(net5190),
    .Y(_04788_));
 sg13g2_a21oi_1 _21471_ (.A1(net5680),
    .A2(net5190),
    .Y(_00399_),
    .B1(_04788_));
 sg13g2_nor2_1 _21472_ (.A(net3634),
    .B(net5190),
    .Y(_04789_));
 sg13g2_a21oi_1 _21473_ (.A1(net5601),
    .A2(net5190),
    .Y(_00400_),
    .B1(_04789_));
 sg13g2_nor2_1 _21474_ (.A(net3006),
    .B(net5190),
    .Y(_04790_));
 sg13g2_a21oi_1 _21475_ (.A1(net5663),
    .A2(net5190),
    .Y(_00401_),
    .B1(_04790_));
 sg13g2_nor2_1 _21476_ (.A(net3450),
    .B(net5190),
    .Y(_04791_));
 sg13g2_a21oi_1 _21477_ (.A1(net5639),
    .A2(net5190),
    .Y(_00402_),
    .B1(_04791_));
 sg13g2_nand2_1 _21478_ (.Y(_04792_),
    .A(_09337_),
    .B(_03026_));
 sg13g2_nor2_1 _21479_ (.A(_04779_),
    .B(net5248),
    .Y(_04793_));
 sg13g2_nor2_1 _21480_ (.A(net3198),
    .B(net5187),
    .Y(_04794_));
 sg13g2_a21oi_1 _21481_ (.A1(net5769),
    .A2(net5187),
    .Y(_00403_),
    .B1(_04794_));
 sg13g2_nor2_1 _21482_ (.A(net3527),
    .B(net5187),
    .Y(_04795_));
 sg13g2_a21oi_1 _21483_ (.A1(net5788),
    .A2(net5187),
    .Y(_00404_),
    .B1(_04795_));
 sg13g2_nor2_1 _21484_ (.A(net3167),
    .B(net5188),
    .Y(_04796_));
 sg13g2_a21oi_1 _21485_ (.A1(net5719),
    .A2(net5188),
    .Y(_00405_),
    .B1(_04796_));
 sg13g2_nor2_1 _21486_ (.A(net3056),
    .B(net5187),
    .Y(_04797_));
 sg13g2_a21oi_1 _21487_ (.A1(net5696),
    .A2(net5187),
    .Y(_00406_),
    .B1(_04797_));
 sg13g2_nor2_1 _21488_ (.A(net3021),
    .B(net5187),
    .Y(_04798_));
 sg13g2_a21oi_1 _21489_ (.A1(net5682),
    .A2(net5187),
    .Y(_00407_),
    .B1(_04798_));
 sg13g2_nor2_1 _21490_ (.A(net3904),
    .B(net5188),
    .Y(_04799_));
 sg13g2_a21oi_1 _21491_ (.A1(net5601),
    .A2(_04793_),
    .Y(_00408_),
    .B1(_04799_));
 sg13g2_nor2_1 _21492_ (.A(net3355),
    .B(net5188),
    .Y(_04800_));
 sg13g2_a21oi_1 _21493_ (.A1(net5659),
    .A2(net5188),
    .Y(_00409_),
    .B1(_04800_));
 sg13g2_nor2_1 _21494_ (.A(net3733),
    .B(net5188),
    .Y(_04801_));
 sg13g2_a21oi_1 _21495_ (.A1(net5636),
    .A2(net5188),
    .Y(_00410_),
    .B1(_04801_));
 sg13g2_nor2_1 _21496_ (.A(net5254),
    .B(_04779_),
    .Y(_04802_));
 sg13g2_nor2_1 _21497_ (.A(net3902),
    .B(net5185),
    .Y(_04803_));
 sg13g2_a21oi_1 _21498_ (.A1(net5774),
    .A2(net5185),
    .Y(_00411_),
    .B1(_04803_));
 sg13g2_nor2_1 _21499_ (.A(net3406),
    .B(net5185),
    .Y(_04804_));
 sg13g2_a21oi_1 _21500_ (.A1(net5795),
    .A2(net5185),
    .Y(_00412_),
    .B1(_04804_));
 sg13g2_nor2_1 _21501_ (.A(net3207),
    .B(net5185),
    .Y(_04805_));
 sg13g2_a21oi_1 _21502_ (.A1(net5725),
    .A2(net5185),
    .Y(_00413_),
    .B1(_04805_));
 sg13g2_nor2_1 _21503_ (.A(net3139),
    .B(net5185),
    .Y(_04806_));
 sg13g2_a21oi_1 _21504_ (.A1(net5700),
    .A2(net5185),
    .Y(_00414_),
    .B1(_04806_));
 sg13g2_nor2_1 _21505_ (.A(net3565),
    .B(net5186),
    .Y(_04807_));
 sg13g2_a21oi_1 _21506_ (.A1(net5684),
    .A2(net5186),
    .Y(_00415_),
    .B1(_04807_));
 sg13g2_nor2_1 _21507_ (.A(net3405),
    .B(net5186),
    .Y(_04808_));
 sg13g2_a21oi_1 _21508_ (.A1(net5603),
    .A2(net5186),
    .Y(_00416_),
    .B1(_04808_));
 sg13g2_nor2_1 _21509_ (.A(net3403),
    .B(net5186),
    .Y(_04809_));
 sg13g2_a21oi_1 _21510_ (.A1(net5663),
    .A2(net5186),
    .Y(_00417_),
    .B1(_04809_));
 sg13g2_nor2_1 _21511_ (.A(net3474),
    .B(net5186),
    .Y(_04810_));
 sg13g2_a21oi_1 _21512_ (.A1(net5639),
    .A2(net5186),
    .Y(_00418_),
    .B1(_04810_));
 sg13g2_nor2_1 _21513_ (.A(net5236),
    .B(_04779_),
    .Y(_04811_));
 sg13g2_nor2_1 _21514_ (.A(net3116),
    .B(net5183),
    .Y(_04812_));
 sg13g2_a21oi_1 _21515_ (.A1(net5768),
    .A2(net5183),
    .Y(_00419_),
    .B1(_04812_));
 sg13g2_nor2_1 _21516_ (.A(net3156),
    .B(net5183),
    .Y(_04813_));
 sg13g2_a21oi_1 _21517_ (.A1(net5788),
    .A2(net5183),
    .Y(_00420_),
    .B1(_04813_));
 sg13g2_nor2_1 _21518_ (.A(net3449),
    .B(net5184),
    .Y(_04814_));
 sg13g2_a21oi_1 _21519_ (.A1(net5718),
    .A2(net5183),
    .Y(_00421_),
    .B1(_04814_));
 sg13g2_nor2_1 _21520_ (.A(net3182),
    .B(_04811_),
    .Y(_04815_));
 sg13g2_a21oi_1 _21521_ (.A1(net5700),
    .A2(net5183),
    .Y(_00422_),
    .B1(_04815_));
 sg13g2_nor2_1 _21522_ (.A(net3024),
    .B(net5183),
    .Y(_04816_));
 sg13g2_a21oi_1 _21523_ (.A1(net5682),
    .A2(net5183),
    .Y(_00423_),
    .B1(_04816_));
 sg13g2_nor2_1 _21524_ (.A(net3649),
    .B(net5184),
    .Y(_04817_));
 sg13g2_a21oi_1 _21525_ (.A1(net5601),
    .A2(net5184),
    .Y(_00424_),
    .B1(_04817_));
 sg13g2_nor2_1 _21526_ (.A(net3131),
    .B(net5184),
    .Y(_04818_));
 sg13g2_a21oi_1 _21527_ (.A1(net5657),
    .A2(net5184),
    .Y(_00425_),
    .B1(_04818_));
 sg13g2_nor2_1 _21528_ (.A(net3329),
    .B(net5184),
    .Y(_04819_));
 sg13g2_a21oi_1 _21529_ (.A1(net5636),
    .A2(net5184),
    .Y(_00426_),
    .B1(_04819_));
 sg13g2_nor2_1 _21530_ (.A(net5256),
    .B(_04779_),
    .Y(_04820_));
 sg13g2_nor2_1 _21531_ (.A(net4061),
    .B(net5181),
    .Y(_04821_));
 sg13g2_a21oi_1 _21532_ (.A1(net5775),
    .A2(net5181),
    .Y(_00427_),
    .B1(_04821_));
 sg13g2_nor2_1 _21533_ (.A(net4197),
    .B(net5181),
    .Y(_04822_));
 sg13g2_a21oi_1 _21534_ (.A1(net5794),
    .A2(net5181),
    .Y(_00428_),
    .B1(_04822_));
 sg13g2_nor2_1 _21535_ (.A(net3583),
    .B(net5181),
    .Y(_04823_));
 sg13g2_a21oi_1 _21536_ (.A1(net5725),
    .A2(net5181),
    .Y(_00429_),
    .B1(_04823_));
 sg13g2_nor2_1 _21537_ (.A(net3636),
    .B(net5181),
    .Y(_04824_));
 sg13g2_a21oi_1 _21538_ (.A1(net5702),
    .A2(net5181),
    .Y(_00430_),
    .B1(_04824_));
 sg13g2_nor2_1 _21539_ (.A(net4215),
    .B(net5182),
    .Y(_04825_));
 sg13g2_a21oi_1 _21540_ (.A1(net5684),
    .A2(net5182),
    .Y(_00431_),
    .B1(_04825_));
 sg13g2_nor2_1 _21541_ (.A(net4256),
    .B(net5182),
    .Y(_04826_));
 sg13g2_a21oi_1 _21542_ (.A1(net5603),
    .A2(net5182),
    .Y(_00432_),
    .B1(_04826_));
 sg13g2_nor2_1 _21543_ (.A(net3300),
    .B(net5182),
    .Y(_04827_));
 sg13g2_a21oi_1 _21544_ (.A1(net5663),
    .A2(net5182),
    .Y(_00433_),
    .B1(_04827_));
 sg13g2_nor2_1 _21545_ (.A(net3741),
    .B(net5182),
    .Y(_04828_));
 sg13g2_a21oi_1 _21546_ (.A1(net5639),
    .A2(net5182),
    .Y(_00434_),
    .B1(_04828_));
 sg13g2_nor2_1 _21547_ (.A(net5258),
    .B(_04779_),
    .Y(_04829_));
 sg13g2_nor2_1 _21548_ (.A(net4384),
    .B(net5180),
    .Y(_04830_));
 sg13g2_a21oi_1 _21549_ (.A1(net5768),
    .A2(net5180),
    .Y(_00435_),
    .B1(_04830_));
 sg13g2_nor2_1 _21550_ (.A(net3187),
    .B(net5179),
    .Y(_04831_));
 sg13g2_a21oi_1 _21551_ (.A1(net5788),
    .A2(net5179),
    .Y(_00436_),
    .B1(_04831_));
 sg13g2_nor2_1 _21552_ (.A(net3966),
    .B(net5179),
    .Y(_04832_));
 sg13g2_a21oi_1 _21553_ (.A1(net5718),
    .A2(net5179),
    .Y(_00437_),
    .B1(_04832_));
 sg13g2_nor2_1 _21554_ (.A(net3719),
    .B(net5180),
    .Y(_04833_));
 sg13g2_a21oi_1 _21555_ (.A1(net5700),
    .A2(net5180),
    .Y(_00438_),
    .B1(_04833_));
 sg13g2_nor2_1 _21556_ (.A(net3745),
    .B(net5180),
    .Y(_04834_));
 sg13g2_a21oi_1 _21557_ (.A1(net5682),
    .A2(net5180),
    .Y(_00439_),
    .B1(_04834_));
 sg13g2_nor2_1 _21558_ (.A(net3667),
    .B(net5180),
    .Y(_04835_));
 sg13g2_a21oi_1 _21559_ (.A1(net5601),
    .A2(_04829_),
    .Y(_00440_),
    .B1(_04835_));
 sg13g2_nor2_1 _21560_ (.A(net3221),
    .B(net5179),
    .Y(_04836_));
 sg13g2_a21oi_1 _21561_ (.A1(net5657),
    .A2(net5179),
    .Y(_00441_),
    .B1(_04836_));
 sg13g2_nor2_1 _21562_ (.A(net3530),
    .B(net5179),
    .Y(_04837_));
 sg13g2_a21oi_1 _21563_ (.A1(net5636),
    .A2(net5179),
    .Y(_00442_),
    .B1(_04837_));
 sg13g2_nor2_1 _21564_ (.A(_09331_),
    .B(net5238),
    .Y(_04838_));
 sg13g2_nor2_1 _21565_ (.A(net3703),
    .B(_04838_),
    .Y(_04839_));
 sg13g2_a21oi_1 _21566_ (.A1(net5763),
    .A2(net5070),
    .Y(_00443_),
    .B1(_04839_));
 sg13g2_nor2_1 _21567_ (.A(net3153),
    .B(net5069),
    .Y(_04840_));
 sg13g2_a21oi_1 _21568_ (.A1(net5782),
    .A2(net5069),
    .Y(_00444_),
    .B1(_04840_));
 sg13g2_nor2_1 _21569_ (.A(net3173),
    .B(net5070),
    .Y(_04841_));
 sg13g2_a21oi_1 _21570_ (.A1(net5712),
    .A2(net5070),
    .Y(_00445_),
    .B1(_04841_));
 sg13g2_nor2_1 _21571_ (.A(net3602),
    .B(net5069),
    .Y(_04842_));
 sg13g2_a21oi_1 _21572_ (.A1(net5690),
    .A2(net5069),
    .Y(_00446_),
    .B1(_04842_));
 sg13g2_nor2_1 _21573_ (.A(net3185),
    .B(net5070),
    .Y(_04843_));
 sg13g2_a21oi_1 _21574_ (.A1(net5669),
    .A2(net5070),
    .Y(_00447_),
    .B1(_04843_));
 sg13g2_nor2_1 _21575_ (.A(net3190),
    .B(net5069),
    .Y(_04844_));
 sg13g2_a21oi_1 _21576_ (.A1(net5591),
    .A2(net5069),
    .Y(_00448_),
    .B1(_04844_));
 sg13g2_nor2_1 _21577_ (.A(net3053),
    .B(net5069),
    .Y(_04845_));
 sg13g2_a21oi_1 _21578_ (.A1(net5650),
    .A2(net5069),
    .Y(_00449_),
    .B1(_04845_));
 sg13g2_nor2_1 _21579_ (.A(net3695),
    .B(net5070),
    .Y(_04846_));
 sg13g2_a21oi_1 _21580_ (.A1(net5629),
    .A2(net5070),
    .Y(_00450_),
    .B1(_04846_));
 sg13g2_nor2_1 _21581_ (.A(_03091_),
    .B(net5254),
    .Y(_04847_));
 sg13g2_nor2_1 _21582_ (.A(net3083),
    .B(net5177),
    .Y(_04848_));
 sg13g2_a21oi_1 _21583_ (.A1(net5772),
    .A2(net5177),
    .Y(_00451_),
    .B1(_04848_));
 sg13g2_nor2_1 _21584_ (.A(net3324),
    .B(net5178),
    .Y(_04849_));
 sg13g2_a21oi_1 _21585_ (.A1(net5792),
    .A2(net5178),
    .Y(_00452_),
    .B1(_04849_));
 sg13g2_nor2_1 _21586_ (.A(net3430),
    .B(net5178),
    .Y(_04850_));
 sg13g2_a21oi_1 _21587_ (.A1(net5722),
    .A2(net5178),
    .Y(_00453_),
    .B1(_04850_));
 sg13g2_nor2_1 _21588_ (.A(net3205),
    .B(net5178),
    .Y(_04851_));
 sg13g2_a21oi_1 _21589_ (.A1(net5699),
    .A2(net5178),
    .Y(_00454_),
    .B1(_04851_));
 sg13g2_nor2_1 _21590_ (.A(net3842),
    .B(net5177),
    .Y(_04852_));
 sg13g2_a21oi_1 _21591_ (.A1(net5679),
    .A2(net5178),
    .Y(_00455_),
    .B1(_04852_));
 sg13g2_nor2_1 _21592_ (.A(net3771),
    .B(net5177),
    .Y(_04853_));
 sg13g2_a21oi_1 _21593_ (.A1(net5598),
    .A2(_04847_),
    .Y(_00456_),
    .B1(_04853_));
 sg13g2_nor2_1 _21594_ (.A(net3005),
    .B(net5177),
    .Y(_04854_));
 sg13g2_a21oi_1 _21595_ (.A1(net5661),
    .A2(net5177),
    .Y(_00457_),
    .B1(_04854_));
 sg13g2_nor2_1 _21596_ (.A(net3976),
    .B(net5177),
    .Y(_04855_));
 sg13g2_a21oi_1 _21597_ (.A1(net5632),
    .A2(net5177),
    .Y(_00458_),
    .B1(_04855_));
 sg13g2_nor3_2 _21598_ (.A(net5995),
    .B(_09044_),
    .C(_09071_),
    .Y(_04856_));
 sg13g2_nand4_1 _21599_ (.B(_08803_),
    .C(_08823_),
    .A(_08796_),
    .Y(_04857_),
    .D(_08920_));
 sg13g2_a21oi_1 _21600_ (.A1(net6515),
    .A2(net6513),
    .Y(_04858_),
    .B1(net6521));
 sg13g2_nand2b_1 _21601_ (.Y(_04859_),
    .B(net6521),
    .A_N(net6515));
 sg13g2_xnor2_1 _21602_ (.Y(_04860_),
    .A(net6514),
    .B(_04859_));
 sg13g2_nor2_1 _21603_ (.A(net6515),
    .B(net6103),
    .Y(_04861_));
 sg13g2_a21oi_1 _21604_ (.A1(net6515),
    .A2(net6109),
    .Y(_04862_),
    .B1(_04861_));
 sg13g2_o21ai_1 _21605_ (.B1(\atari2600.cpu.state[1] ),
    .Y(_04863_),
    .A1(_04860_),
    .A2(_04862_));
 sg13g2_o21ai_1 _21606_ (.B1(_04863_),
    .Y(_04864_),
    .A1(_08797_),
    .A2(_04858_));
 sg13g2_nand4_1 _21607_ (.B(net5990),
    .C(_09074_),
    .A(_08847_),
    .Y(_04865_),
    .D(_04864_));
 sg13g2_nor4_1 _21608_ (.A(_08818_),
    .B(_09070_),
    .C(_04857_),
    .D(_04865_),
    .Y(_04866_));
 sg13g2_nand2_1 _21609_ (.Y(_04867_),
    .A(_04856_),
    .B(_04866_));
 sg13g2_and2_2 _21610_ (.A(_08879_),
    .B(_08939_),
    .X(_04868_));
 sg13g2_nand4_1 _21611_ (.B(_09011_),
    .C(_04867_),
    .A(net5856),
    .Y(_04869_),
    .D(_04868_));
 sg13g2_mux2_1 _21612_ (.A0(_09270_),
    .A1(net7431),
    .S(net5815),
    .X(_00459_));
 sg13g2_mux2_1 _21613_ (.A0(_09275_),
    .A1(net7399),
    .S(net5815),
    .X(_00460_));
 sg13g2_mux2_1 _21614_ (.A0(_09281_),
    .A1(net7398),
    .S(net5815),
    .X(_00461_));
 sg13g2_mux2_1 _21615_ (.A0(_09288_),
    .A1(net7425),
    .S(net5813),
    .X(_00462_));
 sg13g2_mux2_1 _21616_ (.A0(_09124_),
    .A1(net7356),
    .S(net5813),
    .X(_00463_));
 sg13g2_nand3_1 _21617_ (.B(_09345_),
    .C(net5253),
    .A(_09262_),
    .Y(_04870_));
 sg13g2_mux2_1 _21618_ (.A0(net5742),
    .A1(net6763),
    .S(_04870_),
    .X(_00464_));
 sg13g2_mux2_1 _21619_ (.A0(net5747),
    .A1(net4673),
    .S(_04870_),
    .X(_00465_));
 sg13g2_mux2_1 _21620_ (.A0(net5619),
    .A1(net4887),
    .S(_04870_),
    .X(_00466_));
 sg13g2_mux2_1 _21621_ (.A0(net5613),
    .A1(net4667),
    .S(_04870_),
    .X(_00467_));
 sg13g2_mux2_1 _21622_ (.A0(net5609),
    .A1(net4737),
    .S(_04870_),
    .X(_00468_));
 sg13g2_mux2_1 _21623_ (.A0(net5583),
    .A1(net7107),
    .S(_04870_),
    .X(_00469_));
 sg13g2_mux2_1 _21624_ (.A0(net5579),
    .A1(net4813),
    .S(_04870_),
    .X(_00470_));
 sg13g2_mux2_1 _21625_ (.A0(net5645),
    .A1(net6676),
    .S(_04870_),
    .X(_00471_));
 sg13g2_nor2_1 _21626_ (.A(_09331_),
    .B(net5255),
    .Y(_04871_));
 sg13g2_nor2_1 _21627_ (.A(net4345),
    .B(net5067),
    .Y(_04872_));
 sg13g2_a21oi_1 _21628_ (.A1(net5763),
    .A2(net5067),
    .Y(_00472_),
    .B1(_04872_));
 sg13g2_nor2_1 _21629_ (.A(net3142),
    .B(_04871_),
    .Y(_04873_));
 sg13g2_a21oi_1 _21630_ (.A1(net5782),
    .A2(net5068),
    .Y(_00473_),
    .B1(_04873_));
 sg13g2_nor2_1 _21631_ (.A(net3762),
    .B(net5067),
    .Y(_04874_));
 sg13g2_a21oi_1 _21632_ (.A1(net5713),
    .A2(net5067),
    .Y(_00474_),
    .B1(_04874_));
 sg13g2_nor2_1 _21633_ (.A(net3308),
    .B(net5068),
    .Y(_04875_));
 sg13g2_a21oi_1 _21634_ (.A1(net5690),
    .A2(net5068),
    .Y(_00475_),
    .B1(_04875_));
 sg13g2_nor2_1 _21635_ (.A(net3586),
    .B(net5067),
    .Y(_04876_));
 sg13g2_a21oi_1 _21636_ (.A1(net5669),
    .A2(net5067),
    .Y(_00476_),
    .B1(_04876_));
 sg13g2_nor2_1 _21637_ (.A(net3057),
    .B(net5068),
    .Y(_04877_));
 sg13g2_a21oi_1 _21638_ (.A1(net5591),
    .A2(net5068),
    .Y(_00477_),
    .B1(_04877_));
 sg13g2_nor2_1 _21639_ (.A(net3342),
    .B(net5068),
    .Y(_04878_));
 sg13g2_a21oi_1 _21640_ (.A1(net5650),
    .A2(net5068),
    .Y(_00478_),
    .B1(_04878_));
 sg13g2_nor2_1 _21641_ (.A(net3770),
    .B(net5067),
    .Y(_04879_));
 sg13g2_a21oi_1 _21642_ (.A1(net5629),
    .A2(net5067),
    .Y(_00479_),
    .B1(_04879_));
 sg13g2_nor2_1 _21643_ (.A(net5268),
    .B(_03123_),
    .Y(_04880_));
 sg13g2_nand2_2 _21644_ (.Y(_04881_),
    .A(_09301_),
    .B(_03122_));
 sg13g2_nor2_1 _21645_ (.A(net5248),
    .B(_04881_),
    .Y(_04882_));
 sg13g2_nor2_1 _21646_ (.A(net3039),
    .B(net5175),
    .Y(_04883_));
 sg13g2_a21oi_1 _21647_ (.A1(net5771),
    .A2(net5175),
    .Y(_00480_),
    .B1(_04883_));
 sg13g2_nor2_1 _21648_ (.A(net3111),
    .B(net5175),
    .Y(_04884_));
 sg13g2_a21oi_1 _21649_ (.A1(net5793),
    .A2(net5175),
    .Y(_00481_),
    .B1(_04884_));
 sg13g2_nor2_1 _21650_ (.A(net3567),
    .B(net5176),
    .Y(_04885_));
 sg13g2_a21oi_1 _21651_ (.A1(net5721),
    .A2(net5176),
    .Y(_00482_),
    .B1(_04885_));
 sg13g2_nor2_1 _21652_ (.A(net3310),
    .B(net5176),
    .Y(_04886_));
 sg13g2_a21oi_1 _21653_ (.A1(net5701),
    .A2(net5176),
    .Y(_00483_),
    .B1(_04886_));
 sg13g2_nor2_1 _21654_ (.A(net3100),
    .B(net5175),
    .Y(_04887_));
 sg13g2_a21oi_1 _21655_ (.A1(net5678),
    .A2(net5175),
    .Y(_00484_),
    .B1(_04887_));
 sg13g2_nor2_1 _21656_ (.A(net3582),
    .B(net5175),
    .Y(_04888_));
 sg13g2_a21oi_1 _21657_ (.A1(net5597),
    .A2(net5175),
    .Y(_00485_),
    .B1(_04888_));
 sg13g2_nor2_1 _21658_ (.A(net4689),
    .B(net5176),
    .Y(_04889_));
 sg13g2_a21oi_1 _21659_ (.A1(net5658),
    .A2(net5176),
    .Y(_00486_),
    .B1(_04889_));
 sg13g2_nor2_1 _21660_ (.A(net3674),
    .B(_04882_),
    .Y(_04890_));
 sg13g2_a21oi_1 _21661_ (.A1(net5635),
    .A2(net5176),
    .Y(_00487_),
    .B1(_04890_));
 sg13g2_nor2_1 _21662_ (.A(net5236),
    .B(_04881_),
    .Y(_04891_));
 sg13g2_nor2_1 _21663_ (.A(net4158),
    .B(net5173),
    .Y(_04892_));
 sg13g2_a21oi_1 _21664_ (.A1(net5771),
    .A2(net5173),
    .Y(_00488_),
    .B1(_04892_));
 sg13g2_nor2_1 _21665_ (.A(net3420),
    .B(net5173),
    .Y(_04893_));
 sg13g2_a21oi_1 _21666_ (.A1(net5793),
    .A2(net5173),
    .Y(_00489_),
    .B1(_04893_));
 sg13g2_nor2_1 _21667_ (.A(net3879),
    .B(net5174),
    .Y(_04894_));
 sg13g2_a21oi_1 _21668_ (.A1(net5721),
    .A2(net5174),
    .Y(_00490_),
    .B1(_04894_));
 sg13g2_nor2_1 _21669_ (.A(net3206),
    .B(net5174),
    .Y(_04895_));
 sg13g2_a21oi_1 _21670_ (.A1(net5701),
    .A2(net5174),
    .Y(_00491_),
    .B1(_04895_));
 sg13g2_nor2_1 _21671_ (.A(net3264),
    .B(net5173),
    .Y(_04896_));
 sg13g2_a21oi_1 _21672_ (.A1(net5678),
    .A2(net5173),
    .Y(_00492_),
    .B1(_04896_));
 sg13g2_nor2_1 _21673_ (.A(net3295),
    .B(net5173),
    .Y(_04897_));
 sg13g2_a21oi_1 _21674_ (.A1(net5597),
    .A2(net5173),
    .Y(_00493_),
    .B1(_04897_));
 sg13g2_nor2_1 _21675_ (.A(net4360),
    .B(net5174),
    .Y(_04898_));
 sg13g2_a21oi_1 _21676_ (.A1(net5658),
    .A2(net5174),
    .Y(_00494_),
    .B1(_04898_));
 sg13g2_nor2_1 _21677_ (.A(net3390),
    .B(net5174),
    .Y(_04899_));
 sg13g2_a21oi_1 _21678_ (.A1(net5637),
    .A2(net5174),
    .Y(_00495_),
    .B1(_04899_));
 sg13g2_nor2_1 _21679_ (.A(net5258),
    .B(_04881_),
    .Y(_04900_));
 sg13g2_nor2_1 _21680_ (.A(net3376),
    .B(net5171),
    .Y(_04901_));
 sg13g2_a21oi_1 _21681_ (.A1(net5771),
    .A2(net5171),
    .Y(_00496_),
    .B1(_04901_));
 sg13g2_nor2_1 _21682_ (.A(net3348),
    .B(net5171),
    .Y(_04902_));
 sg13g2_a21oi_1 _21683_ (.A1(net5791),
    .A2(net5171),
    .Y(_00497_),
    .B1(_04902_));
 sg13g2_nor2_1 _21684_ (.A(net3683),
    .B(net5172),
    .Y(_04903_));
 sg13g2_a21oi_1 _21685_ (.A1(net5721),
    .A2(net5172),
    .Y(_00498_),
    .B1(_04903_));
 sg13g2_nor2_1 _21686_ (.A(net3373),
    .B(net5172),
    .Y(_04904_));
 sg13g2_a21oi_1 _21687_ (.A1(net5701),
    .A2(net5172),
    .Y(_00499_),
    .B1(_04904_));
 sg13g2_nor2_1 _21688_ (.A(net3523),
    .B(net5171),
    .Y(_04905_));
 sg13g2_a21oi_1 _21689_ (.A1(net5678),
    .A2(net5171),
    .Y(_00500_),
    .B1(_04905_));
 sg13g2_nor2_1 _21690_ (.A(net4121),
    .B(net5171),
    .Y(_04906_));
 sg13g2_a21oi_1 _21691_ (.A1(net5596),
    .A2(net5171),
    .Y(_00501_),
    .B1(_04906_));
 sg13g2_nor2_1 _21692_ (.A(net3352),
    .B(net5172),
    .Y(_04907_));
 sg13g2_a21oi_1 _21693_ (.A1(net5658),
    .A2(net5172),
    .Y(_00502_),
    .B1(_04907_));
 sg13g2_nor2_1 _21694_ (.A(net3412),
    .B(net5172),
    .Y(_04908_));
 sg13g2_a21oi_1 _21695_ (.A1(net5637),
    .A2(net5172),
    .Y(_00503_),
    .B1(_04908_));
 sg13g2_nor2_1 _21696_ (.A(net5203),
    .B(net5249),
    .Y(_04909_));
 sg13g2_nor2_1 _21697_ (.A(net3037),
    .B(net5066),
    .Y(_04910_));
 sg13g2_a21oi_1 _21698_ (.A1(net5762),
    .A2(net5066),
    .Y(_00504_),
    .B1(_04910_));
 sg13g2_nor2_1 _21699_ (.A(net3117),
    .B(net5066),
    .Y(_04911_));
 sg13g2_a21oi_1 _21700_ (.A1(net5782),
    .A2(net5066),
    .Y(_00505_),
    .B1(_04911_));
 sg13g2_nor2_1 _21701_ (.A(net3041),
    .B(net5065),
    .Y(_04912_));
 sg13g2_a21oi_1 _21702_ (.A1(net5712),
    .A2(net5065),
    .Y(_00506_),
    .B1(_04912_));
 sg13g2_nor2_1 _21703_ (.A(net3702),
    .B(net5066),
    .Y(_04913_));
 sg13g2_a21oi_1 _21704_ (.A1(net5690),
    .A2(net5066),
    .Y(_00507_),
    .B1(_04913_));
 sg13g2_nor2_1 _21705_ (.A(net3265),
    .B(net5065),
    .Y(_04914_));
 sg13g2_a21oi_1 _21706_ (.A1(net5668),
    .A2(net5065),
    .Y(_00508_),
    .B1(_04914_));
 sg13g2_nor2_1 _21707_ (.A(net3233),
    .B(net5066),
    .Y(_04915_));
 sg13g2_a21oi_1 _21708_ (.A1(net5591),
    .A2(net5066),
    .Y(_00509_),
    .B1(_04915_));
 sg13g2_nor2_1 _21709_ (.A(net3957),
    .B(net5065),
    .Y(_04916_));
 sg13g2_a21oi_1 _21710_ (.A1(net5650),
    .A2(net5065),
    .Y(_00510_),
    .B1(_04916_));
 sg13g2_nor2_1 _21711_ (.A(net3038),
    .B(net5065),
    .Y(_04917_));
 sg13g2_a21oi_1 _21712_ (.A1(net5629),
    .A2(net5065),
    .Y(_00511_),
    .B1(_04917_));
 sg13g2_nor2_1 _21713_ (.A(net5239),
    .B(_04881_),
    .Y(_04918_));
 sg13g2_nor2_1 _21714_ (.A(net4218),
    .B(net5170),
    .Y(_04919_));
 sg13g2_a21oi_1 _21715_ (.A1(net5770),
    .A2(net5170),
    .Y(_00512_),
    .B1(_04919_));
 sg13g2_nor2_1 _21716_ (.A(net3941),
    .B(net5170),
    .Y(_04920_));
 sg13g2_a21oi_1 _21717_ (.A1(net5791),
    .A2(net5170),
    .Y(_00513_),
    .B1(_04920_));
 sg13g2_nor2_1 _21718_ (.A(net3340),
    .B(net5169),
    .Y(_04921_));
 sg13g2_a21oi_1 _21719_ (.A1(net5721),
    .A2(net5169),
    .Y(_00514_),
    .B1(_04921_));
 sg13g2_nor2_1 _21720_ (.A(net3540),
    .B(net5170),
    .Y(_04922_));
 sg13g2_a21oi_1 _21721_ (.A1(net5698),
    .A2(net5170),
    .Y(_00515_),
    .B1(_04922_));
 sg13g2_nor2_1 _21722_ (.A(net3159),
    .B(net5169),
    .Y(_04923_));
 sg13g2_a21oi_1 _21723_ (.A1(net5677),
    .A2(net5169),
    .Y(_00516_),
    .B1(_04923_));
 sg13g2_nor2_1 _21724_ (.A(net3258),
    .B(net5169),
    .Y(_04924_));
 sg13g2_a21oi_1 _21725_ (.A1(net5596),
    .A2(net5169),
    .Y(_00517_),
    .B1(_04924_));
 sg13g2_nor2_1 _21726_ (.A(net3133),
    .B(net5169),
    .Y(_04925_));
 sg13g2_a21oi_1 _21727_ (.A1(net5660),
    .A2(net5169),
    .Y(_00518_),
    .B1(_04925_));
 sg13g2_nor2_1 _21728_ (.A(net4254),
    .B(net5170),
    .Y(_04926_));
 sg13g2_a21oi_1 _21729_ (.A1(net5634),
    .A2(_04918_),
    .Y(_00519_),
    .B1(_04926_));
 sg13g2_nor2_1 _21730_ (.A(net5254),
    .B(_04881_),
    .Y(_04927_));
 sg13g2_nor2_1 _21731_ (.A(net3013),
    .B(net5167),
    .Y(_04928_));
 sg13g2_a21oi_1 _21732_ (.A1(net5770),
    .A2(net5167),
    .Y(_00520_),
    .B1(_04928_));
 sg13g2_nor2_1 _21733_ (.A(net3992),
    .B(net5168),
    .Y(_04929_));
 sg13g2_a21oi_1 _21734_ (.A1(net5791),
    .A2(net5168),
    .Y(_00521_),
    .B1(_04929_));
 sg13g2_nor2_1 _21735_ (.A(net3353),
    .B(net5168),
    .Y(_04930_));
 sg13g2_a21oi_1 _21736_ (.A1(net5723),
    .A2(net5168),
    .Y(_00522_),
    .B1(_04930_));
 sg13g2_nor2_1 _21737_ (.A(net3979),
    .B(net5167),
    .Y(_04931_));
 sg13g2_a21oi_1 _21738_ (.A1(net5698),
    .A2(net5167),
    .Y(_00523_),
    .B1(_04931_));
 sg13g2_nor2_1 _21739_ (.A(net3418),
    .B(net5167),
    .Y(_04932_));
 sg13g2_a21oi_1 _21740_ (.A1(net5677),
    .A2(net5167),
    .Y(_00524_),
    .B1(_04932_));
 sg13g2_nor2_1 _21741_ (.A(net3345),
    .B(net5168),
    .Y(_04933_));
 sg13g2_a21oi_1 _21742_ (.A1(net5596),
    .A2(net5168),
    .Y(_00525_),
    .B1(_04933_));
 sg13g2_nor2_1 _21743_ (.A(net3136),
    .B(net5167),
    .Y(_04934_));
 sg13g2_a21oi_1 _21744_ (.A1(net5660),
    .A2(net5167),
    .Y(_00526_),
    .B1(_04934_));
 sg13g2_nor2_1 _21745_ (.A(net3073),
    .B(net5168),
    .Y(_04935_));
 sg13g2_a21oi_1 _21746_ (.A1(net5634),
    .A2(net5168),
    .Y(_00527_),
    .B1(_04935_));
 sg13g2_nor2_1 _21747_ (.A(net5256),
    .B(_04881_),
    .Y(_04936_));
 sg13g2_nor2_1 _21748_ (.A(net4119),
    .B(net5165),
    .Y(_04937_));
 sg13g2_a21oi_1 _21749_ (.A1(net5770),
    .A2(net5165),
    .Y(_00528_),
    .B1(_04937_));
 sg13g2_nor2_1 _21750_ (.A(net3575),
    .B(net5166),
    .Y(_04938_));
 sg13g2_a21oi_1 _21751_ (.A1(net5791),
    .A2(net5166),
    .Y(_00529_),
    .B1(_04938_));
 sg13g2_nor2_1 _21752_ (.A(net3350),
    .B(net5166),
    .Y(_04939_));
 sg13g2_a21oi_1 _21753_ (.A1(net5723),
    .A2(net5166),
    .Y(_00530_),
    .B1(_04939_));
 sg13g2_nor2_1 _21754_ (.A(net3289),
    .B(net5165),
    .Y(_04940_));
 sg13g2_a21oi_1 _21755_ (.A1(net5698),
    .A2(net5165),
    .Y(_00531_),
    .B1(_04940_));
 sg13g2_nor2_1 _21756_ (.A(net4461),
    .B(net5165),
    .Y(_04941_));
 sg13g2_a21oi_1 _21757_ (.A1(net5685),
    .A2(net5165),
    .Y(_00532_),
    .B1(_04941_));
 sg13g2_nor2_1 _21758_ (.A(net4288),
    .B(net5166),
    .Y(_04942_));
 sg13g2_a21oi_1 _21759_ (.A1(net5596),
    .A2(net5166),
    .Y(_00533_),
    .B1(_04942_));
 sg13g2_nor2_1 _21760_ (.A(net4083),
    .B(net5165),
    .Y(_04943_));
 sg13g2_a21oi_1 _21761_ (.A1(net5660),
    .A2(net5165),
    .Y(_00534_),
    .B1(_04943_));
 sg13g2_nor2_1 _21762_ (.A(net4403),
    .B(net5166),
    .Y(_04944_));
 sg13g2_a21oi_1 _21763_ (.A1(net5634),
    .A2(net5166),
    .Y(_00535_),
    .B1(_04944_));
 sg13g2_nand2_2 _21764_ (.Y(_04945_),
    .A(net5253),
    .B(_04880_));
 sg13g2_mux2_1 _21765_ (.A0(net5741),
    .A1(net4656),
    .S(_04945_),
    .X(_00536_));
 sg13g2_mux2_1 _21766_ (.A0(net5746),
    .A1(net7014),
    .S(_04945_),
    .X(_00537_));
 sg13g2_mux2_1 _21767_ (.A0(net5620),
    .A1(net7087),
    .S(_04945_),
    .X(_00538_));
 sg13g2_mux2_1 _21768_ (.A0(net5614),
    .A1(net4791),
    .S(_04945_),
    .X(_00539_));
 sg13g2_mux2_1 _21769_ (.A0(net5608),
    .A1(net4454),
    .S(_04945_),
    .X(_00540_));
 sg13g2_mux2_1 _21770_ (.A0(net5583),
    .A1(net4652),
    .S(_04945_),
    .X(_00541_));
 sg13g2_mux2_1 _21771_ (.A0(net5577),
    .A1(net6661),
    .S(_04945_),
    .X(_00542_));
 sg13g2_mux2_1 _21772_ (.A0(net5643),
    .A1(net4677),
    .S(_04945_),
    .X(_00543_));
 sg13g2_nor2_2 _21773_ (.A(net5549),
    .B(_09397_),
    .Y(_04946_));
 sg13g2_nand3_1 _21774_ (.B(net5555),
    .C(_09261_),
    .A(net5281),
    .Y(_04947_));
 sg13g2_nor2_1 _21775_ (.A(net5248),
    .B(_04947_),
    .Y(_04948_));
 sg13g2_nor2_1 _21776_ (.A(net4253),
    .B(net5234),
    .Y(_04949_));
 sg13g2_a21oi_1 _21777_ (.A1(net5771),
    .A2(net5234),
    .Y(_00544_),
    .B1(_04949_));
 sg13g2_nor2_1 _21778_ (.A(net3063),
    .B(net5234),
    .Y(_04950_));
 sg13g2_a21oi_1 _21779_ (.A1(net5787),
    .A2(net5234),
    .Y(_00545_),
    .B1(_04950_));
 sg13g2_nor2_1 _21780_ (.A(net3781),
    .B(net5235),
    .Y(_04951_));
 sg13g2_a21oi_1 _21781_ (.A1(net5715),
    .A2(net5235),
    .Y(_00546_),
    .B1(_04951_));
 sg13g2_nor2_1 _21782_ (.A(net3972),
    .B(net5235),
    .Y(_04952_));
 sg13g2_a21oi_1 _21783_ (.A1(net5695),
    .A2(net5235),
    .Y(_00547_),
    .B1(_04952_));
 sg13g2_nor2_1 _21784_ (.A(net3626),
    .B(net5234),
    .Y(_04953_));
 sg13g2_a21oi_1 _21785_ (.A1(net5678),
    .A2(net5234),
    .Y(_00548_),
    .B1(_04953_));
 sg13g2_nor2_1 _21786_ (.A(net3365),
    .B(net5234),
    .Y(_04954_));
 sg13g2_a21oi_1 _21787_ (.A1(net5597),
    .A2(net5234),
    .Y(_00549_),
    .B1(_04954_));
 sg13g2_nor2_1 _21788_ (.A(net3089),
    .B(net5235),
    .Y(_04955_));
 sg13g2_a21oi_1 _21789_ (.A1(net5657),
    .A2(net5235),
    .Y(_00550_),
    .B1(_04955_));
 sg13g2_nor2_1 _21790_ (.A(net4323),
    .B(net5235),
    .Y(_04956_));
 sg13g2_a21oi_1 _21791_ (.A1(net5635),
    .A2(net5235),
    .Y(_00551_),
    .B1(_04956_));
 sg13g2_nor2_1 _21792_ (.A(net5236),
    .B(_04947_),
    .Y(_04957_));
 sg13g2_nor2_1 _21793_ (.A(net3148),
    .B(net5163),
    .Y(_04958_));
 sg13g2_a21oi_1 _21794_ (.A1(net5770),
    .A2(net5163),
    .Y(_00552_),
    .B1(_04958_));
 sg13g2_nor2_1 _21795_ (.A(net3371),
    .B(net5163),
    .Y(_04959_));
 sg13g2_a21oi_1 _21796_ (.A1(net5787),
    .A2(net5163),
    .Y(_00553_),
    .B1(_04959_));
 sg13g2_nor2_1 _21797_ (.A(net3232),
    .B(net5164),
    .Y(_04960_));
 sg13g2_a21oi_1 _21798_ (.A1(net5721),
    .A2(net5164),
    .Y(_00554_),
    .B1(_04960_));
 sg13g2_nor2_1 _21799_ (.A(net3436),
    .B(net5164),
    .Y(_04961_));
 sg13g2_a21oi_1 _21800_ (.A1(net5693),
    .A2(net5164),
    .Y(_00555_),
    .B1(_04961_));
 sg13g2_nor2_1 _21801_ (.A(net3062),
    .B(net5163),
    .Y(_04962_));
 sg13g2_a21oi_1 _21802_ (.A1(net5677),
    .A2(net5163),
    .Y(_00556_),
    .B1(_04962_));
 sg13g2_nor2_1 _21803_ (.A(net3209),
    .B(net5163),
    .Y(_04963_));
 sg13g2_a21oi_1 _21804_ (.A1(net5597),
    .A2(net5163),
    .Y(_00557_),
    .B1(_04963_));
 sg13g2_nor2_1 _21805_ (.A(net3971),
    .B(net5164),
    .Y(_04964_));
 sg13g2_a21oi_1 _21806_ (.A1(net5657),
    .A2(net5164),
    .Y(_00558_),
    .B1(_04964_));
 sg13g2_nor2_1 _21807_ (.A(net3663),
    .B(net5164),
    .Y(_04965_));
 sg13g2_a21oi_1 _21808_ (.A1(net5635),
    .A2(net5164),
    .Y(_00559_),
    .B1(_04965_));
 sg13g2_nor2_1 _21809_ (.A(net5258),
    .B(_04947_),
    .Y(_04966_));
 sg13g2_nor2_1 _21810_ (.A(net3651),
    .B(net5232),
    .Y(_04967_));
 sg13g2_a21oi_1 _21811_ (.A1(net5770),
    .A2(net5232),
    .Y(_00560_),
    .B1(_04967_));
 sg13g2_nor2_1 _21812_ (.A(net3861),
    .B(net5232),
    .Y(_04968_));
 sg13g2_a21oi_1 _21813_ (.A1(net5787),
    .A2(net5232),
    .Y(_00561_),
    .B1(_04968_));
 sg13g2_nor2_1 _21814_ (.A(net3388),
    .B(net5233),
    .Y(_04969_));
 sg13g2_a21oi_1 _21815_ (.A1(net5723),
    .A2(net5233),
    .Y(_00562_),
    .B1(_04969_));
 sg13g2_nor2_1 _21816_ (.A(net3428),
    .B(net5233),
    .Y(_04970_));
 sg13g2_a21oi_1 _21817_ (.A1(net5693),
    .A2(net5233),
    .Y(_00563_),
    .B1(_04970_));
 sg13g2_nor2_1 _21818_ (.A(net3421),
    .B(net5232),
    .Y(_04971_));
 sg13g2_a21oi_1 _21819_ (.A1(net5676),
    .A2(net5232),
    .Y(_00564_),
    .B1(_04971_));
 sg13g2_nor2_1 _21820_ (.A(net3493),
    .B(net5232),
    .Y(_04972_));
 sg13g2_a21oi_1 _21821_ (.A1(net5597),
    .A2(net5232),
    .Y(_00565_),
    .B1(_04972_));
 sg13g2_nor2_1 _21822_ (.A(net3431),
    .B(net5233),
    .Y(_04973_));
 sg13g2_a21oi_1 _21823_ (.A1(net5657),
    .A2(net5233),
    .Y(_00566_),
    .B1(_04973_));
 sg13g2_nor2_1 _21824_ (.A(net3331),
    .B(net5233),
    .Y(_04974_));
 sg13g2_a21oi_1 _21825_ (.A1(net5635),
    .A2(net5233),
    .Y(_00567_),
    .B1(_04974_));
 sg13g2_nand2_2 _21826_ (.Y(_04975_),
    .A(net5251),
    .B(_04946_));
 sg13g2_mux2_1 _21827_ (.A0(net5741),
    .A1(net4877),
    .S(_04975_),
    .X(_00568_));
 sg13g2_mux2_1 _21828_ (.A0(net5746),
    .A1(net6695),
    .S(_04975_),
    .X(_00569_));
 sg13g2_mux2_1 _21829_ (.A0(net5617),
    .A1(net4488),
    .S(_04975_),
    .X(_00570_));
 sg13g2_mux2_1 _21830_ (.A0(net5613),
    .A1(net6851),
    .S(_04975_),
    .X(_00571_));
 sg13g2_mux2_1 _21831_ (.A0(net5608),
    .A1(net6910),
    .S(_04975_),
    .X(_00572_));
 sg13g2_mux2_1 _21832_ (.A0(net5583),
    .A1(net4464),
    .S(_04975_),
    .X(_00573_));
 sg13g2_mux2_1 _21833_ (.A0(net5578),
    .A1(net4646),
    .S(_04975_),
    .X(_00574_));
 sg13g2_mux2_1 _21834_ (.A0(net5644),
    .A1(net4563),
    .S(_04975_),
    .X(_00575_));
 sg13g2_nor2_1 _21835_ (.A(net5239),
    .B(_04947_),
    .Y(_04976_));
 sg13g2_nor2_1 _21836_ (.A(net3157),
    .B(net5161),
    .Y(_04977_));
 sg13g2_a21oi_1 _21837_ (.A1(net5770),
    .A2(net5161),
    .Y(_00576_),
    .B1(_04977_));
 sg13g2_nor2_1 _21838_ (.A(net3359),
    .B(net5162),
    .Y(_04978_));
 sg13g2_a21oi_1 _21839_ (.A1(net5791),
    .A2(net5162),
    .Y(_00577_),
    .B1(_04978_));
 sg13g2_nor2_1 _21840_ (.A(net3432),
    .B(net5162),
    .Y(_04979_));
 sg13g2_a21oi_1 _21841_ (.A1(net5721),
    .A2(net5162),
    .Y(_00578_),
    .B1(_04979_));
 sg13g2_nor2_1 _21842_ (.A(net3084),
    .B(net5161),
    .Y(_04980_));
 sg13g2_a21oi_1 _21843_ (.A1(net5698),
    .A2(net5161),
    .Y(_00579_),
    .B1(_04980_));
 sg13g2_nor2_1 _21844_ (.A(net3155),
    .B(net5161),
    .Y(_04981_));
 sg13g2_a21oi_1 _21845_ (.A1(net5677),
    .A2(net5161),
    .Y(_00580_),
    .B1(_04981_));
 sg13g2_nor2_1 _21846_ (.A(net4465),
    .B(net5161),
    .Y(_04982_));
 sg13g2_a21oi_1 _21847_ (.A1(net5596),
    .A2(net5161),
    .Y(_00581_),
    .B1(_04982_));
 sg13g2_nor2_1 _21848_ (.A(net3134),
    .B(net5162),
    .Y(_04983_));
 sg13g2_a21oi_1 _21849_ (.A1(net5660),
    .A2(net5162),
    .Y(_00582_),
    .B1(_04983_));
 sg13g2_nor2_1 _21850_ (.A(net3611),
    .B(net5162),
    .Y(_04984_));
 sg13g2_a21oi_1 _21851_ (.A1(net5634),
    .A2(net5162),
    .Y(_00583_),
    .B1(_04984_));
 sg13g2_nor2_1 _21852_ (.A(_09331_),
    .B(net5259),
    .Y(_04985_));
 sg13g2_nor2_1 _21853_ (.A(net3440),
    .B(net5063),
    .Y(_04986_));
 sg13g2_a21oi_1 _21854_ (.A1(net5761),
    .A2(net5063),
    .Y(_00584_),
    .B1(_04986_));
 sg13g2_nor2_1 _21855_ (.A(net3343),
    .B(net5063),
    .Y(_04987_));
 sg13g2_a21oi_1 _21856_ (.A1(net5781),
    .A2(net5063),
    .Y(_00585_),
    .B1(_04987_));
 sg13g2_nor2_1 _21857_ (.A(net3382),
    .B(net5063),
    .Y(_04988_));
 sg13g2_a21oi_1 _21858_ (.A1(net5711),
    .A2(net5063),
    .Y(_00586_),
    .B1(_04988_));
 sg13g2_nor2_1 _21859_ (.A(net4376),
    .B(net5064),
    .Y(_04989_));
 sg13g2_a21oi_1 _21860_ (.A1(net5686),
    .A2(net5064),
    .Y(_00587_),
    .B1(_04989_));
 sg13g2_nor2_1 _21861_ (.A(net3525),
    .B(net5064),
    .Y(_04990_));
 sg13g2_a21oi_1 _21862_ (.A1(net5667),
    .A2(_04985_),
    .Y(_00588_),
    .B1(_04990_));
 sg13g2_nor2_1 _21863_ (.A(net3496),
    .B(net5064),
    .Y(_04991_));
 sg13g2_a21oi_1 _21864_ (.A1(net5587),
    .A2(net5064),
    .Y(_00589_),
    .B1(_04991_));
 sg13g2_nor2_1 _21865_ (.A(net4263),
    .B(net5064),
    .Y(_04992_));
 sg13g2_a21oi_1 _21866_ (.A1(net5649),
    .A2(net5064),
    .Y(_00590_),
    .B1(_04992_));
 sg13g2_nor2_1 _21867_ (.A(net3655),
    .B(net5063),
    .Y(_04993_));
 sg13g2_a21oi_1 _21868_ (.A1(net5624),
    .A2(net5063),
    .Y(_00591_),
    .B1(_04993_));
 sg13g2_nor2_1 _21869_ (.A(net5256),
    .B(_04947_),
    .Y(_04994_));
 sg13g2_nor2_1 _21870_ (.A(net4181),
    .B(net5230),
    .Y(_04995_));
 sg13g2_a21oi_1 _21871_ (.A1(net5770),
    .A2(net5230),
    .Y(_00592_),
    .B1(_04995_));
 sg13g2_nor2_1 _21872_ (.A(net4294),
    .B(net5231),
    .Y(_04996_));
 sg13g2_a21oi_1 _21873_ (.A1(net5791),
    .A2(net5231),
    .Y(_00593_),
    .B1(_04996_));
 sg13g2_nor2_1 _21874_ (.A(net4059),
    .B(net5231),
    .Y(_04997_));
 sg13g2_a21oi_1 _21875_ (.A1(net5721),
    .A2(net5231),
    .Y(_00594_),
    .B1(_04997_));
 sg13g2_nor2_1 _21876_ (.A(net4064),
    .B(net5230),
    .Y(_04998_));
 sg13g2_a21oi_1 _21877_ (.A1(net5698),
    .A2(net5230),
    .Y(_00595_),
    .B1(_04998_));
 sg13g2_nor2_1 _21878_ (.A(net3574),
    .B(net5230),
    .Y(_04999_));
 sg13g2_a21oi_1 _21879_ (.A1(net5677),
    .A2(net5230),
    .Y(_00596_),
    .B1(_04999_));
 sg13g2_nor2_1 _21880_ (.A(net3384),
    .B(net5230),
    .Y(_05000_));
 sg13g2_a21oi_1 _21881_ (.A1(net5596),
    .A2(net5230),
    .Y(_00597_),
    .B1(_05000_));
 sg13g2_nor2_1 _21882_ (.A(net4407),
    .B(net5231),
    .Y(_05001_));
 sg13g2_a21oi_1 _21883_ (.A1(net5660),
    .A2(net5231),
    .Y(_00598_),
    .B1(_05001_));
 sg13g2_nor2_1 _21884_ (.A(net4238),
    .B(net5231),
    .Y(_05002_));
 sg13g2_a21oi_1 _21885_ (.A1(net5634),
    .A2(net5231),
    .Y(_00599_),
    .B1(_05002_));
 sg13g2_nand2_2 _21886_ (.Y(_05003_),
    .A(net5253),
    .B(_04946_));
 sg13g2_mux2_1 _21887_ (.A0(net5741),
    .A1(net4910),
    .S(_05003_),
    .X(_00600_));
 sg13g2_mux2_1 _21888_ (.A0(net5746),
    .A1(net4741),
    .S(_05003_),
    .X(_00601_));
 sg13g2_mux2_1 _21889_ (.A0(net5617),
    .A1(net6999),
    .S(_05003_),
    .X(_00602_));
 sg13g2_mux2_1 _21890_ (.A0(net5614),
    .A1(net4820),
    .S(_05003_),
    .X(_00603_));
 sg13g2_mux2_1 _21891_ (.A0(net5608),
    .A1(net6692),
    .S(_05003_),
    .X(_00604_));
 sg13g2_mux2_1 _21892_ (.A0(net5583),
    .A1(net4814),
    .S(_05003_),
    .X(_00605_));
 sg13g2_mux2_1 _21893_ (.A0(net5577),
    .A1(net6651),
    .S(_05003_),
    .X(_00606_));
 sg13g2_mux2_1 _21894_ (.A0(net5643),
    .A1(net7043),
    .S(_05003_),
    .X(_00607_));
 sg13g2_nor2_2 _21895_ (.A(_09361_),
    .B(_03123_),
    .Y(_05004_));
 sg13g2_nand3_1 _21896_ (.B(net5551),
    .C(_09261_),
    .A(net5276),
    .Y(_05005_));
 sg13g2_nor2_1 _21897_ (.A(net5248),
    .B(_05005_),
    .Y(_05006_));
 sg13g2_nor2_1 _21898_ (.A(net3110),
    .B(net5229),
    .Y(_05007_));
 sg13g2_a21oi_1 _21899_ (.A1(net5765),
    .A2(net5229),
    .Y(_00608_),
    .B1(_05007_));
 sg13g2_nor2_1 _21900_ (.A(net4424),
    .B(net5228),
    .Y(_05008_));
 sg13g2_a21oi_1 _21901_ (.A1(net5786),
    .A2(net5228),
    .Y(_00609_),
    .B1(_05008_));
 sg13g2_nor2_1 _21902_ (.A(net3064),
    .B(net5229),
    .Y(_05009_));
 sg13g2_a21oi_1 _21903_ (.A1(net5716),
    .A2(net5229),
    .Y(_00610_),
    .B1(_05009_));
 sg13g2_nor2_1 _21904_ (.A(net3872),
    .B(net5229),
    .Y(_05010_));
 sg13g2_a21oi_1 _21905_ (.A1(net5693),
    .A2(net5229),
    .Y(_00611_),
    .B1(_05010_));
 sg13g2_nor2_1 _21906_ (.A(net4070),
    .B(net5229),
    .Y(_05011_));
 sg13g2_a21oi_1 _21907_ (.A1(net5673),
    .A2(net5229),
    .Y(_00612_),
    .B1(_05011_));
 sg13g2_nor2_1 _21908_ (.A(net4252),
    .B(net5228),
    .Y(_05012_));
 sg13g2_a21oi_1 _21909_ (.A1(net5589),
    .A2(net5228),
    .Y(_00613_),
    .B1(_05012_));
 sg13g2_nor2_1 _21910_ (.A(net3169),
    .B(net5228),
    .Y(_05013_));
 sg13g2_a21oi_1 _21911_ (.A1(net5653),
    .A2(net5228),
    .Y(_00614_),
    .B1(_05013_));
 sg13g2_nor2_1 _21912_ (.A(net3407),
    .B(net5228),
    .Y(_05014_));
 sg13g2_a21oi_1 _21913_ (.A1(net5627),
    .A2(net5228),
    .Y(_00615_),
    .B1(_05014_));
 sg13g2_nor2_1 _21914_ (.A(net5236),
    .B(_05005_),
    .Y(_05015_));
 sg13g2_nor2_1 _21915_ (.A(net4062),
    .B(net5160),
    .Y(_05016_));
 sg13g2_a21oi_1 _21916_ (.A1(net5766),
    .A2(net5160),
    .Y(_00616_),
    .B1(_05016_));
 sg13g2_nor2_1 _21917_ (.A(net3271),
    .B(net5159),
    .Y(_05017_));
 sg13g2_a21oi_1 _21918_ (.A1(net5784),
    .A2(net5159),
    .Y(_00617_),
    .B1(_05017_));
 sg13g2_nor2_1 _21919_ (.A(net3920),
    .B(net5160),
    .Y(_05018_));
 sg13g2_a21oi_1 _21920_ (.A1(net5716),
    .A2(net5160),
    .Y(_00618_),
    .B1(_05018_));
 sg13g2_nor2_1 _21921_ (.A(net3750),
    .B(net5160),
    .Y(_05019_));
 sg13g2_a21oi_1 _21922_ (.A1(net5692),
    .A2(net5160),
    .Y(_00619_),
    .B1(_05019_));
 sg13g2_nor2_1 _21923_ (.A(net3286),
    .B(net5160),
    .Y(_05020_));
 sg13g2_a21oi_1 _21924_ (.A1(net5673),
    .A2(net5160),
    .Y(_00620_),
    .B1(_05020_));
 sg13g2_nor2_1 _21925_ (.A(net4195),
    .B(net5159),
    .Y(_05021_));
 sg13g2_a21oi_1 _21926_ (.A1(net5589),
    .A2(net5159),
    .Y(_00621_),
    .B1(_05021_));
 sg13g2_nor2_1 _21927_ (.A(net3272),
    .B(net5159),
    .Y(_05022_));
 sg13g2_a21oi_1 _21928_ (.A1(net5653),
    .A2(net5159),
    .Y(_00622_),
    .B1(_05022_));
 sg13g2_nor2_1 _21929_ (.A(net3273),
    .B(net5159),
    .Y(_05023_));
 sg13g2_a21oi_1 _21930_ (.A1(net5627),
    .A2(net5159),
    .Y(_00623_),
    .B1(_05023_));
 sg13g2_nor2_1 _21931_ (.A(net5258),
    .B(_05005_),
    .Y(_05024_));
 sg13g2_nor2_1 _21932_ (.A(net4216),
    .B(net5227),
    .Y(_05025_));
 sg13g2_a21oi_1 _21933_ (.A1(net5766),
    .A2(net5227),
    .Y(_00624_),
    .B1(_05025_));
 sg13g2_nor2_1 _21934_ (.A(net3434),
    .B(net5226),
    .Y(_05026_));
 sg13g2_a21oi_1 _21935_ (.A1(net5784),
    .A2(net5226),
    .Y(_00625_),
    .B1(_05026_));
 sg13g2_nor2_1 _21936_ (.A(net3366),
    .B(net5227),
    .Y(_05027_));
 sg13g2_a21oi_1 _21937_ (.A1(net5716),
    .A2(net5227),
    .Y(_00626_),
    .B1(_05027_));
 sg13g2_nor2_1 _21938_ (.A(net3535),
    .B(net5227),
    .Y(_05028_));
 sg13g2_a21oi_1 _21939_ (.A1(net5692),
    .A2(net5227),
    .Y(_00627_),
    .B1(_05028_));
 sg13g2_nor2_1 _21940_ (.A(net3274),
    .B(net5227),
    .Y(_05029_));
 sg13g2_a21oi_1 _21941_ (.A1(net5673),
    .A2(net5227),
    .Y(_00628_),
    .B1(_05029_));
 sg13g2_nor2_1 _21942_ (.A(net4188),
    .B(net5226),
    .Y(_05030_));
 sg13g2_a21oi_1 _21943_ (.A1(net5589),
    .A2(net5226),
    .Y(_00629_),
    .B1(_05030_));
 sg13g2_nor2_1 _21944_ (.A(net4391),
    .B(net5226),
    .Y(_05031_));
 sg13g2_a21oi_1 _21945_ (.A1(net5653),
    .A2(net5226),
    .Y(_00630_),
    .B1(_05031_));
 sg13g2_nor2_1 _21946_ (.A(net3317),
    .B(net5226),
    .Y(_05032_));
 sg13g2_a21oi_1 _21947_ (.A1(net5627),
    .A2(net5226),
    .Y(_00631_),
    .B1(_05032_));
 sg13g2_nand2_2 _21948_ (.Y(_05033_),
    .A(net5251),
    .B(_05004_));
 sg13g2_mux2_1 _21949_ (.A0(net5739),
    .A1(net4690),
    .S(_05033_),
    .X(_00632_));
 sg13g2_mux2_1 _21950_ (.A0(net5744),
    .A1(net6807),
    .S(_05033_),
    .X(_00633_));
 sg13g2_mux2_1 _21951_ (.A0(net5617),
    .A1(net6644),
    .S(_05033_),
    .X(_00634_));
 sg13g2_mux2_1 _21952_ (.A0(net5614),
    .A1(net6749),
    .S(_05033_),
    .X(_00635_));
 sg13g2_mux2_1 _21953_ (.A0(net5606),
    .A1(net4635),
    .S(_05033_),
    .X(_00636_));
 sg13g2_mux2_1 _21954_ (.A0(net5581),
    .A1(net4835),
    .S(_05033_),
    .X(_00637_));
 sg13g2_mux2_1 _21955_ (.A0(net5576),
    .A1(net4711),
    .S(_05033_),
    .X(_00638_));
 sg13g2_mux2_1 _21956_ (.A0(net5642),
    .A1(net7016),
    .S(_05033_),
    .X(_00639_));
 sg13g2_nor2_1 _21957_ (.A(net5239),
    .B(_05005_),
    .Y(_05034_));
 sg13g2_nor2_1 _21958_ (.A(net3411),
    .B(net5158),
    .Y(_05035_));
 sg13g2_a21oi_1 _21959_ (.A1(net5766),
    .A2(net5158),
    .Y(_00640_),
    .B1(_05035_));
 sg13g2_nor2_1 _21960_ (.A(net3531),
    .B(net5158),
    .Y(_05036_));
 sg13g2_a21oi_1 _21961_ (.A1(net5791),
    .A2(net5158),
    .Y(_00641_),
    .B1(_05036_));
 sg13g2_nor2_1 _21962_ (.A(net3375),
    .B(net5158),
    .Y(_05037_));
 sg13g2_a21oi_1 _21963_ (.A1(net5716),
    .A2(net5158),
    .Y(_00642_),
    .B1(_05037_));
 sg13g2_nor2_1 _21964_ (.A(net3711),
    .B(net5157),
    .Y(_05038_));
 sg13g2_a21oi_1 _21965_ (.A1(net5692),
    .A2(net5157),
    .Y(_00643_),
    .B1(_05038_));
 sg13g2_nor2_1 _21966_ (.A(net3054),
    .B(net5158),
    .Y(_05039_));
 sg13g2_a21oi_1 _21967_ (.A1(net5676),
    .A2(net5158),
    .Y(_00644_),
    .B1(_05039_));
 sg13g2_nor2_1 _21968_ (.A(net4404),
    .B(net5157),
    .Y(_05040_));
 sg13g2_a21oi_1 _21969_ (.A1(net5590),
    .A2(net5157),
    .Y(_00645_),
    .B1(_05040_));
 sg13g2_nor2_1 _21970_ (.A(net3047),
    .B(net5157),
    .Y(_05041_));
 sg13g2_a21oi_1 _21971_ (.A1(net5652),
    .A2(net5157),
    .Y(_00646_),
    .B1(_05041_));
 sg13g2_nor2_1 _21972_ (.A(net3615),
    .B(net5157),
    .Y(_05042_));
 sg13g2_a21oi_1 _21973_ (.A1(net5626),
    .A2(net5157),
    .Y(_00647_),
    .B1(_05042_));
 sg13g2_nor2_1 _21974_ (.A(net5254),
    .B(_05005_),
    .Y(_05043_));
 sg13g2_nor2_1 _21975_ (.A(net3715),
    .B(net5225),
    .Y(_05044_));
 sg13g2_a21oi_1 _21976_ (.A1(net5765),
    .A2(net5225),
    .Y(_00648_),
    .B1(_05044_));
 sg13g2_nor2_1 _21977_ (.A(net3374),
    .B(net5225),
    .Y(_05045_));
 sg13g2_a21oi_1 _21978_ (.A1(net5787),
    .A2(net5225),
    .Y(_00649_),
    .B1(_05045_));
 sg13g2_nor2_1 _21979_ (.A(net3055),
    .B(net5225),
    .Y(_05046_));
 sg13g2_a21oi_1 _21980_ (.A1(net5715),
    .A2(net5225),
    .Y(_00650_),
    .B1(_05046_));
 sg13g2_nor2_1 _21981_ (.A(net4328),
    .B(net5224),
    .Y(_05047_));
 sg13g2_a21oi_1 _21982_ (.A1(net5692),
    .A2(net5224),
    .Y(_00651_),
    .B1(_05047_));
 sg13g2_nor2_1 _21983_ (.A(net3460),
    .B(net5225),
    .Y(_05048_));
 sg13g2_a21oi_1 _21984_ (.A1(net5676),
    .A2(net5225),
    .Y(_00652_),
    .B1(_05048_));
 sg13g2_nor2_1 _21985_ (.A(net3759),
    .B(net5224),
    .Y(_05049_));
 sg13g2_a21oi_1 _21986_ (.A1(net5589),
    .A2(net5224),
    .Y(_00653_),
    .B1(_05049_));
 sg13g2_nor2_1 _21987_ (.A(net3990),
    .B(net5224),
    .Y(_05050_));
 sg13g2_a21oi_1 _21988_ (.A1(net5652),
    .A2(net5224),
    .Y(_00654_),
    .B1(_05050_));
 sg13g2_nor2_1 _21989_ (.A(net3862),
    .B(net5224),
    .Y(_05051_));
 sg13g2_a21oi_1 _21990_ (.A1(net5626),
    .A2(net5224),
    .Y(_00655_),
    .B1(_05051_));
 sg13g2_nor2_1 _21991_ (.A(net5256),
    .B(_05005_),
    .Y(_05052_));
 sg13g2_nor2_1 _21992_ (.A(net3558),
    .B(net5223),
    .Y(_05053_));
 sg13g2_a21oi_1 _21993_ (.A1(net5766),
    .A2(net5223),
    .Y(_00656_),
    .B1(_05053_));
 sg13g2_nor2_1 _21994_ (.A(net3410),
    .B(net5221),
    .Y(_05054_));
 sg13g2_a21oi_1 _21995_ (.A1(net5787),
    .A2(net5221),
    .Y(_00657_),
    .B1(_05054_));
 sg13g2_nor2_1 _21996_ (.A(net4413),
    .B(net5222),
    .Y(_05055_));
 sg13g2_a21oi_1 _21997_ (.A1(net5715),
    .A2(net5222),
    .Y(_00658_),
    .B1(_05055_));
 sg13g2_nor2_1 _21998_ (.A(net4284),
    .B(net5221),
    .Y(_05056_));
 sg13g2_a21oi_1 _21999_ (.A1(net5692),
    .A2(net5221),
    .Y(_00659_),
    .B1(_05056_));
 sg13g2_nor2_1 _22000_ (.A(net3183),
    .B(net5222),
    .Y(_05057_));
 sg13g2_a21oi_1 _22001_ (.A1(net5676),
    .A2(net5222),
    .Y(_00660_),
    .B1(_05057_));
 sg13g2_nor2_1 _22002_ (.A(net3947),
    .B(net5223),
    .Y(_05058_));
 sg13g2_a21oi_1 _22003_ (.A1(net5589),
    .A2(net5223),
    .Y(_00661_),
    .B1(_05058_));
 sg13g2_nor2_1 _22004_ (.A(net3486),
    .B(net5221),
    .Y(_05059_));
 sg13g2_a21oi_1 _22005_ (.A1(net5652),
    .A2(net5221),
    .Y(_00662_),
    .B1(_05059_));
 sg13g2_nor2_1 _22006_ (.A(net3095),
    .B(net5221),
    .Y(_05060_));
 sg13g2_a21oi_1 _22007_ (.A1(net5626),
    .A2(net5221),
    .Y(_00663_),
    .B1(_05060_));
 sg13g2_nand3_1 _22008_ (.B(_09329_),
    .C(net5250),
    .A(net5556),
    .Y(_05061_));
 sg13g2_mux2_1 _22009_ (.A0(net5740),
    .A1(net7070),
    .S(_05061_),
    .X(_00664_));
 sg13g2_mux2_1 _22010_ (.A0(net5745),
    .A1(net6767),
    .S(_05061_),
    .X(_00665_));
 sg13g2_mux2_1 _22011_ (.A0(net5616),
    .A1(net4569),
    .S(_05061_),
    .X(_00666_));
 sg13g2_mux2_1 _22012_ (.A0(net5611),
    .A1(net6963),
    .S(_05061_),
    .X(_00667_));
 sg13g2_mux2_1 _22013_ (.A0(net5607),
    .A1(net7030),
    .S(_05061_),
    .X(_00668_));
 sg13g2_mux2_1 _22014_ (.A0(net5580),
    .A1(net6825),
    .S(_05061_),
    .X(_00669_));
 sg13g2_mux2_1 _22015_ (.A0(net5575),
    .A1(net4921),
    .S(_05061_),
    .X(_00670_));
 sg13g2_mux2_1 _22016_ (.A0(net5641),
    .A1(net4494),
    .S(_05061_),
    .X(_00671_));
 sg13g2_nor2_1 _22017_ (.A(_09265_),
    .B(net5248),
    .Y(_05062_));
 sg13g2_nor2_1 _22018_ (.A(net3101),
    .B(net5155),
    .Y(_05063_));
 sg13g2_a21oi_1 _22019_ (.A1(net5765),
    .A2(_05062_),
    .Y(_00672_),
    .B1(_05063_));
 sg13g2_nor2_1 _22020_ (.A(net4164),
    .B(net5156),
    .Y(_05064_));
 sg13g2_a21oi_1 _22021_ (.A1(net5786),
    .A2(net5156),
    .Y(_00673_),
    .B1(_05064_));
 sg13g2_nor2_1 _22022_ (.A(net3162),
    .B(net5155),
    .Y(_05065_));
 sg13g2_a21oi_1 _22023_ (.A1(net5715),
    .A2(net5155),
    .Y(_00674_),
    .B1(_05065_));
 sg13g2_nor2_1 _22024_ (.A(net3031),
    .B(net5155),
    .Y(_05066_));
 sg13g2_a21oi_1 _22025_ (.A1(net5693),
    .A2(net5155),
    .Y(_00675_),
    .B1(_05066_));
 sg13g2_nor2_1 _22026_ (.A(net3186),
    .B(net5155),
    .Y(_05067_));
 sg13g2_a21oi_1 _22027_ (.A1(net5679),
    .A2(net5156),
    .Y(_00676_),
    .B1(_05067_));
 sg13g2_nor2_1 _22028_ (.A(net3791),
    .B(net5155),
    .Y(_05068_));
 sg13g2_a21oi_1 _22029_ (.A1(net5589),
    .A2(net5155),
    .Y(_00677_),
    .B1(_05068_));
 sg13g2_nor2_1 _22030_ (.A(net3393),
    .B(net5156),
    .Y(_05069_));
 sg13g2_a21oi_1 _22031_ (.A1(net5653),
    .A2(net5156),
    .Y(_00678_),
    .B1(_05069_));
 sg13g2_nor2_1 _22032_ (.A(net3788),
    .B(net5156),
    .Y(_05070_));
 sg13g2_a21oi_1 _22033_ (.A1(net5627),
    .A2(net5156),
    .Y(_00679_),
    .B1(_05070_));
 sg13g2_nor2_1 _22034_ (.A(_09265_),
    .B(net5236),
    .Y(_05071_));
 sg13g2_nor2_1 _22035_ (.A(net3899),
    .B(net5154),
    .Y(_05072_));
 sg13g2_a21oi_1 _22036_ (.A1(net5765),
    .A2(net5154),
    .Y(_00680_),
    .B1(_05072_));
 sg13g2_nor2_1 _22037_ (.A(net3170),
    .B(net5153),
    .Y(_05073_));
 sg13g2_a21oi_1 _22038_ (.A1(net5785),
    .A2(net5153),
    .Y(_00681_),
    .B1(_05073_));
 sg13g2_nor2_1 _22039_ (.A(net3473),
    .B(net5154),
    .Y(_05074_));
 sg13g2_a21oi_1 _22040_ (.A1(net5716),
    .A2(net5154),
    .Y(_00682_),
    .B1(_05074_));
 sg13g2_nor2_1 _22041_ (.A(net3882),
    .B(net5154),
    .Y(_05075_));
 sg13g2_a21oi_1 _22042_ (.A1(net5693),
    .A2(net5154),
    .Y(_00683_),
    .B1(_05075_));
 sg13g2_nor2_1 _22043_ (.A(net3413),
    .B(net5154),
    .Y(_05076_));
 sg13g2_a21oi_1 _22044_ (.A1(net5678),
    .A2(net5154),
    .Y(_00684_),
    .B1(_05076_));
 sg13g2_nor2_1 _22045_ (.A(net4319),
    .B(net5153),
    .Y(_05077_));
 sg13g2_a21oi_1 _22046_ (.A1(net5589),
    .A2(net5153),
    .Y(_00685_),
    .B1(_05077_));
 sg13g2_nor2_1 _22047_ (.A(net3143),
    .B(net5153),
    .Y(_05078_));
 sg13g2_a21oi_1 _22048_ (.A1(net5653),
    .A2(net5153),
    .Y(_00686_),
    .B1(_05078_));
 sg13g2_nor2_1 _22049_ (.A(net3396),
    .B(net5153),
    .Y(_05079_));
 sg13g2_a21oi_1 _22050_ (.A1(net5627),
    .A2(net5153),
    .Y(_00687_),
    .B1(_05079_));
 sg13g2_nor2_1 _22051_ (.A(_09265_),
    .B(net5258),
    .Y(_05080_));
 sg13g2_nor2_1 _22052_ (.A(net4186),
    .B(net5152),
    .Y(_05081_));
 sg13g2_a21oi_1 _22053_ (.A1(net5765),
    .A2(net5152),
    .Y(_00688_),
    .B1(_05081_));
 sg13g2_nor2_1 _22054_ (.A(net4279),
    .B(net5151),
    .Y(_05082_));
 sg13g2_a21oi_1 _22055_ (.A1(net5785),
    .A2(net5151),
    .Y(_00689_),
    .B1(_05082_));
 sg13g2_nor2_1 _22056_ (.A(net4378),
    .B(net5152),
    .Y(_05083_));
 sg13g2_a21oi_1 _22057_ (.A1(net5715),
    .A2(net5152),
    .Y(_00690_),
    .B1(_05083_));
 sg13g2_nor2_1 _22058_ (.A(net3419),
    .B(net5152),
    .Y(_05084_));
 sg13g2_a21oi_1 _22059_ (.A1(net5693),
    .A2(net5152),
    .Y(_00691_),
    .B1(_05084_));
 sg13g2_nor2_1 _22060_ (.A(net3891),
    .B(net5152),
    .Y(_05085_));
 sg13g2_a21oi_1 _22061_ (.A1(net5678),
    .A2(net5152),
    .Y(_00692_),
    .B1(_05085_));
 sg13g2_nor2_1 _22062_ (.A(net3462),
    .B(net5151),
    .Y(_05086_));
 sg13g2_a21oi_1 _22063_ (.A1(net5589),
    .A2(net5151),
    .Y(_00693_),
    .B1(_05086_));
 sg13g2_nor2_1 _22064_ (.A(net3217),
    .B(net5151),
    .Y(_05087_));
 sg13g2_a21oi_1 _22065_ (.A1(net5653),
    .A2(net5151),
    .Y(_00694_),
    .B1(_05087_));
 sg13g2_nor2_1 _22066_ (.A(net4301),
    .B(net5151),
    .Y(_05088_));
 sg13g2_a21oi_1 _22067_ (.A1(net5627),
    .A2(net5151),
    .Y(_00695_),
    .B1(_05088_));
 sg13g2_nand2_2 _22068_ (.Y(_05089_),
    .A(_09264_),
    .B(net5250));
 sg13g2_mux2_1 _22069_ (.A0(_09199_),
    .A1(net7216),
    .S(_05089_),
    .X(_00696_));
 sg13g2_mux2_1 _22070_ (.A0(net5744),
    .A1(net7085),
    .S(_05089_),
    .X(_00697_));
 sg13g2_mux2_1 _22071_ (.A0(net5618),
    .A1(net7099),
    .S(_05089_),
    .X(_00698_));
 sg13g2_mux2_1 _22072_ (.A0(net5614),
    .A1(net4527),
    .S(_05089_),
    .X(_00699_));
 sg13g2_mux2_1 _22073_ (.A0(net5608),
    .A1(net6619),
    .S(_05089_),
    .X(_00700_));
 sg13g2_mux2_1 _22074_ (.A0(net5581),
    .A1(net6662),
    .S(_05089_),
    .X(_00701_));
 sg13g2_mux2_1 _22075_ (.A0(net5578),
    .A1(net6900),
    .S(_05089_),
    .X(_00702_));
 sg13g2_mux2_1 _22076_ (.A0(net5642),
    .A1(net6970),
    .S(_05089_),
    .X(_00703_));
 sg13g2_nor2_1 _22077_ (.A(_09265_),
    .B(net5239),
    .Y(_05090_));
 sg13g2_nor2_1 _22078_ (.A(net3086),
    .B(net5150),
    .Y(_05091_));
 sg13g2_a21oi_1 _22079_ (.A1(net5765),
    .A2(net5150),
    .Y(_00704_),
    .B1(_05091_));
 sg13g2_nor2_1 _22080_ (.A(net3562),
    .B(net5149),
    .Y(_05092_));
 sg13g2_a21oi_1 _22081_ (.A1(net5787),
    .A2(net5149),
    .Y(_00705_),
    .B1(_05092_));
 sg13g2_nor2_1 _22082_ (.A(net4312),
    .B(net5150),
    .Y(_05093_));
 sg13g2_a21oi_1 _22083_ (.A1(net5715),
    .A2(net5150),
    .Y(_00706_),
    .B1(_05093_));
 sg13g2_nor2_1 _22084_ (.A(net3283),
    .B(net5150),
    .Y(_05094_));
 sg13g2_a21oi_1 _22085_ (.A1(net5692),
    .A2(net5150),
    .Y(_00707_),
    .B1(_05094_));
 sg13g2_nor2_1 _22086_ (.A(net3194),
    .B(net5150),
    .Y(_05095_));
 sg13g2_a21oi_1 _22087_ (.A1(net5676),
    .A2(net5150),
    .Y(_00708_),
    .B1(_05095_));
 sg13g2_nor2_1 _22088_ (.A(net4122),
    .B(net5149),
    .Y(_05096_));
 sg13g2_a21oi_1 _22089_ (.A1(net5590),
    .A2(net5149),
    .Y(_00709_),
    .B1(_05096_));
 sg13g2_nor2_1 _22090_ (.A(net3856),
    .B(net5149),
    .Y(_05097_));
 sg13g2_a21oi_1 _22091_ (.A1(net5652),
    .A2(net5149),
    .Y(_00710_),
    .B1(_05097_));
 sg13g2_nor2_1 _22092_ (.A(net4010),
    .B(net5149),
    .Y(_05098_));
 sg13g2_a21oi_1 _22093_ (.A1(net5626),
    .A2(net5149),
    .Y(_00711_),
    .B1(_05098_));
 sg13g2_nor2_1 _22094_ (.A(_09265_),
    .B(net5254),
    .Y(_05099_));
 sg13g2_nor2_1 _22095_ (.A(net3905),
    .B(net5148),
    .Y(_05100_));
 sg13g2_a21oi_1 _22096_ (.A1(net5765),
    .A2(net5148),
    .Y(_00712_),
    .B1(_05100_));
 sg13g2_nor2_1 _22097_ (.A(net3779),
    .B(net5147),
    .Y(_05101_));
 sg13g2_a21oi_1 _22098_ (.A1(net5790),
    .A2(net5147),
    .Y(_00713_),
    .B1(_05101_));
 sg13g2_nor2_1 _22099_ (.A(net3129),
    .B(net5148),
    .Y(_05102_));
 sg13g2_a21oi_1 _22100_ (.A1(net5715),
    .A2(net5148),
    .Y(_00714_),
    .B1(_05102_));
 sg13g2_nor2_1 _22101_ (.A(net3093),
    .B(net5148),
    .Y(_05103_));
 sg13g2_a21oi_1 _22102_ (.A1(net5692),
    .A2(net5148),
    .Y(_00715_),
    .B1(_05103_));
 sg13g2_nor2_1 _22103_ (.A(net4208),
    .B(net5148),
    .Y(_05104_));
 sg13g2_a21oi_1 _22104_ (.A1(net5676),
    .A2(net5148),
    .Y(_00716_),
    .B1(_05104_));
 sg13g2_nor2_1 _22105_ (.A(net3332),
    .B(net5147),
    .Y(_05105_));
 sg13g2_a21oi_1 _22106_ (.A1(net5590),
    .A2(net5147),
    .Y(_00717_),
    .B1(_05105_));
 sg13g2_nor2_1 _22107_ (.A(net4002),
    .B(net5147),
    .Y(_05106_));
 sg13g2_a21oi_1 _22108_ (.A1(net5652),
    .A2(net5147),
    .Y(_00718_),
    .B1(_05106_));
 sg13g2_nor2_1 _22109_ (.A(net3052),
    .B(net5147),
    .Y(_05107_));
 sg13g2_a21oi_1 _22110_ (.A1(net5626),
    .A2(net5147),
    .Y(_00719_),
    .B1(_05107_));
 sg13g2_nor2_1 _22111_ (.A(_09265_),
    .B(net5256),
    .Y(_05108_));
 sg13g2_nor2_1 _22112_ (.A(net3284),
    .B(net5146),
    .Y(_05109_));
 sg13g2_a21oi_1 _22113_ (.A1(net5765),
    .A2(net5146),
    .Y(_00720_),
    .B1(_05109_));
 sg13g2_nor2_1 _22114_ (.A(net3354),
    .B(net5145),
    .Y(_05110_));
 sg13g2_a21oi_1 _22115_ (.A1(net5787),
    .A2(net5145),
    .Y(_00721_),
    .B1(_05110_));
 sg13g2_nor2_1 _22116_ (.A(net3900),
    .B(net5146),
    .Y(_05111_));
 sg13g2_a21oi_1 _22117_ (.A1(net5715),
    .A2(net5146),
    .Y(_00722_),
    .B1(_05111_));
 sg13g2_nor2_1 _22118_ (.A(net3266),
    .B(net5146),
    .Y(_05112_));
 sg13g2_a21oi_1 _22119_ (.A1(net5692),
    .A2(net5146),
    .Y(_00723_),
    .B1(_05112_));
 sg13g2_nor2_1 _22120_ (.A(net3477),
    .B(net5146),
    .Y(_05113_));
 sg13g2_a21oi_1 _22121_ (.A1(net5676),
    .A2(net5146),
    .Y(_00724_),
    .B1(_05113_));
 sg13g2_nor2_1 _22122_ (.A(net4209),
    .B(net5145),
    .Y(_05114_));
 sg13g2_a21oi_1 _22123_ (.A1(net5590),
    .A2(net5145),
    .Y(_00725_),
    .B1(_05114_));
 sg13g2_nor2_1 _22124_ (.A(net4310),
    .B(net5145),
    .Y(_05115_));
 sg13g2_a21oi_1 _22125_ (.A1(net5652),
    .A2(net5145),
    .Y(_00726_),
    .B1(_05115_));
 sg13g2_nor2_1 _22126_ (.A(net3171),
    .B(net5145),
    .Y(_05116_));
 sg13g2_a21oi_1 _22127_ (.A1(net5626),
    .A2(net5145),
    .Y(_00727_),
    .B1(_05116_));
 sg13g2_nor2_1 _22128_ (.A(_03021_),
    .B(net5239),
    .Y(_05117_));
 sg13g2_nor2_1 _22129_ (.A(net4379),
    .B(net5143),
    .Y(_05118_));
 sg13g2_a21oi_1 _22130_ (.A1(net5774),
    .A2(net5143),
    .Y(_00728_),
    .B1(_05118_));
 sg13g2_nor2_1 _22131_ (.A(net4072),
    .B(net5143),
    .Y(_05119_));
 sg13g2_a21oi_1 _22132_ (.A1(net5794),
    .A2(net5143),
    .Y(_00729_),
    .B1(_05119_));
 sg13g2_nor2_1 _22133_ (.A(net4283),
    .B(net5143),
    .Y(_05120_));
 sg13g2_a21oi_1 _22134_ (.A1(net5724),
    .A2(net5143),
    .Y(_00730_),
    .B1(_05120_));
 sg13g2_nor2_1 _22135_ (.A(net4278),
    .B(net5143),
    .Y(_05121_));
 sg13g2_a21oi_1 _22136_ (.A1(net5701),
    .A2(net5143),
    .Y(_00731_),
    .B1(_05121_));
 sg13g2_nor2_1 _22137_ (.A(net3320),
    .B(net5144),
    .Y(_05122_));
 sg13g2_a21oi_1 _22138_ (.A1(net5682),
    .A2(net5144),
    .Y(_00732_),
    .B1(_05122_));
 sg13g2_nor2_1 _22139_ (.A(net3051),
    .B(net5144),
    .Y(_05123_));
 sg13g2_a21oi_1 _22140_ (.A1(net5604),
    .A2(net5144),
    .Y(_00733_),
    .B1(_05123_));
 sg13g2_nor2_1 _22141_ (.A(net3571),
    .B(net5144),
    .Y(_05124_));
 sg13g2_a21oi_1 _22142_ (.A1(net5658),
    .A2(net5144),
    .Y(_00734_),
    .B1(_05124_));
 sg13g2_nor2_1 _22143_ (.A(net3738),
    .B(net5144),
    .Y(_05125_));
 sg13g2_a21oi_1 _22144_ (.A1(net5635),
    .A2(net5144),
    .Y(_00735_),
    .B1(_05125_));
 sg13g2_nor2_1 _22145_ (.A(net6257),
    .B(_08771_),
    .Y(_05126_));
 sg13g2_a21oi_2 _22146_ (.B1(_09047_),
    .Y(_05127_),
    .A2(_05126_),
    .A1(\atari2600.cpu.load_reg ));
 sg13g2_or2_1 _22147_ (.X(_05128_),
    .B(_05127_),
    .A(net5858));
 sg13g2_inv_1 _22148_ (.Y(_05129_),
    .A(_05128_));
 sg13g2_and2_2 _22149_ (.A(_09058_),
    .B(_05129_),
    .X(_05130_));
 sg13g2_nor2_1 _22150_ (.A(net6253),
    .B(net6033),
    .Y(_05131_));
 sg13g2_a21oi_2 _22151_ (.B1(_05131_),
    .Y(_05132_),
    .A2(_08853_),
    .A1(_08731_));
 sg13g2_mux2_1 _22152_ (.A0(net4095),
    .A1(_05132_),
    .S(_05130_),
    .X(_00736_));
 sg13g2_nor2_1 _22153_ (.A(\atari2600.cpu.adc_bcd ),
    .B(_00163_),
    .Y(_05133_));
 sg13g2_nand2b_1 _22154_ (.Y(_05134_),
    .B(_05133_),
    .A_N(\atari2600.cpu.ALU.HC ));
 sg13g2_nand2_1 _22155_ (.Y(_05135_),
    .A(\atari2600.cpu.adc_bcd ),
    .B(\atari2600.cpu.ALU.HC ));
 sg13g2_o21ai_1 _22156_ (.B1(_05134_),
    .Y(_05136_),
    .A1(_00163_),
    .A2(_05135_));
 sg13g2_xnor2_1 _22157_ (.Y(_05137_),
    .A(_00074_),
    .B(_05136_));
 sg13g2_nor2_1 _22158_ (.A(net6032),
    .B(_05137_),
    .Y(_05138_));
 sg13g2_a21oi_2 _22159_ (.B1(_05138_),
    .Y(_05139_),
    .A2(net6032),
    .A1(_08735_));
 sg13g2_mux2_1 _22160_ (.A0(net4306),
    .A1(_05139_),
    .S(_05130_),
    .X(_00737_));
 sg13g2_nand2_1 _22161_ (.Y(_05140_),
    .A(net5827),
    .B(net6032));
 sg13g2_nand3_1 _22162_ (.B(\atari2600.cpu.adj_bcd ),
    .C(\atari2600.cpu.ALU.HC ),
    .A(\atari2600.cpu.adc_bcd ),
    .Y(_05141_));
 sg13g2_xnor2_1 _22163_ (.Y(_05142_),
    .A(net6251),
    .B(_05141_));
 sg13g2_a21oi_1 _22164_ (.A1(net6252),
    .A2(_05136_),
    .Y(_05143_),
    .B1(_05142_));
 sg13g2_nand3_1 _22165_ (.B(_05136_),
    .C(_05142_),
    .A(net6252),
    .Y(_05144_));
 sg13g2_nand2_1 _22166_ (.Y(_05145_),
    .A(net5997),
    .B(_05144_));
 sg13g2_o21ai_1 _22167_ (.B1(_05140_),
    .Y(_05146_),
    .A1(_05143_),
    .A2(_05145_));
 sg13g2_mux2_1 _22168_ (.A0(net3166),
    .A1(_05146_),
    .S(_05130_),
    .X(_00738_));
 sg13g2_nand2_1 _22169_ (.Y(_05147_),
    .A(net5826),
    .B(net6032));
 sg13g2_o21ai_1 _22170_ (.B1(_05144_),
    .Y(_05148_),
    .A1(_08580_),
    .A2(_05141_));
 sg13g2_xor2_1 _22171_ (.B(_05134_),
    .A(_00090_),
    .X(_05149_));
 sg13g2_xnor2_1 _22172_ (.Y(_05150_),
    .A(_05148_),
    .B(_05149_));
 sg13g2_o21ai_1 _22173_ (.B1(_05147_),
    .Y(_05151_),
    .A1(net6032),
    .A2(_05150_));
 sg13g2_mux2_1 _22174_ (.A0(net3871),
    .A1(_05151_),
    .S(_05130_),
    .X(_00739_));
 sg13g2_nor2_1 _22175_ (.A(\atari2600.cpu.ADD[4] ),
    .B(net6032),
    .Y(_05152_));
 sg13g2_a21oi_2 _22176_ (.B1(_05152_),
    .Y(_05153_),
    .A2(net6032),
    .A1(_08749_));
 sg13g2_mux2_1 _22177_ (.A0(net3334),
    .A1(_05153_),
    .S(_05130_),
    .X(_00740_));
 sg13g2_nand2_1 _22178_ (.Y(_05154_),
    .A(_08592_),
    .B(_05133_));
 sg13g2_nand2_1 _22179_ (.Y(_05155_),
    .A(net6247),
    .B(\atari2600.cpu.adc_bcd ));
 sg13g2_o21ai_1 _22180_ (.B1(_05154_),
    .Y(_05156_),
    .A1(_00163_),
    .A2(_05155_));
 sg13g2_xnor2_1 _22181_ (.Y(_05157_),
    .A(_00086_),
    .B(_05156_));
 sg13g2_nand2_1 _22182_ (.Y(_05158_),
    .A(net5997),
    .B(_05157_));
 sg13g2_o21ai_1 _22183_ (.B1(_05158_),
    .Y(_05159_),
    .A1(_08759_),
    .A2(net5997));
 sg13g2_mux2_1 _22184_ (.A0(net3480),
    .A1(_05159_),
    .S(_05130_),
    .X(_00741_));
 sg13g2_nand2_1 _22185_ (.Y(_05160_),
    .A(net5825),
    .B(net6033));
 sg13g2_nand3_1 _22186_ (.B(\atari2600.cpu.adc_bcd ),
    .C(\atari2600.cpu.adj_bcd ),
    .A(net6247),
    .Y(_05161_));
 sg13g2_xnor2_1 _22187_ (.Y(_05162_),
    .A(net6248),
    .B(_05161_));
 sg13g2_a21oi_1 _22188_ (.A1(net6249),
    .A2(_05156_),
    .Y(_05163_),
    .B1(_05162_));
 sg13g2_nand3_1 _22189_ (.B(_05156_),
    .C(_05162_),
    .A(net6249),
    .Y(_05164_));
 sg13g2_nand2_1 _22190_ (.Y(_05165_),
    .A(net5997),
    .B(_05164_));
 sg13g2_o21ai_1 _22191_ (.B1(_05160_),
    .Y(_05166_),
    .A1(_05163_),
    .A2(_05165_));
 sg13g2_mux2_1 _22192_ (.A0(net3705),
    .A1(_05166_),
    .S(_05130_),
    .X(_00742_));
 sg13g2_nand2_1 _22193_ (.Y(_05167_),
    .A(\atari2600.cpu.DIMUX[7] ),
    .B(net6033));
 sg13g2_o21ai_1 _22194_ (.B1(_05164_),
    .Y(_05168_),
    .A1(_08594_),
    .A2(_05161_));
 sg13g2_xnor2_1 _22195_ (.Y(_05169_),
    .A(_08599_),
    .B(_05154_));
 sg13g2_xnor2_1 _22196_ (.Y(_05170_),
    .A(_05168_),
    .B(_05169_));
 sg13g2_o21ai_1 _22197_ (.B1(_05167_),
    .Y(_05171_),
    .A1(net6032),
    .A2(_05170_));
 sg13g2_mux2_1 _22198_ (.A0(net3338),
    .A1(_05171_),
    .S(_05130_),
    .X(_00743_));
 sg13g2_nand3_1 _22199_ (.B(_09321_),
    .C(net5250),
    .A(net5550),
    .Y(_05172_));
 sg13g2_mux2_1 _22200_ (.A0(net5739),
    .A1(net4750),
    .S(_05172_),
    .X(_00744_));
 sg13g2_mux2_1 _22201_ (.A0(net5749),
    .A1(net6821),
    .S(_05172_),
    .X(_00745_));
 sg13g2_mux2_1 _22202_ (.A0(net5618),
    .A1(net4716),
    .S(_05172_),
    .X(_00746_));
 sg13g2_mux2_1 _22203_ (.A0(net5612),
    .A1(net4600),
    .S(_05172_),
    .X(_00747_));
 sg13g2_mux2_1 _22204_ (.A0(_03045_),
    .A1(net4830),
    .S(_05172_),
    .X(_00748_));
 sg13g2_mux2_1 _22205_ (.A0(net5582),
    .A1(net4697),
    .S(_05172_),
    .X(_00749_));
 sg13g2_mux2_1 _22206_ (.A0(net5576),
    .A1(net4929),
    .S(_05172_),
    .X(_00750_));
 sg13g2_mux2_1 _22207_ (.A0(net5644),
    .A1(net6774),
    .S(_05172_),
    .X(_00751_));
 sg13g2_nor2_1 _22208_ (.A(_09441_),
    .B(net5254),
    .Y(_05173_));
 sg13g2_nor2_1 _22209_ (.A(net3094),
    .B(net5060),
    .Y(_05174_));
 sg13g2_a21oi_1 _22210_ (.A1(net5768),
    .A2(net5061),
    .Y(_00752_),
    .B1(_05174_));
 sg13g2_nor2_1 _22211_ (.A(net3294),
    .B(net5061),
    .Y(_05175_));
 sg13g2_a21oi_1 _22212_ (.A1(net5789),
    .A2(net5061),
    .Y(_00753_),
    .B1(_05175_));
 sg13g2_nor2_1 _22213_ (.A(net3096),
    .B(net5060),
    .Y(_05176_));
 sg13g2_a21oi_1 _22214_ (.A1(net5718),
    .A2(net5060),
    .Y(_00754_),
    .B1(_05176_));
 sg13g2_nor2_1 _22215_ (.A(net3810),
    .B(net5060),
    .Y(_05177_));
 sg13g2_a21oi_1 _22216_ (.A1(net5696),
    .A2(net5060),
    .Y(_00755_),
    .B1(_05177_));
 sg13g2_nor2_1 _22217_ (.A(net3127),
    .B(net5060),
    .Y(_05178_));
 sg13g2_a21oi_1 _22218_ (.A1(net5675),
    .A2(net5061),
    .Y(_00756_),
    .B1(_05178_));
 sg13g2_nor2_1 _22219_ (.A(net3227),
    .B(net5060),
    .Y(_05179_));
 sg13g2_a21oi_1 _22220_ (.A1(net5594),
    .A2(net5060),
    .Y(_00757_),
    .B1(_05179_));
 sg13g2_nor2_1 _22221_ (.A(net3293),
    .B(net5062),
    .Y(_05180_));
 sg13g2_a21oi_1 _22222_ (.A1(net5655),
    .A2(net5062),
    .Y(_00758_),
    .B1(_05180_));
 sg13g2_nor2_1 _22223_ (.A(net3004),
    .B(net5062),
    .Y(_05181_));
 sg13g2_a21oi_1 _22224_ (.A1(net5630),
    .A2(net5062),
    .Y(_00759_),
    .B1(_05181_));
 sg13g2_nand3_1 _22225_ (.B(_09421_),
    .C(net5252),
    .A(net5548),
    .Y(_05182_));
 sg13g2_mux2_1 _22226_ (.A0(net5740),
    .A1(net7073),
    .S(_05182_),
    .X(_00760_));
 sg13g2_mux2_1 _22227_ (.A0(net5745),
    .A1(net6641),
    .S(_05182_),
    .X(_00761_));
 sg13g2_mux2_1 _22228_ (.A0(net5616),
    .A1(net4838),
    .S(_05182_),
    .X(_00762_));
 sg13g2_mux2_1 _22229_ (.A0(net5611),
    .A1(net4545),
    .S(_05182_),
    .X(_00763_));
 sg13g2_mux2_1 _22230_ (.A0(net5607),
    .A1(net4506),
    .S(_05182_),
    .X(_00764_));
 sg13g2_mux2_1 _22231_ (.A0(net5580),
    .A1(net4590),
    .S(_05182_),
    .X(_00765_));
 sg13g2_mux2_1 _22232_ (.A0(net5575),
    .A1(net4595),
    .S(_05182_),
    .X(_00766_));
 sg13g2_mux2_1 _22233_ (.A0(net5641),
    .A1(net4478),
    .S(_05182_),
    .X(_00767_));
 sg13g2_nor2_1 _22234_ (.A(net5263),
    .B(net5237),
    .Y(_05183_));
 sg13g2_nor2_1 _22235_ (.A(net3112),
    .B(net5142),
    .Y(_05184_));
 sg13g2_a21oi_1 _22236_ (.A1(net5761),
    .A2(net5142),
    .Y(_00768_),
    .B1(_05184_));
 sg13g2_nor2_1 _22237_ (.A(net3644),
    .B(net5142),
    .Y(_05185_));
 sg13g2_a21oi_1 _22238_ (.A1(net5784),
    .A2(net5142),
    .Y(_00769_),
    .B1(_05185_));
 sg13g2_nor2_1 _22239_ (.A(net4198),
    .B(net5142),
    .Y(_05186_));
 sg13g2_a21oi_1 _22240_ (.A1(net5710),
    .A2(net5142),
    .Y(_00770_),
    .B1(_05186_));
 sg13g2_nor2_1 _22241_ (.A(net3015),
    .B(net5141),
    .Y(_05187_));
 sg13g2_a21oi_1 _22242_ (.A1(net5687),
    .A2(net5141),
    .Y(_00771_),
    .B1(_05187_));
 sg13g2_nor2_1 _22243_ (.A(net4290),
    .B(net5142),
    .Y(_05188_));
 sg13g2_a21oi_1 _22244_ (.A1(net5671),
    .A2(net5142),
    .Y(_00772_),
    .B1(_05188_));
 sg13g2_nor2_1 _22245_ (.A(net4438),
    .B(net5141),
    .Y(_05189_));
 sg13g2_a21oi_1 _22246_ (.A1(net5588),
    .A2(net5141),
    .Y(_00773_),
    .B1(_05189_));
 sg13g2_nor2_1 _22247_ (.A(net3048),
    .B(net5141),
    .Y(_05190_));
 sg13g2_a21oi_1 _22248_ (.A1(net5648),
    .A2(net5141),
    .Y(_00774_),
    .B1(_05190_));
 sg13g2_nor2_1 _22249_ (.A(net3491),
    .B(net5141),
    .Y(_05191_));
 sg13g2_a21oi_1 _22250_ (.A1(net5624),
    .A2(net5141),
    .Y(_00775_),
    .B1(_05191_));
 sg13g2_nand3_1 _22251_ (.B(_09318_),
    .C(net5250),
    .A(_09262_),
    .Y(_05192_));
 sg13g2_mux2_1 _22252_ (.A0(net5739),
    .A1(net4873),
    .S(_05192_),
    .X(_00776_));
 sg13g2_mux2_1 _22253_ (.A0(net5744),
    .A1(net4696),
    .S(_05192_),
    .X(_00777_));
 sg13g2_mux2_1 _22254_ (.A0(net5616),
    .A1(net4908),
    .S(_05192_),
    .X(_00778_));
 sg13g2_mux2_1 _22255_ (.A0(net5611),
    .A1(net4819),
    .S(_05192_),
    .X(_00779_));
 sg13g2_mux2_1 _22256_ (.A0(net5606),
    .A1(net4519),
    .S(_05192_),
    .X(_00780_));
 sg13g2_mux2_1 _22257_ (.A0(net5580),
    .A1(net6646),
    .S(_05192_),
    .X(_00781_));
 sg13g2_mux2_1 _22258_ (.A0(net5576),
    .A1(net4660),
    .S(_05192_),
    .X(_00782_));
 sg13g2_mux2_1 _22259_ (.A0(net5641),
    .A1(net4513),
    .S(_05192_),
    .X(_00783_));
 sg13g2_nor2_1 _22260_ (.A(net5254),
    .B(_03124_),
    .Y(_05193_));
 sg13g2_nor2_1 _22261_ (.A(net3045),
    .B(net5139),
    .Y(_05194_));
 sg13g2_a21oi_1 _22262_ (.A1(net5775),
    .A2(net5139),
    .Y(_00784_),
    .B1(_05194_));
 sg13g2_nor2_1 _22263_ (.A(net3160),
    .B(net5140),
    .Y(_05195_));
 sg13g2_a21oi_1 _22264_ (.A1(net5795),
    .A2(net5140),
    .Y(_00785_),
    .B1(_05195_));
 sg13g2_nor2_1 _22265_ (.A(net3241),
    .B(net5140),
    .Y(_05196_));
 sg13g2_a21oi_1 _22266_ (.A1(net5724),
    .A2(net5140),
    .Y(_00786_),
    .B1(_05196_));
 sg13g2_nor2_1 _22267_ (.A(net3172),
    .B(net5140),
    .Y(_05197_));
 sg13g2_a21oi_1 _22268_ (.A1(net5701),
    .A2(net5140),
    .Y(_00787_),
    .B1(_05197_));
 sg13g2_nor2_1 _22269_ (.A(net3453),
    .B(net5139),
    .Y(_05198_));
 sg13g2_a21oi_1 _22270_ (.A1(net5680),
    .A2(net5140),
    .Y(_00788_),
    .B1(_05198_));
 sg13g2_nor2_1 _22271_ (.A(net3505),
    .B(net5139),
    .Y(_05199_));
 sg13g2_a21oi_1 _22272_ (.A1(net5602),
    .A2(net5139),
    .Y(_00789_),
    .B1(_05199_));
 sg13g2_nor2_1 _22273_ (.A(net3495),
    .B(net5139),
    .Y(_05200_));
 sg13g2_a21oi_1 _22274_ (.A1(net5663),
    .A2(net5139),
    .Y(_00790_),
    .B1(_05200_));
 sg13g2_nor2_1 _22275_ (.A(net3630),
    .B(net5139),
    .Y(_05201_));
 sg13g2_a21oi_1 _22276_ (.A1(net5638),
    .A2(_05193_),
    .Y(_00791_),
    .B1(_05201_));
 sg13g2_nand2b_2 _22277_ (.Y(_05202_),
    .B(net5253),
    .A_N(_03091_));
 sg13g2_mux2_1 _22278_ (.A0(net5741),
    .A1(net4804),
    .S(_05202_),
    .X(_00792_));
 sg13g2_mux2_1 _22279_ (.A0(net5746),
    .A1(net6911),
    .S(_05202_),
    .X(_00793_));
 sg13g2_mux2_1 _22280_ (.A0(net5617),
    .A1(net4859),
    .S(_05202_),
    .X(_00794_));
 sg13g2_mux2_1 _22281_ (.A0(net5614),
    .A1(net4530),
    .S(_05202_),
    .X(_00795_));
 sg13g2_mux2_1 _22282_ (.A0(net5609),
    .A1(net6838),
    .S(_05202_),
    .X(_00796_));
 sg13g2_mux2_1 _22283_ (.A0(net5583),
    .A1(net4568),
    .S(_05202_),
    .X(_00797_));
 sg13g2_mux2_1 _22284_ (.A0(net5577),
    .A1(net4837),
    .S(_05202_),
    .X(_00798_));
 sg13g2_mux2_1 _22285_ (.A0(net5643),
    .A1(net6691),
    .S(_05202_),
    .X(_00799_));
 sg13g2_nor2_1 _22286_ (.A(_03021_),
    .B(net5236),
    .Y(_05203_));
 sg13g2_nor2_1 _22287_ (.A(net4329),
    .B(net5138),
    .Y(_05204_));
 sg13g2_a21oi_1 _22288_ (.A1(net5774),
    .A2(net5138),
    .Y(_00800_),
    .B1(_05204_));
 sg13g2_nor2_1 _22289_ (.A(net3210),
    .B(net5138),
    .Y(_05205_));
 sg13g2_a21oi_1 _22290_ (.A1(net5794),
    .A2(net5138),
    .Y(_00801_),
    .B1(_05205_));
 sg13g2_nor2_1 _22291_ (.A(net3224),
    .B(net5138),
    .Y(_05206_));
 sg13g2_a21oi_1 _22292_ (.A1(net5724),
    .A2(net5138),
    .Y(_00802_),
    .B1(_05206_));
 sg13g2_nor2_1 _22293_ (.A(net3466),
    .B(net5138),
    .Y(_05207_));
 sg13g2_a21oi_1 _22294_ (.A1(net5700),
    .A2(_05203_),
    .Y(_00803_),
    .B1(_05207_));
 sg13g2_nor2_1 _22295_ (.A(net4415),
    .B(net5137),
    .Y(_05208_));
 sg13g2_a21oi_1 _22296_ (.A1(net5681),
    .A2(net5137),
    .Y(_00804_),
    .B1(_05208_));
 sg13g2_nor2_1 _22297_ (.A(net3268),
    .B(net5137),
    .Y(_05209_));
 sg13g2_a21oi_1 _22298_ (.A1(net5601),
    .A2(net5137),
    .Y(_00805_),
    .B1(_05209_));
 sg13g2_nor2_1 _22299_ (.A(net3168),
    .B(net5137),
    .Y(_05210_));
 sg13g2_a21oi_1 _22300_ (.A1(net5658),
    .A2(net5137),
    .Y(_00806_),
    .B1(_05210_));
 sg13g2_nor2_1 _22301_ (.A(net3305),
    .B(net5137),
    .Y(_05211_));
 sg13g2_a21oi_1 _22302_ (.A1(net5636),
    .A2(net5137),
    .Y(_00807_),
    .B1(_05211_));
 sg13g2_nand2_2 _22303_ (.Y(_05212_),
    .A(net5251),
    .B(_04880_));
 sg13g2_mux2_1 _22304_ (.A0(net5741),
    .A1(net6794),
    .S(_05212_),
    .X(_00808_));
 sg13g2_mux2_1 _22305_ (.A0(net5746),
    .A1(net4596),
    .S(_05212_),
    .X(_00809_));
 sg13g2_mux2_1 _22306_ (.A0(net5619),
    .A1(net6915),
    .S(_05212_),
    .X(_00810_));
 sg13g2_mux2_1 _22307_ (.A0(net5612),
    .A1(net4628),
    .S(_05212_),
    .X(_00811_));
 sg13g2_mux2_1 _22308_ (.A0(net5608),
    .A1(net6725),
    .S(_05212_),
    .X(_00812_));
 sg13g2_mux2_1 _22309_ (.A0(net5583),
    .A1(net6919),
    .S(_05212_),
    .X(_00813_));
 sg13g2_mux2_1 _22310_ (.A0(net5577),
    .A1(net6762),
    .S(_05212_),
    .X(_00814_));
 sg13g2_mux2_1 _22311_ (.A0(net5645),
    .A1(net6947),
    .S(_05212_),
    .X(_00815_));
 sg13g2_nor2_1 _22312_ (.A(net5254),
    .B(_04947_),
    .Y(_05213_));
 sg13g2_nor2_1 _22313_ (.A(net3903),
    .B(net5220),
    .Y(_05214_));
 sg13g2_a21oi_1 _22314_ (.A1(net5770),
    .A2(net5220),
    .Y(_00816_),
    .B1(_05214_));
 sg13g2_nor2_1 _22315_ (.A(net3757),
    .B(_05213_),
    .Y(_05215_));
 sg13g2_a21oi_1 _22316_ (.A1(net5791),
    .A2(net5219),
    .Y(_00817_),
    .B1(_05215_));
 sg13g2_nor2_1 _22317_ (.A(net3135),
    .B(net5219),
    .Y(_05216_));
 sg13g2_a21oi_1 _22318_ (.A1(net5721),
    .A2(net5219),
    .Y(_00818_),
    .B1(_05216_));
 sg13g2_nor2_1 _22319_ (.A(net3275),
    .B(net5219),
    .Y(_05217_));
 sg13g2_a21oi_1 _22320_ (.A1(net5698),
    .A2(net5220),
    .Y(_00819_),
    .B1(_05217_));
 sg13g2_nor2_1 _22321_ (.A(net3147),
    .B(net5220),
    .Y(_05218_));
 sg13g2_a21oi_1 _22322_ (.A1(net5676),
    .A2(net5220),
    .Y(_00820_),
    .B1(_05218_));
 sg13g2_nor2_1 _22323_ (.A(net3319),
    .B(net5220),
    .Y(_05219_));
 sg13g2_a21oi_1 _22324_ (.A1(net5596),
    .A2(net5220),
    .Y(_00821_),
    .B1(_05219_));
 sg13g2_nor2_1 _22325_ (.A(net3773),
    .B(net5219),
    .Y(_05220_));
 sg13g2_a21oi_1 _22326_ (.A1(net5660),
    .A2(net5219),
    .Y(_00822_),
    .B1(_05220_));
 sg13g2_nor2_1 _22327_ (.A(net4015),
    .B(net5219),
    .Y(_05221_));
 sg13g2_a21oi_1 _22328_ (.A1(net5634),
    .A2(net5219),
    .Y(_00823_),
    .B1(_05221_));
 sg13g2_nand2_2 _22329_ (.Y(_05222_),
    .A(net5253),
    .B(_05004_));
 sg13g2_mux2_1 _22330_ (.A0(net5741),
    .A1(net4875),
    .S(_05222_),
    .X(_00824_));
 sg13g2_mux2_1 _22331_ (.A0(net5746),
    .A1(net6950),
    .S(_05222_),
    .X(_00825_));
 sg13g2_mux2_1 _22332_ (.A0(net5617),
    .A1(net4917),
    .S(_05222_),
    .X(_00826_));
 sg13g2_mux2_1 _22333_ (.A0(net5614),
    .A1(net6896),
    .S(_05222_),
    .X(_00827_));
 sg13g2_mux2_1 _22334_ (.A0(net5608),
    .A1(net4850),
    .S(_05222_),
    .X(_00828_));
 sg13g2_mux2_1 _22335_ (.A0(net5581),
    .A1(net4955),
    .S(_05222_),
    .X(_00829_));
 sg13g2_mux2_1 _22336_ (.A0(net5578),
    .A1(net6610),
    .S(_05222_),
    .X(_00830_));
 sg13g2_mux2_1 _22337_ (.A0(net5644),
    .A1(net4900),
    .S(_05222_),
    .X(_00831_));
 sg13g2_nor2_1 _22338_ (.A(net5258),
    .B(_03091_),
    .Y(_05223_));
 sg13g2_nor2_1 _22339_ (.A(net4214),
    .B(net5135),
    .Y(_05224_));
 sg13g2_a21oi_1 _22340_ (.A1(net5772),
    .A2(net5135),
    .Y(_00832_),
    .B1(_05224_));
 sg13g2_nor2_1 _22341_ (.A(net4184),
    .B(net5136),
    .Y(_05225_));
 sg13g2_a21oi_1 _22342_ (.A1(net5793),
    .A2(net5136),
    .Y(_00833_),
    .B1(_05225_));
 sg13g2_nor2_1 _22343_ (.A(net4273),
    .B(net5136),
    .Y(_05226_));
 sg13g2_a21oi_1 _22344_ (.A1(net5723),
    .A2(net5136),
    .Y(_00834_),
    .B1(_05226_));
 sg13g2_nor2_1 _22345_ (.A(net4287),
    .B(net5136),
    .Y(_05227_));
 sg13g2_a21oi_1 _22346_ (.A1(net5699),
    .A2(net5136),
    .Y(_00835_),
    .B1(_05227_));
 sg13g2_nor2_1 _22347_ (.A(net4296),
    .B(net5136),
    .Y(_05228_));
 sg13g2_a21oi_1 _22348_ (.A1(net5679),
    .A2(_05223_),
    .Y(_00836_),
    .B1(_05228_));
 sg13g2_nor2_1 _22349_ (.A(net3349),
    .B(net5135),
    .Y(_05229_));
 sg13g2_a21oi_1 _22350_ (.A1(net5599),
    .A2(net5135),
    .Y(_00837_),
    .B1(_05229_));
 sg13g2_nor2_1 _22351_ (.A(net3391),
    .B(net5135),
    .Y(_05230_));
 sg13g2_a21oi_1 _22352_ (.A1(net5661),
    .A2(net5135),
    .Y(_00838_),
    .B1(_05230_));
 sg13g2_nor2_1 _22353_ (.A(net3873),
    .B(net5135),
    .Y(_05231_));
 sg13g2_a21oi_1 _22354_ (.A1(net5633),
    .A2(net5135),
    .Y(_00839_),
    .B1(_05231_));
 sg13g2_nand2b_2 _22355_ (.Y(_05232_),
    .B(net5251),
    .A_N(_03091_));
 sg13g2_mux2_1 _22356_ (.A0(net5741),
    .A1(net4629),
    .S(_05232_),
    .X(_00840_));
 sg13g2_mux2_1 _22357_ (.A0(net5746),
    .A1(net6593),
    .S(_05232_),
    .X(_00841_));
 sg13g2_mux2_1 _22358_ (.A0(net5617),
    .A1(net7012),
    .S(_05232_),
    .X(_00842_));
 sg13g2_mux2_1 _22359_ (.A0(net5614),
    .A1(net4515),
    .S(_05232_),
    .X(_00843_));
 sg13g2_mux2_1 _22360_ (.A0(net5608),
    .A1(net6958),
    .S(_05232_),
    .X(_00844_));
 sg13g2_mux2_1 _22361_ (.A0(net5584),
    .A1(net4576),
    .S(_05232_),
    .X(_00845_));
 sg13g2_mux2_1 _22362_ (.A0(net5577),
    .A1(net4748),
    .S(_05232_),
    .X(_00846_));
 sg13g2_mux2_1 _22363_ (.A0(net5643),
    .A1(net4911),
    .S(_05232_),
    .X(_00847_));
 sg13g2_nand3_1 _22364_ (.B(_09421_),
    .C(net5250),
    .A(net5548),
    .Y(_05233_));
 sg13g2_mux2_1 _22365_ (.A0(net5740),
    .A1(net4825),
    .S(_05233_),
    .X(_00848_));
 sg13g2_mux2_1 _22366_ (.A0(net5745),
    .A1(net4580),
    .S(_05233_),
    .X(_00849_));
 sg13g2_mux2_1 _22367_ (.A0(net5616),
    .A1(net6628),
    .S(_05233_),
    .X(_00850_));
 sg13g2_mux2_1 _22368_ (.A0(net5611),
    .A1(net4632),
    .S(_05233_),
    .X(_00851_));
 sg13g2_mux2_1 _22369_ (.A0(net5607),
    .A1(net4676),
    .S(_05233_),
    .X(_00852_));
 sg13g2_mux2_1 _22370_ (.A0(net5580),
    .A1(net7064),
    .S(_05233_),
    .X(_00853_));
 sg13g2_mux2_1 _22371_ (.A0(net5575),
    .A1(net4566),
    .S(_05233_),
    .X(_00854_));
 sg13g2_mux2_1 _22372_ (.A0(net5641),
    .A1(net4738),
    .S(_05233_),
    .X(_00855_));
 sg13g2_nand2_1 _22373_ (.Y(_05234_),
    .A(net3203),
    .B(net5858));
 sg13g2_nand2_2 _22374_ (.Y(_05235_),
    .A(_08796_),
    .B(_09066_));
 sg13g2_nand2_2 _22375_ (.Y(_05236_),
    .A(\atari2600.cpu.op[3] ),
    .B(_05235_));
 sg13g2_nand2_2 _22376_ (.Y(_05237_),
    .A(_08891_),
    .B(_08920_));
 sg13g2_inv_1 _22377_ (.Y(_05238_),
    .A(_05237_));
 sg13g2_and3_1 _22378_ (.X(_05239_),
    .A(_08939_),
    .B(_09068_),
    .C(_05238_));
 sg13g2_nand3_1 _22379_ (.B(_08995_),
    .C(_09042_),
    .A(_08792_),
    .Y(_05240_));
 sg13g2_nand3_1 _22380_ (.B(_08914_),
    .C(_09069_),
    .A(_08879_),
    .Y(_05241_));
 sg13g2_nor2_1 _22381_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sg13g2_and3_2 _22382_ (.X(_05243_),
    .A(_04856_),
    .B(_05239_),
    .C(_05242_));
 sg13g2_nand3_1 _22383_ (.B(_05239_),
    .C(_05242_),
    .A(_04856_),
    .Y(_05244_));
 sg13g2_nand2_1 _22384_ (.Y(_05245_),
    .A(\atari2600.cpu.PC[7] ),
    .B(net5991));
 sg13g2_o21ai_1 _22385_ (.B1(_05245_),
    .Y(_05246_),
    .A1(_08744_),
    .A2(_05244_));
 sg13g2_a221oi_1 _22386_ (.B2(\atari2600.cpu.op[2] ),
    .C1(_09108_),
    .B1(_05235_),
    .A1(\atari2600.cpu.backwards ),
    .Y(_05247_),
    .A2(net5995));
 sg13g2_xnor2_1 _22387_ (.Y(_05248_),
    .A(_05246_),
    .B(net5915));
 sg13g2_and2_1 _22388_ (.A(net5917),
    .B(_05248_),
    .X(_05249_));
 sg13g2_a21oi_2 _22389_ (.B1(_08587_),
    .Y(_05250_),
    .A2(_09066_),
    .A1(_08796_));
 sg13g2_o21ai_1 _22390_ (.B1(net6247),
    .Y(_05251_),
    .A1(net5995),
    .A2(_09075_));
 sg13g2_a21oi_2 _22391_ (.B1(\atari2600.cpu.rotate ),
    .Y(_05252_),
    .A2(\atari2600.cpu.inc ),
    .A1(_08590_));
 sg13g2_nor2_1 _22392_ (.A(\atari2600.cpu.C ),
    .B(_08591_),
    .Y(_05253_));
 sg13g2_or3_1 _22393_ (.A(_09066_),
    .B(_05252_),
    .C(_05253_),
    .X(_05254_));
 sg13g2_o21ai_1 _22394_ (.B1(_08591_),
    .Y(_05255_),
    .A1(\atari2600.cpu.load_only ),
    .A2(\atari2600.cpu.shift ));
 sg13g2_a22oi_1 _22395_ (.Y(_05256_),
    .B1(_05255_),
    .B2(_08583_),
    .A2(_08591_),
    .A1(\atari2600.cpu.compare ));
 sg13g2_nor2_1 _22396_ (.A(_08796_),
    .B(_05256_),
    .Y(_05257_));
 sg13g2_nand4_1 _22397_ (.B(_09043_),
    .C(_05251_),
    .A(_08937_),
    .Y(_05258_),
    .D(_05254_));
 sg13g2_nor4_2 _22398_ (.A(_08859_),
    .B(_05241_),
    .C(_05257_),
    .Y(_05259_),
    .D(_05258_));
 sg13g2_nor2b_1 _22399_ (.A(_05259_),
    .B_N(net5934),
    .Y(_05260_));
 sg13g2_nor3_2 _22400_ (.A(net6034),
    .B(_08806_),
    .C(_05235_),
    .Y(_05261_));
 sg13g2_a21oi_2 _22401_ (.B1(_08586_),
    .Y(_05262_),
    .A2(_09066_),
    .A1(_08796_));
 sg13g2_nor2_2 _22402_ (.A(_05261_),
    .B(_05262_),
    .Y(_05263_));
 sg13g2_or2_1 _22403_ (.X(_05264_),
    .B(_05262_),
    .A(_05261_));
 sg13g2_a21oi_2 _22404_ (.B1(_05261_),
    .Y(_05265_),
    .A2(_05235_),
    .A1(\atari2600.cpu.op[0] ));
 sg13g2_nand3_1 _22405_ (.B(_08586_),
    .C(_05235_),
    .A(\atari2600.cpu.op[0] ),
    .Y(_05266_));
 sg13g2_o21ai_1 _22406_ (.B1(_04868_),
    .Y(_05267_),
    .A1(\atari2600.cpu.load_only ),
    .A2(_08796_));
 sg13g2_or4_2 _22407_ (.A(_09044_),
    .B(_09051_),
    .C(_05240_),
    .D(_05267_),
    .X(_05268_));
 sg13g2_a22oi_1 _22408_ (.Y(_05269_),
    .B1(net5928),
    .B2(\atari2600.cpu.ADD[7] ),
    .A2(net5993),
    .A1(\atari2600.cpu.ABH[7] ));
 sg13g2_a22oi_1 _22409_ (.Y(_05270_),
    .B1(_05268_),
    .B2(_09116_),
    .A2(_05237_),
    .A1(\atari2600.cpu.DIMUX[7] ));
 sg13g2_nand2_2 _22410_ (.Y(_05271_),
    .A(_05269_),
    .B(_05270_));
 sg13g2_nand3_1 _22411_ (.B(net5875),
    .C(_05271_),
    .A(_05246_),
    .Y(_05272_));
 sg13g2_a22oi_1 _22412_ (.Y(_05273_),
    .B1(_05266_),
    .B2(_05272_),
    .A2(_05263_),
    .A1(_05246_));
 sg13g2_a21oi_1 _22413_ (.A1(_05246_),
    .A2(net5875),
    .Y(_05274_),
    .B1(_05271_));
 sg13g2_nor3_2 _22414_ (.A(net5934),
    .B(_05273_),
    .C(_05274_),
    .Y(_05275_));
 sg13g2_nor3_2 _22415_ (.A(_05249_),
    .B(_05260_),
    .C(_05275_),
    .Y(_05276_));
 sg13g2_nor2b_1 _22416_ (.A(net5917),
    .B_N(net5916),
    .Y(_05277_));
 sg13g2_nand2b_2 _22417_ (.Y(_05278_),
    .B(net5915),
    .A_N(_05236_));
 sg13g2_nand2b_1 _22418_ (.Y(_05279_),
    .B(_05278_),
    .A_N(_05249_));
 sg13g2_nand2_1 _22419_ (.Y(_05280_),
    .A(net5828),
    .B(_05279_));
 sg13g2_o21ai_1 _22420_ (.B1(_05234_),
    .Y(_00856_),
    .A1(_05276_),
    .A2(_05280_));
 sg13g2_nor3_2 _22421_ (.A(net7447),
    .B(_08679_),
    .C(net5929),
    .Y(_05281_));
 sg13g2_and2_1 _22422_ (.A(net6246),
    .B(_05281_),
    .X(_05282_));
 sg13g2_nand2_2 _22423_ (.Y(_05283_),
    .A(net6246),
    .B(_05281_));
 sg13g2_nor4_1 _22424_ (.A(\atari2600.pia.reset_timer[4] ),
    .B(\atari2600.pia.reset_timer[3] ),
    .C(\atari2600.pia.reset_timer[2] ),
    .D(\atari2600.pia.reset_timer[1] ),
    .Y(_05284_));
 sg13g2_nor4_1 _22425_ (.A(\atari2600.pia.reset_timer[0] ),
    .B(\atari2600.pia.reset_timer[7] ),
    .C(\atari2600.pia.reset_timer[6] ),
    .D(\atari2600.pia.reset_timer[5] ),
    .Y(_05285_));
 sg13g2_and2_2 _22426_ (.A(_05284_),
    .B(_05285_),
    .X(_05286_));
 sg13g2_nand2_1 _22427_ (.Y(_05287_),
    .A(_05284_),
    .B(_05285_));
 sg13g2_nor2_1 _22428_ (.A(\atari2600.pia.underflow ),
    .B(\atari2600.pia.interval[0] ),
    .Y(_05288_));
 sg13g2_nor3_2 _22429_ (.A(\atari2600.pia.interval[3] ),
    .B(\atari2600.pia.underflow ),
    .C(\atari2600.pia.interval[0] ),
    .Y(_05289_));
 sg13g2_nand2b_1 _22430_ (.Y(_05290_),
    .B(_05288_),
    .A_N(\atari2600.pia.interval[3] ));
 sg13g2_nor2_1 _22431_ (.A(\atari2600.pia.interval[6] ),
    .B(_05290_),
    .Y(_05291_));
 sg13g2_nor2b_1 _22432_ (.A(\atari2600.pia.underflow ),
    .B_N(\atari2600.pia.interval[6] ),
    .Y(_05292_));
 sg13g2_a21oi_1 _22433_ (.A1(_05290_),
    .A2(_05292_),
    .Y(_05293_),
    .B1(_05291_));
 sg13g2_nor2_1 _22434_ (.A(net7203),
    .B(net7018),
    .Y(_05294_));
 sg13g2_and2_1 _22435_ (.A(\atari2600.pia.time_counter[9] ),
    .B(\atari2600.pia.time_counter[8] ),
    .X(_05295_));
 sg13g2_mux2_1 _22436_ (.A0(_05294_),
    .A1(_05295_),
    .S(_05291_),
    .X(_05296_));
 sg13g2_nor2b_1 _22437_ (.A(\atari2600.pia.underflow ),
    .B_N(\atari2600.pia.interval[10] ),
    .Y(_05297_));
 sg13g2_nand3b_1 _22438_ (.B(_05289_),
    .C(\atari2600.pia.time_counter[7] ),
    .Y(_05298_),
    .A_N(_05292_));
 sg13g2_and3_1 _22439_ (.X(_05299_),
    .A(_00084_),
    .B(_05297_),
    .C(_05298_));
 sg13g2_and2_1 _22440_ (.A(\atari2600.pia.time_counter[5] ),
    .B(\atari2600.pia.time_counter[4] ),
    .X(_05300_));
 sg13g2_nor3_1 _22441_ (.A(\atari2600.pia.time_counter[5] ),
    .B(\atari2600.pia.time_counter[4] ),
    .C(_05289_),
    .Y(_05301_));
 sg13g2_a21oi_1 _22442_ (.A1(_05289_),
    .A2(_05300_),
    .Y(_05302_),
    .B1(_05301_));
 sg13g2_nand3b_1 _22443_ (.B(\atari2600.pia.interval[0] ),
    .C(\atari2600.pia.interval[3] ),
    .Y(_05303_),
    .A_N(\atari2600.pia.underflow ));
 sg13g2_a21oi_1 _22444_ (.A1(_05290_),
    .A2(_05303_),
    .Y(_05304_),
    .B1(\atari2600.pia.time_counter[3] ));
 sg13g2_nor2_1 _22445_ (.A(\atari2600.pia.time_counter[8] ),
    .B(\atari2600.pia.time_counter[7] ),
    .Y(_05305_));
 sg13g2_a21oi_1 _22446_ (.A1(_00084_),
    .A2(_05297_),
    .Y(_05306_),
    .B1(_05305_));
 sg13g2_nor3_1 _22447_ (.A(\atari2600.pia.time_counter[2] ),
    .B(\atari2600.pia.time_counter[1] ),
    .C(_05288_),
    .Y(_05307_));
 sg13g2_nand3_1 _22448_ (.B(\atari2600.pia.time_counter[1] ),
    .C(_05288_),
    .A(\atari2600.pia.time_counter[2] ),
    .Y(_05308_));
 sg13g2_nand2b_1 _22449_ (.Y(_05309_),
    .B(_05308_),
    .A_N(_05307_));
 sg13g2_nor2_1 _22450_ (.A(\atari2600.pia.time_counter[23] ),
    .B(\atari2600.pia.time_counter[22] ),
    .Y(_05310_));
 sg13g2_nor4_1 _22451_ (.A(\atari2600.pia.time_counter[21] ),
    .B(\atari2600.pia.time_counter[20] ),
    .C(\atari2600.pia.time_counter[19] ),
    .D(\atari2600.pia.time_counter[18] ),
    .Y(_05311_));
 sg13g2_and3_1 _22452_ (.X(_05312_),
    .A(\atari2600.pia.time_counter[3] ),
    .B(_05290_),
    .C(_05303_));
 sg13g2_nor3_1 _22453_ (.A(\atari2600.pia.time_counter[13] ),
    .B(\atari2600.pia.time_counter[12] ),
    .C(\atari2600.pia.time_counter[11] ),
    .Y(_05313_));
 sg13g2_nor4_1 _22454_ (.A(\atari2600.pia.time_counter[17] ),
    .B(\atari2600.pia.time_counter[16] ),
    .C(\atari2600.pia.time_counter[15] ),
    .D(\atari2600.pia.time_counter[14] ),
    .Y(_05314_));
 sg13g2_xor2_1 _22455_ (.B(\atari2600.pia.time_counter[0] ),
    .A(\atari2600.pia.time_counter[1] ),
    .X(_05315_));
 sg13g2_nand4_1 _22456_ (.B(_05311_),
    .C(_05313_),
    .A(_05310_),
    .Y(_05316_),
    .D(_05314_));
 sg13g2_xnor2_1 _22457_ (.Y(_05317_),
    .A(_00083_),
    .B(_05293_));
 sg13g2_o21ai_1 _22458_ (.B1(_05309_),
    .Y(_05318_),
    .A1(_00084_),
    .A2(_05297_));
 sg13g2_nor2_1 _22459_ (.A(_05315_),
    .B(_05318_),
    .Y(_05319_));
 sg13g2_nor3_1 _22460_ (.A(_05304_),
    .B(_05306_),
    .C(_05316_),
    .Y(_05320_));
 sg13g2_nand4_1 _22461_ (.B(_05317_),
    .C(_05319_),
    .A(_05296_),
    .Y(_05321_),
    .D(_05320_));
 sg13g2_nor4_1 _22462_ (.A(_05299_),
    .B(_05302_),
    .C(_05312_),
    .D(_05321_),
    .Y(_05322_));
 sg13g2_nand2b_2 _22463_ (.Y(_05323_),
    .B(_05286_),
    .A_N(net5874));
 sg13g2_a21oi_1 _22464_ (.A1(net5844),
    .A2(_05323_),
    .Y(_05324_),
    .B1(net6526));
 sg13g2_a21o_2 _22465_ (.A2(_05323_),
    .A1(net5844),
    .B1(net6525),
    .X(_05325_));
 sg13g2_nand2_1 _22466_ (.Y(_05326_),
    .A(net7270),
    .B(net5812));
 sg13g2_nand3_1 _22467_ (.B(net5844),
    .C(_05323_),
    .A(net6548),
    .Y(_05327_));
 sg13g2_mux2_2 _22468_ (.A0(\atari2600.pia.reset_timer[0] ),
    .A1(net7270),
    .S(net5873),
    .X(_05328_));
 sg13g2_o21ai_1 _22469_ (.B1(_05326_),
    .Y(_00857_),
    .A1(_05327_),
    .A2(_05328_));
 sg13g2_nand2_1 _22470_ (.Y(_05329_),
    .A(net7276),
    .B(net5812));
 sg13g2_mux2_1 _22471_ (.A0(\atari2600.pia.reset_timer[1] ),
    .A1(\atari2600.pia.diag[1] ),
    .S(net5873),
    .X(_05330_));
 sg13g2_nor2_1 _22472_ (.A(_05328_),
    .B(_05330_),
    .Y(_05331_));
 sg13g2_xor2_1 _22473_ (.B(_05330_),
    .A(_05328_),
    .X(_05332_));
 sg13g2_o21ai_1 _22474_ (.B1(_05329_),
    .Y(_00858_),
    .A1(_05327_),
    .A2(_05332_));
 sg13g2_nand2_1 _22475_ (.Y(_05333_),
    .A(net7313),
    .B(net5812));
 sg13g2_mux2_1 _22476_ (.A0(\atari2600.pia.reset_timer[2] ),
    .A1(\atari2600.pia.diag[2] ),
    .S(net5874),
    .X(_05334_));
 sg13g2_nor3_1 _22477_ (.A(_05328_),
    .B(_05330_),
    .C(_05334_),
    .Y(_05335_));
 sg13g2_xnor2_1 _22478_ (.Y(_05336_),
    .A(_05331_),
    .B(_05334_));
 sg13g2_o21ai_1 _22479_ (.B1(_05333_),
    .Y(_00859_),
    .A1(_05327_),
    .A2(_05336_));
 sg13g2_nand2_1 _22480_ (.Y(_05337_),
    .A(net7108),
    .B(net5812));
 sg13g2_mux2_1 _22481_ (.A0(\atari2600.pia.reset_timer[3] ),
    .A1(\atari2600.pia.diag[3] ),
    .S(net5873),
    .X(_05338_));
 sg13g2_nor2b_1 _22482_ (.A(_05338_),
    .B_N(_05335_),
    .Y(_05339_));
 sg13g2_xnor2_1 _22483_ (.Y(_05340_),
    .A(_05335_),
    .B(_05338_));
 sg13g2_o21ai_1 _22484_ (.B1(_05337_),
    .Y(_00860_),
    .A1(_05327_),
    .A2(_05340_));
 sg13g2_nand2_1 _22485_ (.Y(_05341_),
    .A(net7274),
    .B(net5812));
 sg13g2_mux2_1 _22486_ (.A0(\atari2600.pia.reset_timer[4] ),
    .A1(\atari2600.pia.diag[4] ),
    .S(net5873),
    .X(_05342_));
 sg13g2_nand2b_1 _22487_ (.Y(_05343_),
    .B(_05339_),
    .A_N(_05342_));
 sg13g2_xnor2_1 _22488_ (.Y(_05344_),
    .A(_05339_),
    .B(_05342_));
 sg13g2_o21ai_1 _22489_ (.B1(_05341_),
    .Y(_00861_),
    .A1(_05327_),
    .A2(_05344_));
 sg13g2_nand2_1 _22490_ (.Y(_05345_),
    .A(net7159),
    .B(net5812));
 sg13g2_nor2_1 _22491_ (.A(\atari2600.pia.reset_timer[5] ),
    .B(net5873),
    .Y(_05346_));
 sg13g2_a21oi_1 _22492_ (.A1(_08567_),
    .A2(net5873),
    .Y(_05347_),
    .B1(_05346_));
 sg13g2_or2_1 _22493_ (.X(_05348_),
    .B(_05347_),
    .A(_05343_));
 sg13g2_xor2_1 _22494_ (.B(_05347_),
    .A(_05343_),
    .X(_05349_));
 sg13g2_o21ai_1 _22495_ (.B1(_05345_),
    .Y(_00862_),
    .A1(_05327_),
    .A2(_05349_));
 sg13g2_nand2_1 _22496_ (.Y(_05350_),
    .A(net7277),
    .B(net5812));
 sg13g2_mux2_1 _22497_ (.A0(\atari2600.pia.reset_timer[6] ),
    .A1(\atari2600.pia.diag[6] ),
    .S(net5873),
    .X(_05351_));
 sg13g2_nor2_1 _22498_ (.A(_05348_),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_xor2_1 _22499_ (.B(_05351_),
    .A(_05348_),
    .X(_05353_));
 sg13g2_o21ai_1 _22500_ (.B1(_05350_),
    .Y(_00863_),
    .A1(_05327_),
    .A2(_05353_));
 sg13g2_nand2_1 _22501_ (.Y(_05354_),
    .A(net7283),
    .B(net5812));
 sg13g2_mux2_1 _22502_ (.A0(net4467),
    .A1(\atari2600.pia.diag[7] ),
    .S(net5874),
    .X(_05355_));
 sg13g2_xnor2_1 _22503_ (.Y(_05356_),
    .A(_05352_),
    .B(_05355_));
 sg13g2_o21ai_1 _22504_ (.B1(_05354_),
    .Y(_00864_),
    .A1(_05327_),
    .A2(_05356_));
 sg13g2_nand2_1 _22505_ (.Y(_05357_),
    .A(_05282_),
    .B(_05287_));
 sg13g2_a21oi_1 _22506_ (.A1(net5844),
    .A2(_05287_),
    .Y(_05358_),
    .B1(net6525));
 sg13g2_nand2_2 _22507_ (.Y(_05359_),
    .A(net6547),
    .B(_05357_));
 sg13g2_nand2_1 _22508_ (.Y(_05360_),
    .A(net3726),
    .B(net5809));
 sg13g2_nor4_1 _22509_ (.A(net7313),
    .B(net7276),
    .C(net7270),
    .D(net6527),
    .Y(_05361_));
 sg13g2_nor4_1 _22510_ (.A(net7283),
    .B(net7277),
    .C(net7274),
    .D(net7108),
    .Y(_05362_));
 sg13g2_nand4_1 _22511_ (.B(net5873),
    .C(_05361_),
    .A(_08567_),
    .Y(_05363_),
    .D(_05362_));
 sg13g2_o21ai_1 _22512_ (.B1(_05360_),
    .Y(_00865_),
    .A1(_05283_),
    .A2(_05363_));
 sg13g2_and2_1 _22513_ (.A(_09277_),
    .B(_03025_),
    .X(_05364_));
 sg13g2_nor2_1 _22514_ (.A(net6532),
    .B(_08712_),
    .Y(_05365_));
 sg13g2_nand2_2 _22515_ (.Y(_05366_),
    .A(net6576),
    .B(net5913));
 sg13g2_nand2_1 _22516_ (.Y(_05367_),
    .A(net5274),
    .B(net5808));
 sg13g2_nor2_1 _22517_ (.A(_09113_),
    .B(net5247),
    .Y(_05368_));
 sg13g2_and3_1 _22518_ (.X(_05369_),
    .A(_09303_),
    .B(_09413_),
    .C(_05368_));
 sg13g2_nand2b_1 _22519_ (.Y(_05370_),
    .B(_09337_),
    .A_N(_04683_));
 sg13g2_and2_1 _22520_ (.A(_05369_),
    .B(_05370_),
    .X(_05371_));
 sg13g2_a21oi_1 _22521_ (.A1(\gamepad_pmod.decoder.data_reg[8] ),
    .A2(_04681_),
    .Y(_05372_),
    .B1(_04676_));
 sg13g2_o21ai_1 _22522_ (.B1(_03072_),
    .Y(_05373_),
    .A1(net8),
    .A2(_05372_));
 sg13g2_nor2_2 _22523_ (.A(net5432),
    .B(net5506),
    .Y(_05374_));
 sg13g2_and2_2 _22524_ (.A(_09329_),
    .B(_05374_),
    .X(_05375_));
 sg13g2_nor2_2 _22525_ (.A(_09212_),
    .B(_09330_),
    .Y(_05376_));
 sg13g2_a22oi_1 _22526_ (.Y(_05377_),
    .B1(net5134),
    .B2(net7270),
    .A2(_05375_),
    .A1(net3234));
 sg13g2_nand3_1 _22527_ (.B(_05373_),
    .C(_05377_),
    .A(_05371_),
    .Y(_05378_));
 sg13g2_nand3_1 _22528_ (.B(_09338_),
    .C(_09413_),
    .A(_09303_),
    .Y(_05379_));
 sg13g2_nor3_1 _22529_ (.A(_09113_),
    .B(_09414_),
    .C(net5247),
    .Y(_05380_));
 sg13g2_nand2_1 _22530_ (.Y(_05381_),
    .A(_09303_),
    .B(_05380_));
 sg13g2_o21ai_1 _22531_ (.B1(_05378_),
    .Y(_05382_),
    .A1(net7327),
    .A2(_05369_));
 sg13g2_inv_1 _22532_ (.Y(_00866_),
    .A(_05382_));
 sg13g2_nand3_1 _22533_ (.B(_04675_),
    .C(_04681_),
    .A(\gamepad_pmod.decoder.data_reg[9] ),
    .Y(_05383_));
 sg13g2_o21ai_1 _22534_ (.B1(_05383_),
    .Y(_05384_),
    .A1(net6),
    .A2(_04675_));
 sg13g2_nor2_1 _22535_ (.A(_03073_),
    .B(_05384_),
    .Y(_05385_));
 sg13g2_a221oi_1 _22536_ (.B2(\atari2600.pia.diag[1] ),
    .C1(_05385_),
    .B1(net5134),
    .A1(net4409),
    .Y(_05386_),
    .A2(_05375_));
 sg13g2_nand2b_1 _22537_ (.Y(_05387_),
    .B(_05379_),
    .A_N(_04688_));
 sg13g2_nor2b_1 _22538_ (.A(net4991),
    .B_N(_05387_),
    .Y(_05388_));
 sg13g2_a22oi_1 _22539_ (.Y(_00867_),
    .B1(_05386_),
    .B2(_05388_),
    .A2(net4991),
    .A1(_08663_));
 sg13g2_nor2_2 _22540_ (.A(net5203),
    .B(_09437_),
    .Y(_05389_));
 sg13g2_a21o_1 _22541_ (.A2(_05375_),
    .A1(net3288),
    .B1(_03072_),
    .X(_05390_));
 sg13g2_a221oi_1 _22542_ (.B2(net4191),
    .C1(_05390_),
    .B1(_05389_),
    .A1(\atari2600.pia.diag[2] ),
    .Y(_05391_),
    .A2(net5134));
 sg13g2_nand2b_1 _22543_ (.Y(_05392_),
    .B(_05379_),
    .A_N(_04691_));
 sg13g2_nor2b_1 _22544_ (.A(net4991),
    .B_N(_05392_),
    .Y(_05393_));
 sg13g2_a22oi_1 _22545_ (.Y(_00868_),
    .B1(_05391_),
    .B2(_05393_),
    .A2(net4991),
    .A1(_08664_));
 sg13g2_and2_1 _22546_ (.A(net4249),
    .B(_05375_),
    .X(_05394_));
 sg13g2_a221oi_1 _22547_ (.B2(net7108),
    .C1(_05394_),
    .B1(net5134),
    .A1(\atari2600.input_switches[2] ),
    .Y(_05395_),
    .A2(_03072_));
 sg13g2_nand2b_1 _22548_ (.Y(_05396_),
    .B(_09337_),
    .A_N(_04694_));
 sg13g2_and2_1 _22549_ (.A(_05369_),
    .B(_05396_),
    .X(_05397_));
 sg13g2_a22oi_1 _22550_ (.Y(_00869_),
    .B1(_05395_),
    .B2(_05397_),
    .A2(_05381_),
    .A1(_08665_));
 sg13g2_a21o_1 _22551_ (.A2(_05375_),
    .A1(net4089),
    .B1(_03072_),
    .X(_05398_));
 sg13g2_a221oi_1 _22552_ (.B2(net3199),
    .C1(_05398_),
    .B1(_05389_),
    .A1(\atari2600.pia.diag[4] ),
    .Y(_05399_),
    .A2(net5134));
 sg13g2_a22oi_1 _22553_ (.Y(_00870_),
    .B1(_05399_),
    .B2(_05371_),
    .A2(net4991),
    .A1(_08666_));
 sg13g2_a21o_1 _22554_ (.A2(_05389_),
    .A1(net3888),
    .B1(_03072_),
    .X(_05400_));
 sg13g2_a221oi_1 _22555_ (.B2(\atari2600.pia.diag[5] ),
    .C1(_05400_),
    .B1(net5134),
    .A1(net3709),
    .Y(_05401_),
    .A2(_05375_));
 sg13g2_a22oi_1 _22556_ (.Y(_00871_),
    .B1(_05388_),
    .B2(_05401_),
    .A2(net4991),
    .A1(_08667_));
 sg13g2_and2_1 _22557_ (.A(_09353_),
    .B(_09413_),
    .X(_05402_));
 sg13g2_nand2_1 _22558_ (.Y(_05403_),
    .A(\atari2600.pia.diag[6] ),
    .B(_05376_));
 sg13g2_o21ai_1 _22559_ (.B1(_05403_),
    .Y(_05404_),
    .A1(\atari2600.input_switches[0] ),
    .A2(_03073_));
 sg13g2_a221oi_1 _22560_ (.B2(net3121),
    .C1(_05404_),
    .B1(_05402_),
    .A1(net3230),
    .Y(_05405_),
    .A2(_05375_));
 sg13g2_a22oi_1 _22561_ (.Y(_00872_),
    .B1(_05393_),
    .B2(_05405_),
    .A2(net4991),
    .A1(_08668_));
 sg13g2_nand2_1 _22562_ (.Y(_05406_),
    .A(net3726),
    .B(_05402_));
 sg13g2_o21ai_1 _22563_ (.B1(_05406_),
    .Y(_05407_),
    .A1(\atari2600.input_switches[1] ),
    .A2(_03073_));
 sg13g2_a221oi_1 _22564_ (.B2(\atari2600.pia.diag[7] ),
    .C1(_05407_),
    .B1(net5134),
    .A1(\atari2600.pia.swa_dir[7] ),
    .Y(_05408_),
    .A2(_05375_));
 sg13g2_a22oi_1 _22565_ (.Y(_00873_),
    .B1(_05397_),
    .B2(_05408_),
    .A2(net4991),
    .A1(_08669_));
 sg13g2_nor2_2 _22566_ (.A(_05283_),
    .B(_05323_),
    .Y(_05409_));
 sg13g2_xnor2_1 _22567_ (.Y(_05410_),
    .A(net7405),
    .B(net5844));
 sg13g2_nor2_1 _22568_ (.A(_05325_),
    .B(_05410_),
    .Y(_00874_));
 sg13g2_a21oi_1 _22569_ (.A1(\atari2600.pia.time_counter[0] ),
    .A2(net5844),
    .Y(_05411_),
    .B1(net7348));
 sg13g2_and3_1 _22570_ (.X(_05412_),
    .A(\atari2600.pia.time_counter[1] ),
    .B(net7599),
    .C(net5844));
 sg13g2_nor3_1 _22571_ (.A(_05359_),
    .B(net7349),
    .C(_05412_),
    .Y(_00875_));
 sg13g2_o21ai_1 _22572_ (.B1(net5810),
    .Y(_05413_),
    .A1(net7294),
    .A2(_05412_));
 sg13g2_a21oi_1 _22573_ (.A1(net7294),
    .A2(_05412_),
    .Y(_00876_),
    .B1(_05413_));
 sg13g2_a21oi_1 _22574_ (.A1(\atari2600.pia.time_counter[2] ),
    .A2(_05412_),
    .Y(_05414_),
    .B1(net7184));
 sg13g2_and3_1 _22575_ (.X(_05415_),
    .A(net7184),
    .B(net7597),
    .C(_05412_));
 sg13g2_nor3_1 _22576_ (.A(_05325_),
    .B(net7185),
    .C(_05415_),
    .Y(_00877_));
 sg13g2_a21oi_1 _22577_ (.A1(net7414),
    .A2(_05415_),
    .Y(_05416_),
    .B1(_05359_));
 sg13g2_o21ai_1 _22578_ (.B1(_05416_),
    .Y(_05417_),
    .A1(net7414),
    .A2(_05415_));
 sg13g2_inv_1 _22579_ (.Y(_00878_),
    .A(net7415));
 sg13g2_a21oi_1 _22580_ (.A1(\atari2600.pia.time_counter[4] ),
    .A2(_05415_),
    .Y(_05418_),
    .B1(net4151));
 sg13g2_and4_1 _22581_ (.A(\atari2600.pia.time_counter[3] ),
    .B(\atari2600.pia.time_counter[2] ),
    .C(\atari2600.pia.time_counter[1] ),
    .D(\atari2600.pia.time_counter[0] ),
    .X(_05419_));
 sg13g2_and2_2 _22582_ (.A(_05300_),
    .B(_05419_),
    .X(_05420_));
 sg13g2_and2_1 _22583_ (.A(net5844),
    .B(_05420_),
    .X(_05421_));
 sg13g2_nor3_1 _22584_ (.A(_05359_),
    .B(net4152),
    .C(_05421_),
    .Y(_00879_));
 sg13g2_xnor2_1 _22585_ (.Y(_05422_),
    .A(_00083_),
    .B(_05420_));
 sg13g2_a22oi_1 _22586_ (.Y(_05423_),
    .B1(_05409_),
    .B2(_05422_),
    .A2(_05283_),
    .A1(net7343));
 sg13g2_nor2_1 _22587_ (.A(net6525),
    .B(net7344),
    .Y(_00880_));
 sg13g2_a21oi_1 _22588_ (.A1(\atari2600.pia.time_counter[6] ),
    .A2(_05421_),
    .Y(_05424_),
    .B1(net7337));
 sg13g2_and2_1 _22589_ (.A(\atari2600.pia.time_counter[7] ),
    .B(\atari2600.pia.time_counter[6] ),
    .X(_05425_));
 sg13g2_and3_1 _22590_ (.X(_05426_),
    .A(net7337),
    .B(\atari2600.pia.time_counter[6] ),
    .C(_05421_));
 sg13g2_nor3_1 _22591_ (.A(_05325_),
    .B(net7338),
    .C(_05426_),
    .Y(_00881_));
 sg13g2_o21ai_1 _22592_ (.B1(_05324_),
    .Y(_05427_),
    .A1(net7018),
    .A2(_05426_));
 sg13g2_a21oi_1 _22593_ (.A1(net7018),
    .A2(_05426_),
    .Y(_00882_),
    .B1(_05427_));
 sg13g2_and3_1 _22594_ (.X(_05428_),
    .A(_05295_),
    .B(_05420_),
    .C(_05425_));
 sg13g2_a21oi_1 _22595_ (.A1(_05420_),
    .A2(_05425_),
    .Y(_05429_),
    .B1(net7203));
 sg13g2_nor3_1 _22596_ (.A(_05294_),
    .B(_05428_),
    .C(_05429_),
    .Y(_05430_));
 sg13g2_and4_1 _22597_ (.A(\atari2600.pia.time_counter[7] ),
    .B(\atari2600.pia.time_counter[6] ),
    .C(_05295_),
    .D(_05420_),
    .X(_05431_));
 sg13g2_a22oi_1 _22598_ (.Y(_05432_),
    .B1(_05409_),
    .B2(_05430_),
    .A2(_05283_),
    .A1(net7203));
 sg13g2_nor2_1 _22599_ (.A(net6526),
    .B(_05432_),
    .Y(_00883_));
 sg13g2_xnor2_1 _22600_ (.Y(_05433_),
    .A(_00084_),
    .B(_05428_));
 sg13g2_a22oi_1 _22601_ (.Y(_05434_),
    .B1(_05409_),
    .B2(_05433_),
    .A2(_05283_),
    .A1(net4476));
 sg13g2_nor2_1 _22602_ (.A(net6525),
    .B(net4477),
    .Y(_00884_));
 sg13g2_nand3_1 _22603_ (.B(_05282_),
    .C(_05428_),
    .A(net4476),
    .Y(_05435_));
 sg13g2_nor2_1 _22604_ (.A(_08566_),
    .B(_05435_),
    .Y(_05436_));
 sg13g2_and4_1 _22605_ (.A(net7487),
    .B(net4476),
    .C(_05282_),
    .D(_05431_),
    .X(_05437_));
 sg13g2_a21oi_1 _22606_ (.A1(_08566_),
    .A2(_05435_),
    .Y(_05438_),
    .B1(_05325_));
 sg13g2_nor2b_1 _22607_ (.A(_05437_),
    .B_N(_05438_),
    .Y(_00885_));
 sg13g2_nor2_1 _22608_ (.A(net7207),
    .B(_05437_),
    .Y(_05439_));
 sg13g2_and2_1 _22609_ (.A(net7207),
    .B(_05436_),
    .X(_05440_));
 sg13g2_nor3_1 _22610_ (.A(_05359_),
    .B(net7208),
    .C(_05440_),
    .Y(_00886_));
 sg13g2_a21o_1 _22611_ (.A2(_05357_),
    .A1(net7549),
    .B1(_05440_),
    .X(_05441_));
 sg13g2_o21ai_1 _22612_ (.B1(_05440_),
    .Y(_05442_),
    .A1(net7549),
    .A2(_05287_));
 sg13g2_and3_1 _22613_ (.X(_00887_),
    .A(net6547),
    .B(_05441_),
    .C(_05442_));
 sg13g2_a21o_1 _22614_ (.A2(_05440_),
    .A1(\atari2600.pia.time_counter[13] ),
    .B1(net7490),
    .X(_05443_));
 sg13g2_nand4_1 _22615_ (.B(net7598),
    .C(net7207),
    .A(net7490),
    .Y(_05444_),
    .D(_05437_));
 sg13g2_and3_1 _22616_ (.X(_00888_),
    .A(net5811),
    .B(net7491),
    .C(_05444_));
 sg13g2_nand4_1 _22617_ (.B(\atari2600.pia.time_counter[14] ),
    .C(\atari2600.pia.time_counter[13] ),
    .A(net6597),
    .Y(_05445_),
    .D(_05440_));
 sg13g2_nand2_1 _22618_ (.Y(_05446_),
    .A(net5811),
    .B(_05445_));
 sg13g2_a21oi_1 _22619_ (.A1(_08565_),
    .A2(_05444_),
    .Y(_00889_),
    .B1(_05446_));
 sg13g2_nor3_1 _22620_ (.A(_08564_),
    .B(_08565_),
    .C(_05444_),
    .Y(_05447_));
 sg13g2_nand2b_1 _22621_ (.Y(_05448_),
    .B(net5811),
    .A_N(_05447_));
 sg13g2_a21oi_1 _22622_ (.A1(_08564_),
    .A2(_05445_),
    .Y(_00890_),
    .B1(_05448_));
 sg13g2_nand2_1 _22623_ (.Y(_05449_),
    .A(_08563_),
    .B(net6548));
 sg13g2_a21oi_1 _22624_ (.A1(_05286_),
    .A2(_05447_),
    .Y(_05450_),
    .B1(net4324));
 sg13g2_a21oi_1 _22625_ (.A1(_05448_),
    .A2(_05449_),
    .Y(_00891_),
    .B1(net4325));
 sg13g2_nor3_1 _22626_ (.A(_08563_),
    .B(_08564_),
    .C(_05445_),
    .Y(_05451_));
 sg13g2_and3_1 _22627_ (.X(_05452_),
    .A(net7391),
    .B(net4324),
    .C(_05447_));
 sg13g2_o21ai_1 _22628_ (.B1(net5811),
    .Y(_05453_),
    .A1(net7391),
    .A2(_05451_));
 sg13g2_nor2_1 _22629_ (.A(_05452_),
    .B(net7392),
    .Y(_00892_));
 sg13g2_and2_1 _22630_ (.A(net7353),
    .B(_05452_),
    .X(_05454_));
 sg13g2_o21ai_1 _22631_ (.B1(net5811),
    .Y(_05455_),
    .A1(net7353),
    .A2(_05452_));
 sg13g2_nor2_1 _22632_ (.A(_05454_),
    .B(net7354),
    .Y(_00893_));
 sg13g2_nor2_1 _22633_ (.A(net7104),
    .B(_05454_),
    .Y(_05456_));
 sg13g2_and4_1 _22634_ (.A(\atari2600.pia.time_counter[20] ),
    .B(\atari2600.pia.time_counter[19] ),
    .C(\atari2600.pia.time_counter[18] ),
    .D(_05451_),
    .X(_05457_));
 sg13g2_nand2b_1 _22635_ (.Y(_05458_),
    .B(net5811),
    .A_N(_05457_));
 sg13g2_nor2_1 _22636_ (.A(net7105),
    .B(_05458_),
    .Y(_00894_));
 sg13g2_nand2b_1 _22637_ (.Y(_05459_),
    .B(net6548),
    .A_N(net6612));
 sg13g2_a21oi_1 _22638_ (.A1(_05286_),
    .A2(_05457_),
    .Y(_05460_),
    .B1(net6612));
 sg13g2_a21oi_1 _22639_ (.A1(_05458_),
    .A2(_05459_),
    .Y(_00895_),
    .B1(net6613));
 sg13g2_a21oi_1 _22640_ (.A1(\atari2600.pia.time_counter[21] ),
    .A2(_05457_),
    .Y(_05461_),
    .B1(net3617));
 sg13g2_and3_1 _22641_ (.X(_05462_),
    .A(net3617),
    .B(net6612),
    .C(_05457_));
 sg13g2_nor3_1 _22642_ (.A(_05359_),
    .B(net3618),
    .C(_05462_),
    .Y(_00896_));
 sg13g2_a21oi_1 _22643_ (.A1(net7308),
    .A2(_05462_),
    .Y(_05463_),
    .B1(_05359_));
 sg13g2_o21ai_1 _22644_ (.B1(_05463_),
    .Y(_05464_),
    .A1(net7308),
    .A2(_05462_));
 sg13g2_inv_1 _22645_ (.Y(_00897_),
    .A(_05464_));
 sg13g2_nand3_1 _22646_ (.B(net5273),
    .C(net5808),
    .A(_09113_),
    .Y(_05465_));
 sg13g2_nor3_2 _22647_ (.A(net5517),
    .B(_09322_),
    .C(_05465_),
    .Y(_05466_));
 sg13g2_or3_1 _22648_ (.A(net5517),
    .B(_09322_),
    .C(_05465_),
    .X(_05467_));
 sg13g2_nand2_1 _22649_ (.Y(_05468_),
    .A(_05368_),
    .B(net5134));
 sg13g2_nand4_1 _22650_ (.B(net6547),
    .C(net5131),
    .A(net7400),
    .Y(_05469_),
    .D(_05468_));
 sg13g2_o21ai_1 _22651_ (.B1(_05469_),
    .Y(_00898_),
    .A1(_05283_),
    .A2(_05363_));
 sg13g2_nand2_1 _22652_ (.Y(_05470_),
    .A(net7243),
    .B(net6525));
 sg13g2_a21oi_1 _22653_ (.A1(net7243),
    .A2(_05367_),
    .Y(_05471_),
    .B1(_05466_));
 sg13g2_o21ai_1 _22654_ (.B1(net5809),
    .Y(_05472_),
    .A1(net5739),
    .A2(net5131));
 sg13g2_o21ai_1 _22655_ (.B1(_05470_),
    .Y(_00899_),
    .A1(_05471_),
    .A2(_05472_));
 sg13g2_nand2_1 _22656_ (.Y(_05473_),
    .A(net6525),
    .B(net7138));
 sg13g2_a21oi_1 _22657_ (.A1(net7138),
    .A2(_05367_),
    .Y(_05474_),
    .B1(_05466_));
 sg13g2_o21ai_1 _22658_ (.B1(net5810),
    .Y(_05475_),
    .A1(net5749),
    .A2(net5132));
 sg13g2_o21ai_1 _22659_ (.B1(_05473_),
    .Y(_00900_),
    .A1(_05474_),
    .A2(_05475_));
 sg13g2_nand2_1 _22660_ (.Y(_05476_),
    .A(net6527),
    .B(net7124));
 sg13g2_a21oi_1 _22661_ (.A1(net7124),
    .A2(net5247),
    .Y(_05477_),
    .B1(net5133));
 sg13g2_o21ai_1 _22662_ (.B1(net5809),
    .Y(_05478_),
    .A1(net5621),
    .A2(net5131));
 sg13g2_o21ai_1 _22663_ (.B1(_05476_),
    .Y(_00901_),
    .A1(_05477_),
    .A2(_05478_));
 sg13g2_nand2_1 _22664_ (.Y(_05479_),
    .A(net6525),
    .B(net4735));
 sg13g2_a21oi_1 _22665_ (.A1(net4735),
    .A2(net5247),
    .Y(_05480_),
    .B1(net5133));
 sg13g2_o21ai_1 _22666_ (.B1(net5810),
    .Y(_05481_),
    .A1(net5615),
    .A2(net5131));
 sg13g2_o21ai_1 _22667_ (.B1(_05479_),
    .Y(_00902_),
    .A1(_05480_),
    .A2(_05481_));
 sg13g2_nand2_1 _22668_ (.Y(_05482_),
    .A(net6525),
    .B(net4960));
 sg13g2_a21oi_1 _22669_ (.A1(net4960),
    .A2(net5247),
    .Y(_05483_),
    .B1(net5133));
 sg13g2_o21ai_1 _22670_ (.B1(net5809),
    .Y(_05484_),
    .A1(net5606),
    .A2(net5131));
 sg13g2_o21ai_1 _22671_ (.B1(_05482_),
    .Y(_00903_),
    .A1(_05483_),
    .A2(_05484_));
 sg13g2_nand2_1 _22672_ (.Y(_05485_),
    .A(net6527),
    .B(net6941));
 sg13g2_a21oi_1 _22673_ (.A1(net6941),
    .A2(net5247),
    .Y(_05486_),
    .B1(net5133));
 sg13g2_o21ai_1 _22674_ (.B1(net5809),
    .Y(_05487_),
    .A1(net5580),
    .A2(net5131));
 sg13g2_o21ai_1 _22675_ (.B1(_05485_),
    .Y(_00904_),
    .A1(_05486_),
    .A2(_05487_));
 sg13g2_nand2_1 _22676_ (.Y(_05488_),
    .A(net6526),
    .B(net4504));
 sg13g2_a21oi_1 _22677_ (.A1(net4504),
    .A2(net5247),
    .Y(_05489_),
    .B1(net5133));
 sg13g2_o21ai_1 _22678_ (.B1(net5809),
    .Y(_05490_),
    .A1(net5575),
    .A2(net5131));
 sg13g2_o21ai_1 _22679_ (.B1(_05488_),
    .Y(_00905_),
    .A1(_05489_),
    .A2(_05490_));
 sg13g2_nand2_1 _22680_ (.Y(_05491_),
    .A(net6526),
    .B(net4467));
 sg13g2_a21oi_1 _22681_ (.A1(net4467),
    .A2(net5247),
    .Y(_05492_),
    .B1(net5133));
 sg13g2_o21ai_1 _22682_ (.B1(net5809),
    .Y(_05493_),
    .A1(net5642),
    .A2(net5131));
 sg13g2_o21ai_1 _22683_ (.B1(_05491_),
    .Y(_00906_),
    .A1(_05492_),
    .A2(_05493_));
 sg13g2_nor4_2 _22684_ (.A(net5432),
    .B(net5504),
    .C(_09330_),
    .Y(_05494_),
    .D(_05465_));
 sg13g2_nor2_1 _22685_ (.A(net3234),
    .B(net5129),
    .Y(_05495_));
 sg13g2_a21oi_1 _22686_ (.A1(net5763),
    .A2(net5129),
    .Y(_00907_),
    .B1(_05495_));
 sg13g2_nor2_1 _22687_ (.A(net4409),
    .B(_05494_),
    .Y(_05496_));
 sg13g2_a21oi_1 _22688_ (.A1(net5782),
    .A2(net5129),
    .Y(_00908_),
    .B1(_05496_));
 sg13g2_nor2_1 _22689_ (.A(net3288),
    .B(net5130),
    .Y(_05497_));
 sg13g2_a21oi_1 _22690_ (.A1(net5712),
    .A2(net5130),
    .Y(_00909_),
    .B1(_05497_));
 sg13g2_nor2_1 _22691_ (.A(net4249),
    .B(net5129),
    .Y(_05498_));
 sg13g2_a21oi_1 _22692_ (.A1(net5691),
    .A2(net5129),
    .Y(_00910_),
    .B1(_05498_));
 sg13g2_nor2_1 _22693_ (.A(net4089),
    .B(net5129),
    .Y(_05499_));
 sg13g2_a21oi_1 _22694_ (.A1(net5668),
    .A2(net5129),
    .Y(_00911_),
    .B1(_05499_));
 sg13g2_nor2_1 _22695_ (.A(net3709),
    .B(net5130),
    .Y(_05500_));
 sg13g2_a21oi_1 _22696_ (.A1(net5592),
    .A2(net5130),
    .Y(_00912_),
    .B1(_05500_));
 sg13g2_nor2_1 _22697_ (.A(net3230),
    .B(net5130),
    .Y(_05501_));
 sg13g2_a21oi_1 _22698_ (.A1(net5655),
    .A2(net5130),
    .Y(_00913_),
    .B1(_05501_));
 sg13g2_nor2_1 _22699_ (.A(net6989),
    .B(net5130),
    .Y(_05502_));
 sg13g2_a21oi_1 _22700_ (.A1(net5631),
    .A2(net5129),
    .Y(_00914_),
    .B1(_05502_));
 sg13g2_nor2_1 _22701_ (.A(net5533),
    .B(net5267),
    .Y(_05503_));
 sg13g2_nand2b_2 _22702_ (.Y(_05504_),
    .B(_09319_),
    .A_N(net5533));
 sg13g2_nor2_1 _22703_ (.A(net5339),
    .B(net5485),
    .Y(_05505_));
 sg13g2_nand2_2 _22704_ (.Y(_05506_),
    .A(net5368),
    .B(_09340_));
 sg13g2_nor2_1 _22705_ (.A(net5217),
    .B(_05506_),
    .Y(_05507_));
 sg13g2_nand2_2 _22706_ (.Y(_05508_),
    .A(net6551),
    .B(net5127));
 sg13g2_mux2_1 _22707_ (.A0(\atari2600.tia.diag[96] ),
    .A1(net7040),
    .S(_05508_),
    .X(_00915_));
 sg13g2_mux2_1 _22708_ (.A0(net6764),
    .A1(\atari2600.tia.old_grp1[1] ),
    .S(_05508_),
    .X(_00916_));
 sg13g2_mux2_1 _22709_ (.A0(\atari2600.tia.diag[98] ),
    .A1(net7139),
    .S(_05508_),
    .X(_00917_));
 sg13g2_mux2_1 _22710_ (.A0(\atari2600.tia.diag[99] ),
    .A1(net4941),
    .S(_05508_),
    .X(_00918_));
 sg13g2_mux2_1 _22711_ (.A0(\atari2600.tia.diag[100] ),
    .A1(net4525),
    .S(_05508_),
    .X(_00919_));
 sg13g2_mux2_1 _22712_ (.A0(net4346),
    .A1(\atari2600.tia.old_grp1[5] ),
    .S(_05508_),
    .X(_00920_));
 sg13g2_mux2_1 _22713_ (.A0(net4704),
    .A1(\atari2600.tia.old_grp1[6] ),
    .S(_05508_),
    .X(_00921_));
 sg13g2_mux2_1 _22714_ (.A0(net4574),
    .A1(\atari2600.tia.old_grp1[7] ),
    .S(_05508_),
    .X(_00922_));
 sg13g2_o21ai_1 _22715_ (.B1(_09213_),
    .Y(_05509_),
    .A1(_09202_),
    .A2(_09203_));
 sg13g2_nand3_1 _22716_ (.B(net6562),
    .C(_05509_),
    .A(net7440),
    .Y(_05510_));
 sg13g2_o21ai_1 _22717_ (.B1(_05510_),
    .Y(_00923_),
    .A1(_09201_),
    .A2(_09215_));
 sg13g2_nand3_1 _22718_ (.B(_09203_),
    .C(_09213_),
    .A(net6561),
    .Y(_05511_));
 sg13g2_nand3_1 _22719_ (.B(net6561),
    .C(_05509_),
    .A(net7416),
    .Y(_05512_));
 sg13g2_nand2_1 _22720_ (.Y(_00924_),
    .A(_05511_),
    .B(_05512_));
 sg13g2_nand3_1 _22721_ (.B(net5617),
    .C(net5772),
    .A(net5792),
    .Y(_05513_));
 sg13g2_nand3_1 _22722_ (.B(net6562),
    .C(_05509_),
    .A(net7318),
    .Y(_05514_));
 sg13g2_o21ai_1 _22723_ (.B1(_05514_),
    .Y(_00925_),
    .A1(_09215_),
    .A2(_05513_));
 sg13g2_nor2_1 _22724_ (.A(net5726),
    .B(net5776),
    .Y(_05515_));
 sg13g2_o21ai_1 _22725_ (.B1(net6553),
    .Y(_05516_),
    .A1(net7548),
    .A2(_09173_));
 sg13g2_a21oi_1 _22726_ (.A1(_09173_),
    .A2(_05515_),
    .Y(_00926_),
    .B1(_05516_));
 sg13g2_nor4_2 _22727_ (.A(net5080),
    .B(net5748),
    .C(net5726),
    .Y(_05517_),
    .D(net5776));
 sg13g2_a21o_1 _22728_ (.A2(net5079),
    .A1(net7460),
    .B1(_05517_),
    .X(_00927_));
 sg13g2_nor4_2 _22729_ (.A(net5080),
    .B(net5797),
    .C(net5726),
    .Y(_05518_),
    .D(net5776));
 sg13g2_a21o_1 _22730_ (.A2(net5079),
    .A1(net7515),
    .B1(_05518_),
    .X(_00928_));
 sg13g2_a21o_1 _22731_ (.A2(net5079),
    .A1(net6511),
    .B1(_05517_),
    .X(_00929_));
 sg13g2_a21o_1 _22732_ (.A2(net5079),
    .A1(net6510),
    .B1(_05518_),
    .X(_00930_));
 sg13g2_and2_1 _22733_ (.A(_09213_),
    .B(_05515_),
    .X(_05519_));
 sg13g2_a22oi_1 _22734_ (.Y(_05520_),
    .B1(_05519_),
    .B2(net5796),
    .A2(_09214_),
    .A1(net7471));
 sg13g2_nor2_1 _22735_ (.A(net6533),
    .B(_05520_),
    .Y(_00931_));
 sg13g2_and3_1 _22736_ (.X(_05521_),
    .A(net6550),
    .B(net5748),
    .C(_05519_));
 sg13g2_a21o_1 _22737_ (.A2(_09216_),
    .A1(net7489),
    .B1(_05521_),
    .X(_00932_));
 sg13g2_o21ai_1 _22738_ (.B1(net6561),
    .Y(_05522_),
    .A1(net7524),
    .A2(_09213_));
 sg13g2_nor2_1 _22739_ (.A(_05519_),
    .B(_05522_),
    .Y(_00933_));
 sg13g2_a22oi_1 _22740_ (.Y(_05523_),
    .B1(_05519_),
    .B2(net5796),
    .A2(_09214_),
    .A1(net7458));
 sg13g2_nor2_1 _22741_ (.A(net6533),
    .B(_05523_),
    .Y(_00934_));
 sg13g2_a21o_1 _22742_ (.A2(_09216_),
    .A1(net7479),
    .B1(_05521_),
    .X(_00935_));
 sg13g2_o21ai_1 _22743_ (.B1(net6547),
    .Y(_05524_),
    .A1(net7452),
    .A2(net5133));
 sg13g2_a21oi_1 _22744_ (.A1(net5432),
    .A2(net5133),
    .Y(_00936_),
    .B1(_05524_));
 sg13g2_nand3_1 _22745_ (.B(net6547),
    .C(net5132),
    .A(net4627),
    .Y(_05525_));
 sg13g2_o21ai_1 _22746_ (.B1(_05525_),
    .Y(_00937_),
    .A1(_09305_),
    .A2(net5132));
 sg13g2_nand3_1 _22747_ (.B(net6547),
    .C(net5132),
    .A(net3613),
    .Y(_05526_));
 sg13g2_o21ai_1 _22748_ (.B1(_05526_),
    .Y(_00938_),
    .A1(net5338),
    .A2(net5132));
 sg13g2_nand2_1 _22749_ (.Y(_05527_),
    .A(net4353),
    .B(_09205_));
 sg13g2_nand2_2 _22750_ (.Y(_05528_),
    .A(net5683),
    .B(net5599));
 sg13g2_o21ai_1 _22751_ (.B1(_05527_),
    .Y(_00939_),
    .A1(_09174_),
    .A2(_05528_));
 sg13g2_nand2_1 _22752_ (.Y(_05529_),
    .A(net6702),
    .B(_09205_));
 sg13g2_nand2_2 _22753_ (.Y(_05530_),
    .A(net5610),
    .B(net5598));
 sg13g2_o21ai_1 _22754_ (.B1(_05529_),
    .Y(_00940_),
    .A1(_09174_),
    .A2(_05530_));
 sg13g2_nand2_1 _22755_ (.Y(_05531_),
    .A(net4408),
    .B(net5079));
 sg13g2_nand2_2 _22756_ (.Y(_05532_),
    .A(net5683),
    .B(net5584));
 sg13g2_o21ai_1 _22757_ (.B1(_05531_),
    .Y(_00941_),
    .A1(net5080),
    .A2(_05532_));
 sg13g2_nand2_1 _22758_ (.Y(_05533_),
    .A(net4303),
    .B(net5079));
 sg13g2_nand2_2 _22759_ (.Y(_05534_),
    .A(net5610),
    .B(net5584));
 sg13g2_o21ai_1 _22760_ (.B1(_05533_),
    .Y(_00942_),
    .A1(net5080),
    .A2(_05534_));
 sg13g2_nand2_1 _22761_ (.Y(_05535_),
    .A(net4466),
    .B(_09216_));
 sg13g2_o21ai_1 _22762_ (.B1(_05535_),
    .Y(_00943_),
    .A1(_09215_),
    .A2(_05528_));
 sg13g2_nand2_1 _22763_ (.Y(_05536_),
    .A(net6879),
    .B(_09216_));
 sg13g2_o21ai_1 _22764_ (.B1(_05536_),
    .Y(_00944_),
    .A1(_09215_),
    .A2(_05530_));
 sg13g2_nand2_1 _22765_ (.Y(_05537_),
    .A(net4495),
    .B(_09216_));
 sg13g2_o21ai_1 _22766_ (.B1(_05537_),
    .Y(_00945_),
    .A1(_09215_),
    .A2(_05532_));
 sg13g2_nand2_1 _22767_ (.Y(_05538_),
    .A(net4418),
    .B(_09216_));
 sg13g2_o21ai_1 _22768_ (.B1(_05538_),
    .Y(_00946_),
    .A1(_09215_),
    .A2(_05534_));
 sg13g2_nor2_1 _22769_ (.A(net5246),
    .B(_09363_),
    .Y(_05539_));
 sg13g2_o21ai_1 _22770_ (.B1(net6565),
    .Y(_05540_),
    .A1(net7404),
    .A2(net5125));
 sg13g2_a21oi_1 _22771_ (.A1(_05528_),
    .A2(net5125),
    .Y(_00947_),
    .B1(_05540_));
 sg13g2_o21ai_1 _22772_ (.B1(net6565),
    .Y(_05541_),
    .A1(net7411),
    .A2(net5125));
 sg13g2_a21oi_1 _22773_ (.A1(_05530_),
    .A2(net5125),
    .Y(_00948_),
    .B1(_05541_));
 sg13g2_o21ai_1 _22774_ (.B1(net6565),
    .Y(_05542_),
    .A1(net7430),
    .A2(net5126));
 sg13g2_a21oi_1 _22775_ (.A1(_05532_),
    .A2(net5125),
    .Y(_00949_),
    .B1(_05542_));
 sg13g2_o21ai_1 _22776_ (.B1(net6565),
    .Y(_05543_),
    .A1(net7409),
    .A2(net5125));
 sg13g2_a21oi_1 _22777_ (.A1(_05534_),
    .A2(net5125),
    .Y(_00950_),
    .B1(_05543_));
 sg13g2_nor3_1 _22778_ (.A(net6245),
    .B(_00112_),
    .C(_11054_),
    .Y(_05544_));
 sg13g2_nand2b_1 _22779_ (.Y(_05545_),
    .B(_11055_),
    .A_N(_00112_));
 sg13g2_nor2_2 _22780_ (.A(net4988),
    .B(net5977),
    .Y(_05546_));
 sg13g2_a22oi_1 _22781_ (.Y(_05547_),
    .B1(_05546_),
    .B2(net2977),
    .A2(net4987),
    .A1(net5529));
 sg13g2_inv_1 _22782_ (.Y(_00951_),
    .A(_05547_));
 sg13g2_a22oi_1 _22783_ (.Y(_05548_),
    .B1(_05546_),
    .B2(net2985),
    .A2(net4988),
    .A1(net5564));
 sg13g2_inv_1 _22784_ (.Y(_00952_),
    .A(_05548_));
 sg13g2_a22oi_1 _22785_ (.Y(_05549_),
    .B1(_05546_),
    .B2(net2961),
    .A2(net4986),
    .A1(net5563));
 sg13g2_inv_1 _22786_ (.Y(_00953_),
    .A(_05549_));
 sg13g2_a22oi_1 _22787_ (.Y(_05550_),
    .B1(_05546_),
    .B2(net2978),
    .A2(net4986),
    .A1(net5556));
 sg13g2_inv_1 _22788_ (.Y(_00954_),
    .A(_05550_));
 sg13g2_or2_1 _22789_ (.X(_05551_),
    .B(net5977),
    .A(net7418));
 sg13g2_o21ai_1 _22790_ (.B1(_05551_),
    .Y(_05552_),
    .A1(net2977),
    .A2(net5947));
 sg13g2_o21ai_1 _22791_ (.B1(_03218_),
    .Y(_00955_),
    .A1(net4989),
    .A2(_05552_));
 sg13g2_mux2_1 _22792_ (.A0(net7401),
    .A1(net2985),
    .S(net5977),
    .X(_05553_));
 sg13g2_nand2_1 _22793_ (.Y(_05554_),
    .A(net4983),
    .B(_05553_));
 sg13g2_o21ai_1 _22794_ (.B1(_05554_),
    .Y(_00956_),
    .A1(net5570),
    .A2(net4983));
 sg13g2_or2_1 _22795_ (.X(_05555_),
    .B(net5978),
    .A(net7424));
 sg13g2_o21ai_1 _22796_ (.B1(_05555_),
    .Y(_05556_),
    .A1(net2961),
    .A2(net5947));
 sg13g2_o21ai_1 _22797_ (.B1(_03225_),
    .Y(_00957_),
    .A1(net4986),
    .A2(_05556_));
 sg13g2_or2_1 _22798_ (.X(_05557_),
    .B(net5976),
    .A(net7379));
 sg13g2_o21ai_1 _22799_ (.B1(_05557_),
    .Y(_05558_),
    .A1(net2978),
    .A2(net5946));
 sg13g2_o21ai_1 _22800_ (.B1(_03228_),
    .Y(_00958_),
    .A1(net4984),
    .A2(_05558_));
 sg13g2_mux2_1 _22801_ (.A0(net7497),
    .A1(net7418),
    .S(net5977),
    .X(_05559_));
 sg13g2_nand2_1 _22802_ (.Y(_05560_),
    .A(net4983),
    .B(_05559_));
 sg13g2_o21ai_1 _22803_ (.B1(_05560_),
    .Y(_00959_),
    .A1(_09272_),
    .A2(net4982));
 sg13g2_or2_1 _22804_ (.X(_05561_),
    .B(net5977),
    .A(net3256));
 sg13g2_o21ai_1 _22805_ (.B1(_05561_),
    .Y(_05562_),
    .A1(net7401),
    .A2(net5946));
 sg13g2_o21ai_1 _22806_ (.B1(_03234_),
    .Y(_00960_),
    .A1(net4988),
    .A2(_05562_));
 sg13g2_mux2_1 _22807_ (.A0(net7484),
    .A1(net7424),
    .S(net5978),
    .X(_05563_));
 sg13g2_nand2_1 _22808_ (.Y(_05564_),
    .A(net4982),
    .B(_05563_));
 sg13g2_o21ai_1 _22809_ (.B1(_05564_),
    .Y(_00961_),
    .A1(_09283_),
    .A2(net4982));
 sg13g2_or2_1 _22810_ (.X(_05565_),
    .B(net5976),
    .A(net7448));
 sg13g2_o21ai_1 _22811_ (.B1(_05565_),
    .Y(_05566_),
    .A1(net7379),
    .A2(net5946));
 sg13g2_o21ai_1 _22812_ (.B1(_03240_),
    .Y(_00962_),
    .A1(net4984),
    .A2(_05566_));
 sg13g2_nand2b_1 _22813_ (.Y(_05567_),
    .B(net5977),
    .A_N(net2989));
 sg13g2_o21ai_1 _22814_ (.B1(_05567_),
    .Y(_05568_),
    .A1(\flash_rom.addr[16] ),
    .A2(net5978));
 sg13g2_nand2_1 _22815_ (.Y(_05569_),
    .A(net2994),
    .B(net4988));
 sg13g2_o21ai_1 _22816_ (.B1(_05569_),
    .Y(_00963_),
    .A1(net4988),
    .A2(_05568_));
 sg13g2_nand2b_1 _22817_ (.Y(_05570_),
    .B(net5979),
    .A_N(\flash_rom.addr[13] ));
 sg13g2_o21ai_1 _22818_ (.B1(_05570_),
    .Y(_05571_),
    .A1(\flash_rom.addr[17] ),
    .A2(net5979));
 sg13g2_nand2_1 _22819_ (.Y(_05572_),
    .A(net4517),
    .B(net4989));
 sg13g2_o21ai_1 _22820_ (.B1(_05572_),
    .Y(_00964_),
    .A1(net4988),
    .A2(_05571_));
 sg13g2_nand2b_1 _22821_ (.Y(_05573_),
    .B(net5978),
    .A_N(net3049));
 sg13g2_o21ai_1 _22822_ (.B1(_05573_),
    .Y(_05574_),
    .A1(\flash_rom.addr[18] ),
    .A2(net5978));
 sg13g2_nand2_1 _22823_ (.Y(_05575_),
    .A(net7194),
    .B(net4989));
 sg13g2_o21ai_1 _22824_ (.B1(_05575_),
    .Y(_00965_),
    .A1(net4985),
    .A2(_05574_));
 sg13g2_nand2b_1 _22825_ (.Y(_05576_),
    .B(net5979),
    .A_N(net3214));
 sg13g2_o21ai_1 _22826_ (.B1(_05576_),
    .Y(_05577_),
    .A1(\flash_rom.addr[19] ),
    .A2(net5976));
 sg13g2_nand2_1 _22827_ (.Y(_05578_),
    .A(net4425),
    .B(net4984));
 sg13g2_o21ai_1 _22828_ (.B1(_05578_),
    .Y(_00966_),
    .A1(net4984),
    .A2(_05577_));
 sg13g2_nor2_1 _22829_ (.A(net5263),
    .B(net5255),
    .Y(_05579_));
 sg13g2_nor2_1 _22830_ (.A(net3921),
    .B(net5216),
    .Y(_05580_));
 sg13g2_a21oi_1 _22831_ (.A1(net5764),
    .A2(net5216),
    .Y(_00967_),
    .B1(_05580_));
 sg13g2_nor2_1 _22832_ (.A(net3097),
    .B(net5216),
    .Y(_05581_));
 sg13g2_a21oi_1 _22833_ (.A1(net5784),
    .A2(net5216),
    .Y(_00968_),
    .B1(_05581_));
 sg13g2_nor2_1 _22834_ (.A(net4390),
    .B(net5216),
    .Y(_05582_));
 sg13g2_a21oi_1 _22835_ (.A1(net5714),
    .A2(net5216),
    .Y(_00969_),
    .B1(_05582_));
 sg13g2_nor2_1 _22836_ (.A(net3022),
    .B(net5215),
    .Y(_05583_));
 sg13g2_a21oi_1 _22837_ (.A1(net5688),
    .A2(net5215),
    .Y(_00970_),
    .B1(_05583_));
 sg13g2_nor2_1 _22838_ (.A(net3276),
    .B(net5215),
    .Y(_05584_));
 sg13g2_a21oi_1 _22839_ (.A1(net5671),
    .A2(net5215),
    .Y(_00971_),
    .B1(_05584_));
 sg13g2_nor2_1 _22840_ (.A(net3475),
    .B(net5215),
    .Y(_05585_));
 sg13g2_a21oi_1 _22841_ (.A1(net5586),
    .A2(net5215),
    .Y(_00972_),
    .B1(_05585_));
 sg13g2_nor2_1 _22842_ (.A(net3794),
    .B(net5216),
    .Y(_05586_));
 sg13g2_a21oi_1 _22843_ (.A1(net5654),
    .A2(net5216),
    .Y(_00973_),
    .B1(_05586_));
 sg13g2_nor2_1 _22844_ (.A(net3299),
    .B(net5215),
    .Y(_05587_));
 sg13g2_a21oi_1 _22845_ (.A1(net5623),
    .A2(net5215),
    .Y(_00974_),
    .B1(_05587_));
 sg13g2_nand2_1 _22846_ (.Y(_05588_),
    .A(net2989),
    .B(net5947));
 sg13g2_nand2_1 _22847_ (.Y(_05589_),
    .A(\flash_rom.addr[8] ),
    .B(net5977));
 sg13g2_a21oi_1 _22848_ (.A1(_05588_),
    .A2(_05589_),
    .Y(_00975_),
    .B1(net4988));
 sg13g2_nand2_1 _22849_ (.Y(_05590_),
    .A(\flash_rom.addr[13] ),
    .B(net5947));
 sg13g2_nand2_1 _22850_ (.Y(_05591_),
    .A(net3256),
    .B(net5977));
 sg13g2_a21oi_1 _22851_ (.A1(_05590_),
    .A2(_05591_),
    .Y(_00976_),
    .B1(net4989));
 sg13g2_nand2_1 _22852_ (.Y(_05592_),
    .A(net3049),
    .B(net5946));
 sg13g2_nand2_1 _22853_ (.Y(_05593_),
    .A(\flash_rom.addr[10] ),
    .B(net5978));
 sg13g2_a21oi_1 _22854_ (.A1(_05592_),
    .A2(_05593_),
    .Y(_00977_),
    .B1(net4984));
 sg13g2_nand2_1 _22855_ (.Y(_05594_),
    .A(net3214),
    .B(net5946));
 sg13g2_nand2_1 _22856_ (.Y(_05595_),
    .A(\flash_rom.addr[11] ),
    .B(net5976));
 sg13g2_a21oi_1 _22857_ (.A1(_05594_),
    .A2(_05595_),
    .Y(_00978_),
    .B1(net4984));
 sg13g2_nand2_1 _22858_ (.Y(_05596_),
    .A(net7236),
    .B(net5978));
 sg13g2_nand2_1 _22859_ (.Y(_05597_),
    .A(\flash_rom.addr[20] ),
    .B(net5946));
 sg13g2_nand3_1 _22860_ (.B(_05596_),
    .C(_05597_),
    .A(net4982),
    .Y(_00979_));
 sg13g2_nor2_1 _22861_ (.A(\flash_rom.addr[17] ),
    .B(net5947),
    .Y(_05598_));
 sg13g2_nor2_1 _22862_ (.A(net3939),
    .B(net5976),
    .Y(_05599_));
 sg13g2_nor3_1 _22863_ (.A(net4985),
    .B(_05598_),
    .C(_05599_),
    .Y(_00980_));
 sg13g2_nor2_1 _22864_ (.A(\flash_rom.addr[18] ),
    .B(net5946),
    .Y(_05600_));
 sg13g2_nor2_1 _22865_ (.A(net4433),
    .B(net5976),
    .Y(_05601_));
 sg13g2_nor3_1 _22866_ (.A(net4985),
    .B(_05600_),
    .C(_05601_),
    .Y(_00981_));
 sg13g2_nor2_1 _22867_ (.A(\flash_rom.addr[19] ),
    .B(net5946),
    .Y(_05602_));
 sg13g2_nor2_1 _22868_ (.A(net3746),
    .B(net5976),
    .Y(_05603_));
 sg13g2_nor3_1 _22869_ (.A(net4985),
    .B(_05602_),
    .C(_05603_),
    .Y(_00982_));
 sg13g2_nor2_1 _22870_ (.A(_09441_),
    .B(net5256),
    .Y(_05604_));
 sg13g2_nor2_1 _22871_ (.A(net3723),
    .B(net5058),
    .Y(_05605_));
 sg13g2_a21oi_1 _22872_ (.A1(net5768),
    .A2(net5058),
    .Y(_00983_),
    .B1(_05605_));
 sg13g2_nor2_1 _22873_ (.A(net3126),
    .B(net5059),
    .Y(_05606_));
 sg13g2_a21oi_1 _22874_ (.A1(net5788),
    .A2(_05604_),
    .Y(_00984_),
    .B1(_05606_));
 sg13g2_nor2_1 _22875_ (.A(net3870),
    .B(net5058),
    .Y(_05607_));
 sg13g2_a21oi_1 _22876_ (.A1(net5718),
    .A2(net5058),
    .Y(_00985_),
    .B1(_05607_));
 sg13g2_nor2_1 _22877_ (.A(net3752),
    .B(net5058),
    .Y(_05608_));
 sg13g2_a21oi_1 _22878_ (.A1(net5695),
    .A2(net5058),
    .Y(_00986_),
    .B1(_05608_));
 sg13g2_nor2_1 _22879_ (.A(net3360),
    .B(net5058),
    .Y(_05609_));
 sg13g2_a21oi_1 _22880_ (.A1(net5675),
    .A2(net5058),
    .Y(_00987_),
    .B1(_05609_));
 sg13g2_nor2_1 _22881_ (.A(net4298),
    .B(net5059),
    .Y(_05610_));
 sg13g2_a21oi_1 _22882_ (.A1(net5593),
    .A2(net5059),
    .Y(_00988_),
    .B1(_05610_));
 sg13g2_nor2_1 _22883_ (.A(net3784),
    .B(net5059),
    .Y(_05611_));
 sg13g2_a21oi_1 _22884_ (.A1(net5655),
    .A2(net5059),
    .Y(_00989_),
    .B1(_05611_));
 sg13g2_nor2_1 _22885_ (.A(net3200),
    .B(net5059),
    .Y(_05612_));
 sg13g2_a21oi_1 _22886_ (.A1(net5636),
    .A2(net5059),
    .Y(_00990_),
    .B1(_05612_));
 sg13g2_nor2_2 _22887_ (.A(net6541),
    .B(net5913),
    .Y(_05613_));
 sg13g2_nand2_1 _22888_ (.Y(_05614_),
    .A(\atari2600.tia.audio_left_counter[0] ),
    .B(net5838));
 sg13g2_nor2_1 _22889_ (.A(_08509_),
    .B(\atari2600.tia.audc0[0] ),
    .Y(_05615_));
 sg13g2_nand2_1 _22890_ (.Y(_05616_),
    .A(\atari2600.tia.audc0[1] ),
    .B(_08510_));
 sg13g2_and2_1 _22891_ (.A(net6260),
    .B(net6261),
    .X(_05617_));
 sg13g2_nand3_1 _22892_ (.B(\atari2600.tia.audf0[1] ),
    .C(net6261),
    .A(\atari2600.tia.audf0[2] ),
    .Y(_05618_));
 sg13g2_or2_1 _22893_ (.X(_05619_),
    .B(_05618_),
    .A(_08502_));
 sg13g2_inv_1 _22894_ (.Y(_05620_),
    .A(_05619_));
 sg13g2_xor2_1 _22895_ (.B(_05619_),
    .A(_00101_),
    .X(_05621_));
 sg13g2_xnor2_1 _22896_ (.Y(_05622_),
    .A(_08502_),
    .B(_05618_));
 sg13g2_nor2_1 _22897_ (.A(_00101_),
    .B(_05622_),
    .Y(_05623_));
 sg13g2_nor4_2 _22898_ (.A(_08502_),
    .B(\atari2600.tia.audf0[2] ),
    .C(_08503_),
    .Y(_05624_),
    .D(\atari2600.tia.audf0[0] ));
 sg13g2_xor2_1 _22899_ (.B(net6261),
    .A(\atari2600.tia.audf0[1] ),
    .X(_05625_));
 sg13g2_and3_1 _22900_ (.X(_05626_),
    .A(_08502_),
    .B(net6260),
    .C(_05625_));
 sg13g2_nor2_1 _22901_ (.A(net6260),
    .B(\atari2600.tia.audf0[1] ),
    .Y(_05627_));
 sg13g2_a21oi_1 _22902_ (.A1(\atari2600.tia.audf0[1] ),
    .A2(net6261),
    .Y(_05628_),
    .B1(net6260));
 sg13g2_inv_1 _22903_ (.Y(_05629_),
    .A(_05628_));
 sg13g2_nand2_1 _22904_ (.Y(_05630_),
    .A(_05618_),
    .B(_05629_));
 sg13g2_a22oi_1 _22905_ (.Y(_05631_),
    .B1(_05628_),
    .B2(\atari2600.tia.audf0[3] ),
    .A2(_05617_),
    .A1(\atari2600.tia.audf0[1] ));
 sg13g2_xor2_1 _22906_ (.B(_05631_),
    .A(_00101_),
    .X(_05632_));
 sg13g2_nand2_1 _22907_ (.Y(_05633_),
    .A(_05626_),
    .B(_05632_));
 sg13g2_xnor2_1 _22908_ (.Y(_05634_),
    .A(_05626_),
    .B(_05632_));
 sg13g2_xnor2_1 _22909_ (.Y(_05635_),
    .A(_00096_),
    .B(_05634_));
 sg13g2_o21ai_1 _22910_ (.B1(_05633_),
    .Y(_05636_),
    .A1(_08618_),
    .A2(_05634_));
 sg13g2_a21oi_1 _22911_ (.A1(_00101_),
    .A2(_05629_),
    .Y(_05637_),
    .B1(_05622_));
 sg13g2_a21oi_1 _22912_ (.A1(_08502_),
    .A2(_00101_),
    .Y(_05638_),
    .B1(_05637_));
 sg13g2_nand2_1 _22913_ (.Y(_05639_),
    .A(_05625_),
    .B(_05638_));
 sg13g2_xor2_1 _22914_ (.B(_05638_),
    .A(_05625_),
    .X(_05640_));
 sg13g2_a22oi_1 _22915_ (.Y(_05641_),
    .B1(_05636_),
    .B2(_05640_),
    .A2(_05635_),
    .A1(_05624_));
 sg13g2_nand2b_1 _22916_ (.Y(_05642_),
    .B(_05623_),
    .A_N(_05641_));
 sg13g2_a21oi_1 _22917_ (.A1(\atari2600.tia.audf0[4] ),
    .A2(_05620_),
    .Y(_05643_),
    .B1(_05623_));
 sg13g2_nand3_1 _22918_ (.B(_05623_),
    .C(_05629_),
    .A(_05618_),
    .Y(_05644_));
 sg13g2_xnor2_1 _22919_ (.Y(_05645_),
    .A(_05630_),
    .B(_05643_));
 sg13g2_or2_1 _22920_ (.X(_05646_),
    .B(_05645_),
    .A(_05639_));
 sg13g2_o21ai_1 _22921_ (.B1(_05644_),
    .Y(_05647_),
    .A1(_05622_),
    .A2(_05646_));
 sg13g2_nand2b_1 _22922_ (.Y(_05648_),
    .B(_05642_),
    .A_N(_05647_));
 sg13g2_nand2_1 _22923_ (.Y(_05649_),
    .A(_05621_),
    .B(_05648_));
 sg13g2_o21ai_1 _22924_ (.B1(_05649_),
    .Y(_05650_),
    .A1(_00101_),
    .A2(_05619_));
 sg13g2_and2_1 _22925_ (.A(net6010),
    .B(_05650_),
    .X(_05651_));
 sg13g2_xor2_1 _22926_ (.B(_05648_),
    .A(_05621_),
    .X(_05652_));
 sg13g2_and2_2 _22927_ (.A(net6262),
    .B(net6263),
    .X(_05653_));
 sg13g2_nand2_2 _22928_ (.Y(_05654_),
    .A(net6262),
    .B(net6263));
 sg13g2_and2_1 _22929_ (.A(_05639_),
    .B(_05645_),
    .X(_05655_));
 sg13g2_xor2_1 _22930_ (.B(_05645_),
    .A(_05639_),
    .X(_05656_));
 sg13g2_xnor2_1 _22931_ (.Y(_05657_),
    .A(_05641_),
    .B(_05656_));
 sg13g2_nand2_1 _22932_ (.Y(_05658_),
    .A(net6010),
    .B(net5872));
 sg13g2_and2_1 _22933_ (.A(net6010),
    .B(_05652_),
    .X(_05659_));
 sg13g2_nand2_1 _22934_ (.Y(_05660_),
    .A(net6043),
    .B(_05659_));
 sg13g2_nand3_1 _22935_ (.B(net5872),
    .C(_05659_),
    .A(_05653_),
    .Y(_05661_));
 sg13g2_nor2_2 _22936_ (.A(net6262),
    .B(net6263),
    .Y(_05662_));
 sg13g2_nor2_1 _22937_ (.A(net6008),
    .B(_05662_),
    .Y(_05663_));
 sg13g2_nand2b_1 _22938_ (.Y(_05664_),
    .B(net6009),
    .A_N(_05662_));
 sg13g2_nand2_1 _22939_ (.Y(_05665_),
    .A(_05652_),
    .B(_05663_));
 sg13g2_o21ai_1 _22940_ (.B1(_05665_),
    .Y(_05666_),
    .A1(_05654_),
    .A2(_05658_));
 sg13g2_nand2_1 _22941_ (.Y(_05667_),
    .A(_05661_),
    .B(_05666_));
 sg13g2_or2_1 _22942_ (.X(_05668_),
    .B(_05640_),
    .A(_05636_));
 sg13g2_and2_1 _22943_ (.A(_05641_),
    .B(_05668_),
    .X(_05669_));
 sg13g2_nand2b_1 _22944_ (.Y(_05670_),
    .B(_05644_),
    .A_N(_05622_));
 sg13g2_o21ai_1 _22945_ (.B1(_05646_),
    .Y(_05671_),
    .A1(_05641_),
    .A2(_05655_));
 sg13g2_xnor2_1 _22946_ (.Y(_05672_),
    .A(_05670_),
    .B(_05671_));
 sg13g2_and2_1 _22947_ (.A(net6010),
    .B(_05672_),
    .X(_05673_));
 sg13g2_and3_1 _22948_ (.X(_05674_),
    .A(_05653_),
    .B(_05669_),
    .C(_05673_));
 sg13g2_nor2b_1 _22949_ (.A(_05667_),
    .B_N(_05674_),
    .Y(_05675_));
 sg13g2_and2_1 _22950_ (.A(net6010),
    .B(_05669_),
    .X(_05676_));
 sg13g2_xnor2_1 _22951_ (.Y(_05677_),
    .A(_05667_),
    .B(_05674_));
 sg13g2_xnor2_1 _22952_ (.Y(_05678_),
    .A(_05651_),
    .B(_05677_));
 sg13g2_xor2_1 _22953_ (.B(_05635_),
    .A(_05624_),
    .X(_05679_));
 sg13g2_nand2_1 _22954_ (.Y(_05680_),
    .A(net6010),
    .B(_05679_));
 sg13g2_nor2_1 _22955_ (.A(_05654_),
    .B(_05680_),
    .Y(_05681_));
 sg13g2_nand2_1 _22956_ (.Y(_05682_),
    .A(net5872),
    .B(_05681_));
 sg13g2_a22oi_1 _22957_ (.Y(_05683_),
    .B1(_05676_),
    .B2(net6043),
    .A2(_05672_),
    .A1(net5975));
 sg13g2_or2_1 _22958_ (.X(_05684_),
    .B(_05683_),
    .A(_05674_));
 sg13g2_or2_1 _22959_ (.X(_05685_),
    .B(_05684_),
    .A(_05682_));
 sg13g2_xnor2_1 _22960_ (.Y(_05686_),
    .A(_05682_),
    .B(_05684_));
 sg13g2_nand2_2 _22961_ (.Y(_05687_),
    .A(_05616_),
    .B(_05654_));
 sg13g2_a21oi_1 _22962_ (.A1(_05650_),
    .A2(_05687_),
    .Y(_05688_),
    .B1(_05659_));
 sg13g2_or2_1 _22963_ (.X(_05689_),
    .B(_05688_),
    .A(_05686_));
 sg13g2_a21o_1 _22964_ (.A2(_05689_),
    .A1(_05685_),
    .B1(_05678_),
    .X(_05690_));
 sg13g2_nand3_1 _22965_ (.B(_05685_),
    .C(_05689_),
    .A(_05678_),
    .Y(_05691_));
 sg13g2_nand2_1 _22966_ (.Y(_05692_),
    .A(_05690_),
    .B(_05691_));
 sg13g2_a21oi_1 _22967_ (.A1(net6260),
    .A2(_05625_),
    .Y(_05693_),
    .B1(_05627_));
 sg13g2_xnor2_1 _22968_ (.Y(_05694_),
    .A(\atari2600.tia.audf0[3] ),
    .B(_05693_));
 sg13g2_nor2_2 _22969_ (.A(net6008),
    .B(_05694_),
    .Y(_05695_));
 sg13g2_nand3_1 _22970_ (.B(net5871),
    .C(_05695_),
    .A(net6043),
    .Y(_05696_));
 sg13g2_inv_1 _22971_ (.Y(_05697_),
    .A(_05696_));
 sg13g2_a21oi_1 _22972_ (.A1(net5872),
    .A2(net5975),
    .Y(_05698_),
    .B1(_05681_));
 sg13g2_a21oi_1 _22973_ (.A1(net5872),
    .A2(_05681_),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_and2_1 _22974_ (.A(_05697_),
    .B(_05699_),
    .X(_05700_));
 sg13g2_nand2b_1 _22975_ (.Y(_05701_),
    .B(\atari2600.tia.audc0[1] ),
    .A_N(net6262));
 sg13g2_and3_1 _22976_ (.X(_05702_),
    .A(\atari2600.tia.audc0[2] ),
    .B(net6008),
    .C(_05701_));
 sg13g2_nand3_1 _22977_ (.B(net6008),
    .C(_05701_),
    .A(\atari2600.tia.audc0[2] ),
    .Y(_05703_));
 sg13g2_o21ai_1 _22978_ (.B1(net5974),
    .Y(_05704_),
    .A1(net6008),
    .A2(net6043));
 sg13g2_nand2_1 _22979_ (.Y(_05705_),
    .A(_05650_),
    .B(net5945));
 sg13g2_and2_1 _22980_ (.A(_05652_),
    .B(_05673_),
    .X(_05706_));
 sg13g2_o21ai_1 _22981_ (.B1(_05687_),
    .Y(_05707_),
    .A1(_05652_),
    .A2(_05673_));
 sg13g2_o21ai_1 _22982_ (.B1(_05705_),
    .Y(_05708_),
    .A1(_05706_),
    .A2(_05707_));
 sg13g2_xnor2_1 _22983_ (.Y(_05709_),
    .A(_05696_),
    .B(_05699_));
 sg13g2_a21oi_1 _22984_ (.A1(_05708_),
    .A2(_05709_),
    .Y(_05710_),
    .B1(_05700_));
 sg13g2_xnor2_1 _22985_ (.Y(_05711_),
    .A(_05686_),
    .B(_05688_));
 sg13g2_or2_1 _22986_ (.X(_05712_),
    .B(_05711_),
    .A(_05710_));
 sg13g2_xor2_1 _22987_ (.B(_05711_),
    .A(_05710_),
    .X(_05713_));
 sg13g2_nand2_1 _22988_ (.Y(_05714_),
    .A(_05706_),
    .B(_05713_));
 sg13g2_a21oi_1 _22989_ (.A1(_05712_),
    .A2(_05714_),
    .Y(_05715_),
    .B1(_05692_));
 sg13g2_inv_1 _22990_ (.Y(_05716_),
    .A(_05715_));
 sg13g2_a22oi_1 _22991_ (.Y(_05717_),
    .B1(_05673_),
    .B2(net6043),
    .A2(net5975),
    .A1(_05650_));
 sg13g2_nor2_1 _22992_ (.A(_05661_),
    .B(_05717_),
    .Y(_05718_));
 sg13g2_xor2_1 _22993_ (.B(_05717_),
    .A(_05661_),
    .X(_05719_));
 sg13g2_a21oi_1 _22994_ (.A1(_05651_),
    .A2(_05677_),
    .Y(_05720_),
    .B1(_05675_));
 sg13g2_nand2_2 _22995_ (.Y(_05721_),
    .A(_05719_),
    .B(_05720_));
 sg13g2_xor2_1 _22996_ (.B(_05721_),
    .A(_05690_),
    .X(_05722_));
 sg13g2_nor2_1 _22997_ (.A(_05716_),
    .B(_05721_),
    .Y(_05723_));
 sg13g2_or2_1 _22998_ (.X(_05724_),
    .B(_05722_),
    .A(_05715_));
 sg13g2_o21ai_1 _22999_ (.B1(_05724_),
    .Y(_05725_),
    .A1(_05716_),
    .A2(_05721_));
 sg13g2_xnor2_1 _23000_ (.Y(_05726_),
    .A(_05706_),
    .B(_05713_));
 sg13g2_xor2_1 _23001_ (.B(net6261),
    .A(net6260),
    .X(_05727_));
 sg13g2_xnor2_1 _23002_ (.Y(_05728_),
    .A(net6260),
    .B(net6261));
 sg13g2_nand2_1 _23003_ (.Y(_05729_),
    .A(net6009),
    .B(_05727_));
 sg13g2_nor2_2 _23004_ (.A(_05654_),
    .B(_05729_),
    .Y(_05730_));
 sg13g2_nand2_1 _23005_ (.Y(_05731_),
    .A(net5914),
    .B(_05730_));
 sg13g2_a22oi_1 _23006_ (.Y(_05732_),
    .B1(_05695_),
    .B2(net6043),
    .A2(net5871),
    .A1(net5975));
 sg13g2_or2_1 _23007_ (.X(_05733_),
    .B(_05732_),
    .A(_05697_));
 sg13g2_xnor2_1 _23008_ (.Y(_05734_),
    .A(_05731_),
    .B(_05733_));
 sg13g2_nand2_1 _23009_ (.Y(_05735_),
    .A(_05657_),
    .B(_05673_));
 sg13g2_xnor2_1 _23010_ (.Y(_05736_),
    .A(_05658_),
    .B(_05672_));
 sg13g2_nand2_1 _23011_ (.Y(_05737_),
    .A(_05687_),
    .B(_05736_));
 sg13g2_nand2_1 _23012_ (.Y(_05738_),
    .A(_05652_),
    .B(net5945));
 sg13g2_xor2_1 _23013_ (.B(_05738_),
    .A(_05737_),
    .X(_05739_));
 sg13g2_nand2b_1 _23014_ (.Y(_05740_),
    .B(_05739_),
    .A_N(_05734_));
 sg13g2_o21ai_1 _23015_ (.B1(_05740_),
    .Y(_05741_),
    .A1(_05731_),
    .A2(_05733_));
 sg13g2_xor2_1 _23016_ (.B(_05709_),
    .A(_05708_),
    .X(_05742_));
 sg13g2_o21ai_1 _23017_ (.B1(_05735_),
    .Y(_05743_),
    .A1(_05737_),
    .A2(_05738_));
 sg13g2_xnor2_1 _23018_ (.Y(_05744_),
    .A(_05741_),
    .B(_05742_));
 sg13g2_nor2b_1 _23019_ (.A(_05744_),
    .B_N(_05743_),
    .Y(_05745_));
 sg13g2_a21o_1 _23020_ (.A2(_05742_),
    .A1(_05741_),
    .B1(_05745_),
    .X(_05746_));
 sg13g2_nand2b_1 _23021_ (.Y(_05747_),
    .B(_05746_),
    .A_N(_05726_));
 sg13g2_nand3_1 _23022_ (.B(_05712_),
    .C(_05714_),
    .A(_05692_),
    .Y(_05748_));
 sg13g2_nand2_1 _23023_ (.Y(_05749_),
    .A(_05716_),
    .B(_05748_));
 sg13g2_or2_1 _23024_ (.X(_05750_),
    .B(_05749_),
    .A(_05747_));
 sg13g2_xnor2_1 _23025_ (.Y(_05751_),
    .A(_05743_),
    .B(_05744_));
 sg13g2_xnor2_1 _23026_ (.Y(_05752_),
    .A(_08618_),
    .B(_05625_));
 sg13g2_nand2_1 _23027_ (.Y(_05753_),
    .A(net6009),
    .B(net6007));
 sg13g2_nor2_1 _23028_ (.A(_05654_),
    .B(_05753_),
    .Y(_05754_));
 sg13g2_nor2_1 _23029_ (.A(_05664_),
    .B(_05694_),
    .Y(_05755_));
 sg13g2_and2_1 _23030_ (.A(_05695_),
    .B(_05754_),
    .X(_05756_));
 sg13g2_a21oi_1 _23031_ (.A1(net5975),
    .A2(_05679_),
    .Y(_05757_),
    .B1(_05730_));
 sg13g2_a21oi_1 _23032_ (.A1(net5914),
    .A2(_05730_),
    .Y(_05758_),
    .B1(_05757_));
 sg13g2_xnor2_1 _23033_ (.Y(_05759_),
    .A(_05756_),
    .B(_05758_));
 sg13g2_nand2_1 _23034_ (.Y(_05760_),
    .A(_05656_),
    .B(_05676_));
 sg13g2_a22oi_1 _23035_ (.Y(_05761_),
    .B1(_05687_),
    .B2(net5872),
    .A2(net5871),
    .A1(net6010));
 sg13g2_a21oi_1 _23036_ (.A1(_05656_),
    .A2(_05676_),
    .Y(_05762_),
    .B1(_05761_));
 sg13g2_nand2_1 _23037_ (.Y(_05763_),
    .A(_05672_),
    .B(net5945));
 sg13g2_xor2_1 _23038_ (.B(_05763_),
    .A(_05762_),
    .X(_05764_));
 sg13g2_nor2_1 _23039_ (.A(_05759_),
    .B(_05764_),
    .Y(_05765_));
 sg13g2_a21oi_1 _23040_ (.A1(_05756_),
    .A2(_05758_),
    .Y(_05766_),
    .B1(_05765_));
 sg13g2_xnor2_1 _23041_ (.Y(_05767_),
    .A(_05734_),
    .B(_05739_));
 sg13g2_nor2b_1 _23042_ (.A(_05766_),
    .B_N(_05767_),
    .Y(_05768_));
 sg13g2_o21ai_1 _23043_ (.B1(_05760_),
    .Y(_05769_),
    .A1(_05761_),
    .A2(_05763_));
 sg13g2_xnor2_1 _23044_ (.Y(_05770_),
    .A(_05766_),
    .B(_05767_));
 sg13g2_a21oi_1 _23045_ (.A1(_05769_),
    .A2(_05770_),
    .Y(_05771_),
    .B1(_05768_));
 sg13g2_nand2b_1 _23046_ (.Y(_05772_),
    .B(_05751_),
    .A_N(_05771_));
 sg13g2_xnor2_1 _23047_ (.Y(_05773_),
    .A(_05726_),
    .B(_05746_));
 sg13g2_nor2b_1 _23048_ (.A(_05772_),
    .B_N(_05773_),
    .Y(_05774_));
 sg13g2_xnor2_1 _23049_ (.Y(_05775_),
    .A(_05751_),
    .B(_05771_));
 sg13g2_xnor2_1 _23050_ (.Y(_05776_),
    .A(_05754_),
    .B(_05755_));
 sg13g2_nand2_1 _23051_ (.Y(_05777_),
    .A(_00096_),
    .B(_05730_));
 sg13g2_nor2_1 _23052_ (.A(_05776_),
    .B(_05777_),
    .Y(_05778_));
 sg13g2_xor2_1 _23053_ (.B(_05777_),
    .A(_05776_),
    .X(_05779_));
 sg13g2_nand2_1 _23054_ (.Y(_05780_),
    .A(_05676_),
    .B(net5914));
 sg13g2_nand3_1 _23055_ (.B(_05668_),
    .C(_05687_),
    .A(_05641_),
    .Y(_05781_));
 sg13g2_mux2_1 _23056_ (.A0(net5871),
    .A1(_05781_),
    .S(_05680_),
    .X(_05782_));
 sg13g2_nand2_1 _23057_ (.Y(_05783_),
    .A(net5872),
    .B(net5945));
 sg13g2_xor2_1 _23058_ (.B(_05783_),
    .A(_05782_),
    .X(_05784_));
 sg13g2_a21oi_1 _23059_ (.A1(_05779_),
    .A2(_05784_),
    .Y(_05785_),
    .B1(_05778_));
 sg13g2_xnor2_1 _23060_ (.Y(_05786_),
    .A(_05759_),
    .B(_05764_));
 sg13g2_nor2_1 _23061_ (.A(_05785_),
    .B(_05786_),
    .Y(_05787_));
 sg13g2_o21ai_1 _23062_ (.B1(_05780_),
    .Y(_05788_),
    .A1(_05782_),
    .A2(_05783_));
 sg13g2_xor2_1 _23063_ (.B(_05786_),
    .A(_05785_),
    .X(_05789_));
 sg13g2_a21oi_1 _23064_ (.A1(_05788_),
    .A2(_05789_),
    .Y(_05790_),
    .B1(_05787_));
 sg13g2_xnor2_1 _23065_ (.Y(_05791_),
    .A(_05769_),
    .B(_05770_));
 sg13g2_nor2_1 _23066_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sg13g2_and2_1 _23067_ (.A(_05650_),
    .B(_05703_),
    .X(_05793_));
 sg13g2_xor2_1 _23068_ (.B(_05791_),
    .A(_05790_),
    .X(_05794_));
 sg13g2_a21oi_1 _23069_ (.A1(_05793_),
    .A2(_05794_),
    .Y(_05795_),
    .B1(_05792_));
 sg13g2_nand2b_1 _23070_ (.Y(_05796_),
    .B(_05775_),
    .A_N(_05795_));
 sg13g2_nand3_1 _23071_ (.B(net6009),
    .C(net6043),
    .A(_00096_),
    .Y(_05797_));
 sg13g2_o21ai_1 _23072_ (.B1(_05797_),
    .Y(_05798_),
    .A1(_05664_),
    .A2(_05728_));
 sg13g2_nand2_1 _23073_ (.Y(_05799_),
    .A(_05777_),
    .B(_05798_));
 sg13g2_nand2_1 _23074_ (.Y(_05800_),
    .A(_05679_),
    .B(_05695_));
 sg13g2_a21o_1 _23075_ (.A2(_05687_),
    .A1(net5914),
    .B1(_05695_),
    .X(_05801_));
 sg13g2_a22oi_1 _23076_ (.Y(_05802_),
    .B1(_05800_),
    .B2(_05801_),
    .A2(net5945),
    .A1(net5871));
 sg13g2_and4_1 _23077_ (.A(net5871),
    .B(net5944),
    .C(_05800_),
    .D(_05801_),
    .X(_05803_));
 sg13g2_or3_2 _23078_ (.A(_05799_),
    .B(_05802_),
    .C(_05803_),
    .X(_05804_));
 sg13g2_xnor2_1 _23079_ (.Y(_05805_),
    .A(_05779_),
    .B(_05784_));
 sg13g2_nor2_1 _23080_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sg13g2_a21o_1 _23081_ (.A2(_05695_),
    .A1(net5914),
    .B1(_05803_),
    .X(_05807_));
 sg13g2_nand2_1 _23082_ (.Y(_05808_),
    .A(_05804_),
    .B(_05805_));
 sg13g2_xnor2_1 _23083_ (.Y(_05809_),
    .A(_05804_),
    .B(_05805_));
 sg13g2_a21oi_1 _23084_ (.A1(_05807_),
    .A2(_05808_),
    .Y(_05810_),
    .B1(_05806_));
 sg13g2_xnor2_1 _23085_ (.Y(_05811_),
    .A(_05788_),
    .B(_05789_));
 sg13g2_nor2_1 _23086_ (.A(_05810_),
    .B(_05811_),
    .Y(_05812_));
 sg13g2_nand2_1 _23087_ (.Y(_05813_),
    .A(_05652_),
    .B(_05703_));
 sg13g2_xor2_1 _23088_ (.B(_05811_),
    .A(_05810_),
    .X(_05814_));
 sg13g2_nor2b_1 _23089_ (.A(_05813_),
    .B_N(_05814_),
    .Y(_05815_));
 sg13g2_nor2_1 _23090_ (.A(_05812_),
    .B(_05815_),
    .Y(_05816_));
 sg13g2_xnor2_1 _23091_ (.Y(_05817_),
    .A(_05793_),
    .B(_05794_));
 sg13g2_nor2_1 _23092_ (.A(_05816_),
    .B(_05817_),
    .Y(_05818_));
 sg13g2_nand2_1 _23093_ (.Y(_05819_),
    .A(_05695_),
    .B(_05727_));
 sg13g2_a22oi_1 _23094_ (.Y(_05820_),
    .B1(_05694_),
    .B2(_05729_),
    .A2(_05654_),
    .A1(net6008));
 sg13g2_and2_1 _23095_ (.A(_05819_),
    .B(_05820_),
    .X(_05821_));
 sg13g2_a21o_1 _23096_ (.A2(net5944),
    .A1(net5914),
    .B1(_05821_),
    .X(_05822_));
 sg13g2_nand4_1 _23097_ (.B(net5944),
    .C(_05819_),
    .A(net5914),
    .Y(_05823_),
    .D(_05820_));
 sg13g2_and4_1 _23098_ (.A(net5975),
    .B(_05752_),
    .C(_05822_),
    .D(_05823_),
    .X(_05824_));
 sg13g2_o21ai_1 _23099_ (.B1(_05799_),
    .Y(_05825_),
    .A1(_05802_),
    .A2(_05803_));
 sg13g2_nand3_1 _23100_ (.B(_05824_),
    .C(_05825_),
    .A(_05804_),
    .Y(_05826_));
 sg13g2_nand2_1 _23101_ (.Y(_05827_),
    .A(_05819_),
    .B(_05823_));
 sg13g2_a21o_1 _23102_ (.A2(_05825_),
    .A1(_05804_),
    .B1(_05824_),
    .X(_05828_));
 sg13g2_nand3_1 _23103_ (.B(_05827_),
    .C(_05828_),
    .A(_05826_),
    .Y(_05829_));
 sg13g2_nand2_1 _23104_ (.Y(_05830_),
    .A(_05826_),
    .B(_05829_));
 sg13g2_xor2_1 _23105_ (.B(_05809_),
    .A(_05807_),
    .X(_05831_));
 sg13g2_nand2b_1 _23106_ (.Y(_05832_),
    .B(_05830_),
    .A_N(_05831_));
 sg13g2_nand2_1 _23107_ (.Y(_05833_),
    .A(_05672_),
    .B(_05703_));
 sg13g2_xor2_1 _23108_ (.B(_05831_),
    .A(_05830_),
    .X(_05834_));
 sg13g2_o21ai_1 _23109_ (.B1(_05832_),
    .Y(_05835_),
    .A1(_05833_),
    .A2(_05834_));
 sg13g2_xnor2_1 _23110_ (.Y(_05836_),
    .A(_05813_),
    .B(_05814_));
 sg13g2_nand2_1 _23111_ (.Y(_05837_),
    .A(_05835_),
    .B(_05836_));
 sg13g2_nand2_1 _23112_ (.Y(_05838_),
    .A(_00096_),
    .B(net5975));
 sg13g2_nand3_1 _23113_ (.B(_05727_),
    .C(net6007),
    .A(net6009),
    .Y(_05839_));
 sg13g2_nand2_1 _23114_ (.Y(_05840_),
    .A(_05728_),
    .B(_05753_));
 sg13g2_nand3_1 _23115_ (.B(_05839_),
    .C(_05840_),
    .A(_05687_),
    .Y(_05841_));
 sg13g2_nand2b_1 _23116_ (.Y(_05842_),
    .B(net5944),
    .A_N(_05694_));
 sg13g2_xor2_1 _23117_ (.B(_05842_),
    .A(_05841_),
    .X(_05843_));
 sg13g2_nand2b_1 _23118_ (.Y(_05844_),
    .B(_05843_),
    .A_N(_05838_));
 sg13g2_a22oi_1 _23119_ (.Y(_05845_),
    .B1(_05822_),
    .B2(_05823_),
    .A2(net6007),
    .A1(net5975));
 sg13g2_or3_1 _23120_ (.A(_05824_),
    .B(_05844_),
    .C(_05845_),
    .X(_05846_));
 sg13g2_o21ai_1 _23121_ (.B1(_05839_),
    .Y(_05847_),
    .A1(_05841_),
    .A2(_05842_));
 sg13g2_o21ai_1 _23122_ (.B1(_05844_),
    .Y(_05848_),
    .A1(_05824_),
    .A2(_05845_));
 sg13g2_and3_1 _23123_ (.X(_05849_),
    .A(_05846_),
    .B(_05847_),
    .C(_05848_));
 sg13g2_nand3_1 _23124_ (.B(_05847_),
    .C(_05848_),
    .A(_05846_),
    .Y(_05850_));
 sg13g2_nand2_1 _23125_ (.Y(_05851_),
    .A(_05846_),
    .B(_05850_));
 sg13g2_a21o_1 _23126_ (.A2(_05828_),
    .A1(_05826_),
    .B1(_05827_),
    .X(_05852_));
 sg13g2_nand3_1 _23127_ (.B(_05851_),
    .C(_05852_),
    .A(_05829_),
    .Y(_05853_));
 sg13g2_nand2_1 _23128_ (.Y(_05854_),
    .A(net5872),
    .B(net5974));
 sg13g2_inv_1 _23129_ (.Y(_05855_),
    .A(_05854_));
 sg13g2_a21o_1 _23130_ (.A2(_05852_),
    .A1(_05829_),
    .B1(_05851_),
    .X(_05856_));
 sg13g2_nand3_1 _23131_ (.B(_05855_),
    .C(_05856_),
    .A(_05853_),
    .Y(_05857_));
 sg13g2_nand2_1 _23132_ (.Y(_05858_),
    .A(_05853_),
    .B(_05857_));
 sg13g2_xor2_1 _23133_ (.B(_05834_),
    .A(_05833_),
    .X(_05859_));
 sg13g2_and2_1 _23134_ (.A(_05858_),
    .B(_05859_),
    .X(_05860_));
 sg13g2_xnor2_1 _23135_ (.Y(_05861_),
    .A(_05838_),
    .B(_05843_));
 sg13g2_nor2_1 _23136_ (.A(net6261),
    .B(_05753_),
    .Y(_05862_));
 sg13g2_nand3_1 _23137_ (.B(net6009),
    .C(net6007),
    .A(_08504_),
    .Y(_05863_));
 sg13g2_a22oi_1 _23138_ (.Y(_05864_),
    .B1(_05687_),
    .B2(net6007),
    .A2(net6009),
    .A1(_08504_));
 sg13g2_nor2_1 _23139_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sg13g2_nand2_1 _23140_ (.Y(_05866_),
    .A(net5944),
    .B(_05727_));
 sg13g2_o21ai_1 _23141_ (.B1(_05863_),
    .Y(_05867_),
    .A1(_05864_),
    .A2(_05866_));
 sg13g2_nand2_1 _23142_ (.Y(_05868_),
    .A(_05861_),
    .B(_05867_));
 sg13g2_a21oi_1 _23143_ (.A1(_05846_),
    .A2(_05848_),
    .Y(_05869_),
    .B1(_05847_));
 sg13g2_nor3_1 _23144_ (.A(_05849_),
    .B(_05868_),
    .C(_05869_),
    .Y(_05870_));
 sg13g2_or3_1 _23145_ (.A(_05849_),
    .B(_05868_),
    .C(_05869_),
    .X(_05871_));
 sg13g2_o21ai_1 _23146_ (.B1(_05868_),
    .Y(_05872_),
    .A1(_05849_),
    .A2(_05869_));
 sg13g2_and4_1 _23147_ (.A(net5871),
    .B(net5974),
    .C(_05871_),
    .D(_05872_),
    .X(_05873_));
 sg13g2_or2_1 _23148_ (.X(_05874_),
    .B(_05873_),
    .A(_05870_));
 sg13g2_a21o_1 _23149_ (.A2(_05856_),
    .A1(_05853_),
    .B1(_05855_),
    .X(_05875_));
 sg13g2_nand3_1 _23150_ (.B(_05874_),
    .C(_05875_),
    .A(_05857_),
    .Y(_05876_));
 sg13g2_a21oi_1 _23151_ (.A1(net6008),
    .A2(_05654_),
    .Y(_05877_),
    .B1(_08618_));
 sg13g2_nand3_1 _23152_ (.B(net6007),
    .C(_05877_),
    .A(net5944),
    .Y(_05878_));
 sg13g2_xor2_1 _23153_ (.B(_05866_),
    .A(_05865_),
    .X(_05879_));
 sg13g2_or2_1 _23154_ (.X(_05880_),
    .B(_05879_),
    .A(_05878_));
 sg13g2_inv_1 _23155_ (.Y(_05881_),
    .A(_05880_));
 sg13g2_xor2_1 _23156_ (.B(_05867_),
    .A(_05861_),
    .X(_05882_));
 sg13g2_nand2_1 _23157_ (.Y(_05883_),
    .A(net5914),
    .B(net5974));
 sg13g2_xnor2_1 _23158_ (.Y(_05884_),
    .A(_05880_),
    .B(_05882_));
 sg13g2_nor2b_1 _23159_ (.A(_05883_),
    .B_N(_05884_),
    .Y(_05885_));
 sg13g2_a21oi_1 _23160_ (.A1(_05881_),
    .A2(_05882_),
    .Y(_05886_),
    .B1(_05885_));
 sg13g2_a22oi_1 _23161_ (.Y(_05887_),
    .B1(_05871_),
    .B2(_05872_),
    .A2(net5974),
    .A1(net5871));
 sg13g2_nor3_1 _23162_ (.A(_05873_),
    .B(_05886_),
    .C(_05887_),
    .Y(_05888_));
 sg13g2_xnor2_1 _23163_ (.Y(_05889_),
    .A(_05878_),
    .B(_05879_));
 sg13g2_nor2_1 _23164_ (.A(_05694_),
    .B(_05702_),
    .Y(_05890_));
 sg13g2_nor2b_1 _23165_ (.A(_05889_),
    .B_N(_05890_),
    .Y(_05891_));
 sg13g2_xnor2_1 _23166_ (.Y(_05892_),
    .A(_05883_),
    .B(_05884_));
 sg13g2_nand2_1 _23167_ (.Y(_05893_),
    .A(_05891_),
    .B(_05892_));
 sg13g2_and2_1 _23168_ (.A(net5944),
    .B(net6007),
    .X(_05894_));
 sg13g2_o21ai_1 _23169_ (.B1(_05878_),
    .Y(_05895_),
    .A1(_05877_),
    .A2(_05894_));
 sg13g2_nand2_1 _23170_ (.Y(_05896_),
    .A(net5974),
    .B(_05727_));
 sg13g2_or2_1 _23171_ (.X(_05897_),
    .B(_05896_),
    .A(_05895_));
 sg13g2_xnor2_1 _23172_ (.Y(_05898_),
    .A(_05889_),
    .B(_05890_));
 sg13g2_nor2b_1 _23173_ (.A(_05897_),
    .B_N(_05898_),
    .Y(_05899_));
 sg13g2_or4_2 _23174_ (.A(_08618_),
    .B(net6008),
    .C(_05625_),
    .D(net6043),
    .X(_05900_));
 sg13g2_xor2_1 _23175_ (.B(_05896_),
    .A(_05895_),
    .X(_05901_));
 sg13g2_nor2b_1 _23176_ (.A(_05900_),
    .B_N(_05901_),
    .Y(_05902_));
 sg13g2_xnor2_1 _23177_ (.Y(_05903_),
    .A(_05897_),
    .B(_05898_));
 sg13g2_a21oi_1 _23178_ (.A1(_05902_),
    .A2(_05903_),
    .Y(_05904_),
    .B1(_05899_));
 sg13g2_xnor2_1 _23179_ (.Y(_05905_),
    .A(_05891_),
    .B(_05892_));
 sg13g2_o21ai_1 _23180_ (.B1(_05893_),
    .Y(_05906_),
    .A1(_05904_),
    .A2(_05905_));
 sg13g2_o21ai_1 _23181_ (.B1(_05886_),
    .Y(_05907_),
    .A1(_05873_),
    .A2(_05887_));
 sg13g2_nor2b_1 _23182_ (.A(_05888_),
    .B_N(_05907_),
    .Y(_05908_));
 sg13g2_a21oi_1 _23183_ (.A1(_05906_),
    .A2(_05907_),
    .Y(_05909_),
    .B1(_05888_));
 sg13g2_a21oi_1 _23184_ (.A1(_05857_),
    .A2(_05875_),
    .Y(_05910_),
    .B1(_05874_));
 sg13g2_a21o_1 _23185_ (.A2(_05875_),
    .A1(_05857_),
    .B1(_05874_),
    .X(_05911_));
 sg13g2_nand2_1 _23186_ (.Y(_05912_),
    .A(_05876_),
    .B(_05911_));
 sg13g2_o21ai_1 _23187_ (.B1(_05876_),
    .Y(_05913_),
    .A1(_05909_),
    .A2(_05910_));
 sg13g2_or2_1 _23188_ (.X(_05914_),
    .B(_05859_),
    .A(_05858_));
 sg13g2_nand2b_1 _23189_ (.Y(_05915_),
    .B(_05914_),
    .A_N(_05860_));
 sg13g2_a21oi_1 _23190_ (.A1(_05913_),
    .A2(_05914_),
    .Y(_05916_),
    .B1(_05860_));
 sg13g2_xnor2_1 _23191_ (.Y(_05917_),
    .A(_05835_),
    .B(_05836_));
 sg13g2_o21ai_1 _23192_ (.B1(_05837_),
    .Y(_05918_),
    .A1(_05916_),
    .A2(_05917_));
 sg13g2_xor2_1 _23193_ (.B(_05817_),
    .A(_05816_),
    .X(_05919_));
 sg13g2_a21oi_1 _23194_ (.A1(_05918_),
    .A2(_05919_),
    .Y(_05920_),
    .B1(_05818_));
 sg13g2_xor2_1 _23195_ (.B(_05795_),
    .A(_05775_),
    .X(_05921_));
 sg13g2_o21ai_1 _23196_ (.B1(_05796_),
    .Y(_05922_),
    .A1(_05920_),
    .A2(_05921_));
 sg13g2_xnor2_1 _23197_ (.Y(_05923_),
    .A(_05772_),
    .B(_05773_));
 sg13g2_a21oi_1 _23198_ (.A1(_05922_),
    .A2(_05923_),
    .Y(_05924_),
    .B1(_05774_));
 sg13g2_and2_1 _23199_ (.A(_05747_),
    .B(_05749_),
    .X(_05925_));
 sg13g2_xor2_1 _23200_ (.B(_05749_),
    .A(_05747_),
    .X(_05926_));
 sg13g2_o21ai_1 _23201_ (.B1(_05750_),
    .Y(_05927_),
    .A1(_05924_),
    .A2(_05925_));
 sg13g2_a21oi_1 _23202_ (.A1(_05724_),
    .A2(_05927_),
    .Y(_05928_),
    .B1(_05723_));
 sg13g2_o21ai_1 _23203_ (.B1(_05720_),
    .Y(_05929_),
    .A1(_05690_),
    .A2(_05721_));
 sg13g2_nor2_1 _23204_ (.A(_05660_),
    .B(_05718_),
    .Y(_05930_));
 sg13g2_xnor2_1 _23205_ (.Y(_05931_),
    .A(_05929_),
    .B(_05930_));
 sg13g2_xnor2_1 _23206_ (.Y(_05932_),
    .A(_05928_),
    .B(_05931_));
 sg13g2_nor2_1 _23207_ (.A(_08619_),
    .B(_05932_),
    .Y(_05933_));
 sg13g2_xor2_1 _23208_ (.B(_05927_),
    .A(_05725_),
    .X(_05934_));
 sg13g2_xnor2_1 _23209_ (.Y(_05935_),
    .A(_00110_),
    .B(_05934_));
 sg13g2_xnor2_1 _23210_ (.Y(_05936_),
    .A(_05924_),
    .B(_05926_));
 sg13g2_nor2_1 _23211_ (.A(_00109_),
    .B(_05936_),
    .Y(_05937_));
 sg13g2_xor2_1 _23212_ (.B(_05936_),
    .A(_00109_),
    .X(_05938_));
 sg13g2_xor2_1 _23213_ (.B(_05923_),
    .A(_05922_),
    .X(_05939_));
 sg13g2_nand2b_1 _23214_ (.Y(_05940_),
    .B(\atari2600.tia.audio_left_counter[12] ),
    .A_N(_05939_));
 sg13g2_xor2_1 _23215_ (.B(_05921_),
    .A(_05920_),
    .X(_05941_));
 sg13g2_a22oi_1 _23216_ (.Y(_05942_),
    .B1(_05941_),
    .B2(_00107_),
    .A2(_05939_),
    .A1(_00108_));
 sg13g2_o21ai_1 _23217_ (.B1(_05942_),
    .Y(_05943_),
    .A1(_00108_),
    .A2(_05939_));
 sg13g2_xor2_1 _23218_ (.B(_05917_),
    .A(_05916_),
    .X(_05944_));
 sg13g2_xor2_1 _23219_ (.B(_05919_),
    .A(_05918_),
    .X(_05945_));
 sg13g2_a22oi_1 _23220_ (.Y(_05946_),
    .B1(_05945_),
    .B2(_00106_),
    .A2(_05944_),
    .A1(_00105_));
 sg13g2_o21ai_1 _23221_ (.B1(_05946_),
    .Y(_05947_),
    .A1(_00106_),
    .A2(_05945_));
 sg13g2_xnor2_1 _23222_ (.Y(_05948_),
    .A(_05906_),
    .B(_05908_));
 sg13g2_xnor2_1 _23223_ (.Y(_05949_),
    .A(_00102_),
    .B(_05948_));
 sg13g2_xor2_1 _23224_ (.B(_05905_),
    .A(_05904_),
    .X(_05950_));
 sg13g2_or2_1 _23225_ (.X(_05951_),
    .B(_05950_),
    .A(_00100_));
 sg13g2_xnor2_1 _23226_ (.Y(_05952_),
    .A(_05902_),
    .B(_05903_));
 sg13g2_xnor2_1 _23227_ (.Y(_05953_),
    .A(_00099_),
    .B(_05952_));
 sg13g2_xnor2_1 _23228_ (.Y(_05954_),
    .A(_05900_),
    .B(_05901_));
 sg13g2_or2_1 _23229_ (.X(_05955_),
    .B(_05954_),
    .A(_00098_));
 sg13g2_and2_1 _23230_ (.A(_00098_),
    .B(_05954_),
    .X(_05956_));
 sg13g2_nand2_2 _23231_ (.Y(_05957_),
    .A(_00096_),
    .B(net5974));
 sg13g2_nor2_1 _23232_ (.A(\atari2600.tia.audio_left_counter[1] ),
    .B(_05957_),
    .Y(_05958_));
 sg13g2_a22oi_1 _23233_ (.Y(_05959_),
    .B1(net6007),
    .B2(net5974),
    .A2(net5944),
    .A1(_00096_));
 sg13g2_inv_1 _23234_ (.Y(_05960_),
    .A(_05959_));
 sg13g2_nand2_2 _23235_ (.Y(_05961_),
    .A(_05900_),
    .B(_05960_));
 sg13g2_xor2_1 _23236_ (.B(_05961_),
    .A(_00097_),
    .X(_05962_));
 sg13g2_nor2_1 _23237_ (.A(_05958_),
    .B(_05962_),
    .Y(_05963_));
 sg13g2_a21oi_1 _23238_ (.A1(\atari2600.tia.audio_left_counter[2] ),
    .A2(_05961_),
    .Y(_05964_),
    .B1(_05963_));
 sg13g2_o21ai_1 _23239_ (.B1(_05955_),
    .Y(_05965_),
    .A1(_05956_),
    .A2(_05964_));
 sg13g2_a22oi_1 _23240_ (.Y(_05966_),
    .B1(_05953_),
    .B2(_05965_),
    .A2(_05952_),
    .A1(\atari2600.tia.audio_left_counter[4] ));
 sg13g2_nand2_1 _23241_ (.Y(_05967_),
    .A(_05951_),
    .B(_05966_));
 sg13g2_nand2_1 _23242_ (.Y(_05968_),
    .A(_00100_),
    .B(_05950_));
 sg13g2_nand3_1 _23243_ (.B(_05967_),
    .C(_05968_),
    .A(_05949_),
    .Y(_05969_));
 sg13g2_xor2_1 _23244_ (.B(_05912_),
    .A(_05909_),
    .X(_05970_));
 sg13g2_nor2_1 _23245_ (.A(_00103_),
    .B(_05970_),
    .Y(_05971_));
 sg13g2_a21oi_1 _23246_ (.A1(\atari2600.tia.audio_left_counter[6] ),
    .A2(_05948_),
    .Y(_05972_),
    .B1(_05971_));
 sg13g2_xnor2_1 _23247_ (.Y(_05973_),
    .A(_05913_),
    .B(_05915_));
 sg13g2_nand2_1 _23248_ (.Y(_05974_),
    .A(_00103_),
    .B(_05970_));
 sg13g2_xnor2_1 _23249_ (.Y(_05975_),
    .A(_00104_),
    .B(_05973_));
 sg13g2_a221oi_1 _23250_ (.B2(_05969_),
    .C1(_05975_),
    .B1(_05972_),
    .A1(_00103_),
    .Y(_05976_),
    .A2(_05970_));
 sg13g2_nor2_1 _23251_ (.A(_00105_),
    .B(_05944_),
    .Y(_05977_));
 sg13g2_nor2b_1 _23252_ (.A(_05973_),
    .B_N(\atari2600.tia.audio_left_counter[8] ),
    .Y(_05978_));
 sg13g2_nor3_1 _23253_ (.A(_05976_),
    .B(_05977_),
    .C(_05978_),
    .Y(_05979_));
 sg13g2_nor2_1 _23254_ (.A(_05947_),
    .B(_05979_),
    .Y(_05980_));
 sg13g2_nor2_1 _23255_ (.A(_00107_),
    .B(_05941_),
    .Y(_05981_));
 sg13g2_nor2b_1 _23256_ (.A(_05945_),
    .B_N(\atari2600.tia.audio_left_counter[10] ),
    .Y(_05982_));
 sg13g2_nor3_1 _23257_ (.A(_05980_),
    .B(_05981_),
    .C(_05982_),
    .Y(_05983_));
 sg13g2_o21ai_1 _23258_ (.B1(_05940_),
    .Y(_05984_),
    .A1(_05943_),
    .A2(_05983_));
 sg13g2_nand3_1 _23259_ (.B(_05938_),
    .C(_05984_),
    .A(_05935_),
    .Y(_05985_));
 sg13g2_and2_1 _23260_ (.A(\atari2600.tia.audio_left_counter[14] ),
    .B(_05934_),
    .X(_05986_));
 sg13g2_a221oi_1 _23261_ (.B2(_05937_),
    .C1(_05986_),
    .B1(_05935_),
    .A1(_08619_),
    .Y(_05987_),
    .A2(_05932_));
 sg13g2_a21oi_2 _23262_ (.B1(_05933_),
    .Y(_05988_),
    .A2(_05987_),
    .A1(_05985_));
 sg13g2_nor2b_1 _23263_ (.A(net6263),
    .B_N(net6262),
    .Y(_05989_));
 sg13g2_nand2b_1 _23264_ (.Y(_05990_),
    .B(\atari2600.tia.audc0[3] ),
    .A_N(\atari2600.tia.audc0[2] ));
 sg13g2_a22oi_1 _23265_ (.Y(_05991_),
    .B1(_05989_),
    .B2(\atari2600.tia.audc0[1] ),
    .A2(_05662_),
    .A1(_08510_));
 sg13g2_nor2_2 _23266_ (.A(net6009),
    .B(_05991_),
    .Y(_05992_));
 sg13g2_nor3_1 _23267_ (.A(\atari2600.tia.audio_left_counter[0] ),
    .B(_05988_),
    .C(_05992_),
    .Y(_05993_));
 sg13g2_a21oi_1 _23268_ (.A1(net4537),
    .A2(_05992_),
    .Y(_05994_),
    .B1(_05993_));
 sg13g2_o21ai_1 _23269_ (.B1(_05614_),
    .Y(_00991_),
    .A1(_05366_),
    .A2(net4538));
 sg13g2_nand2_1 _23270_ (.Y(_05995_),
    .A(net7306),
    .B(net5838));
 sg13g2_nand2b_1 _23271_ (.Y(_05996_),
    .B(_05988_),
    .A_N(_05992_));
 sg13g2_nand2_1 _23272_ (.Y(_05997_),
    .A(\atari2600.tia.audio_left_counter[1] ),
    .B(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_or2_1 _23273_ (.X(_05998_),
    .B(\atari2600.tia.audio_left_counter[0] ),
    .A(net7306));
 sg13g2_nand4_1 _23274_ (.B(net4965),
    .C(_05997_),
    .A(net5803),
    .Y(_05999_),
    .D(_05998_));
 sg13g2_nand2_1 _23275_ (.Y(_00992_),
    .A(_05995_),
    .B(_05999_));
 sg13g2_nand2_1 _23276_ (.Y(_06000_),
    .A(net3398),
    .B(net5838));
 sg13g2_nor2_1 _23277_ (.A(_00097_),
    .B(_05997_),
    .Y(_06001_));
 sg13g2_xor2_1 _23278_ (.B(_05997_),
    .A(_00097_),
    .X(_06002_));
 sg13g2_nand3_1 _23279_ (.B(net4965),
    .C(_06002_),
    .A(net5803),
    .Y(_06003_));
 sg13g2_nand2_1 _23280_ (.Y(_00993_),
    .A(_06000_),
    .B(_06003_));
 sg13g2_nand2_1 _23281_ (.Y(_06004_),
    .A(net3019),
    .B(net5838));
 sg13g2_xnor2_1 _23282_ (.Y(_06005_),
    .A(_00098_),
    .B(_06001_));
 sg13g2_nand3_1 _23283_ (.B(net4965),
    .C(_06005_),
    .A(net5803),
    .Y(_06006_));
 sg13g2_nand2_1 _23284_ (.Y(_00994_),
    .A(_06004_),
    .B(_06006_));
 sg13g2_nand2_1 _23285_ (.Y(_06007_),
    .A(net3254),
    .B(net5838));
 sg13g2_nand4_1 _23286_ (.B(\atari2600.tia.audio_left_counter[2] ),
    .C(\atari2600.tia.audio_left_counter[1] ),
    .A(net3019),
    .Y(_06008_),
    .D(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_nor2_1 _23287_ (.A(_00099_),
    .B(_06008_),
    .Y(_06009_));
 sg13g2_xor2_1 _23288_ (.B(_06008_),
    .A(_00099_),
    .X(_06010_));
 sg13g2_nand3_1 _23289_ (.B(net4965),
    .C(_06010_),
    .A(net5807),
    .Y(_06011_));
 sg13g2_nand2_1 _23290_ (.Y(_00995_),
    .A(_06007_),
    .B(_06011_));
 sg13g2_nand2_1 _23291_ (.Y(_06012_),
    .A(net3106),
    .B(net5838));
 sg13g2_xnor2_1 _23292_ (.Y(_06013_),
    .A(_00100_),
    .B(_06009_));
 sg13g2_nand3_1 _23293_ (.B(net4965),
    .C(_06013_),
    .A(net5803),
    .Y(_06014_));
 sg13g2_nand2_1 _23294_ (.Y(_00996_),
    .A(_06012_),
    .B(_06014_));
 sg13g2_nand2_1 _23295_ (.Y(_06015_),
    .A(net3137),
    .B(net5839));
 sg13g2_nand2_1 _23296_ (.Y(_06016_),
    .A(\atari2600.tia.audio_left_counter[5] ),
    .B(\atari2600.tia.audio_left_counter[4] ));
 sg13g2_nor2_1 _23297_ (.A(_06008_),
    .B(_06016_),
    .Y(_06017_));
 sg13g2_nor3_1 _23298_ (.A(_00102_),
    .B(_06008_),
    .C(_06016_),
    .Y(_06018_));
 sg13g2_xnor2_1 _23299_ (.Y(_06019_),
    .A(_00102_),
    .B(_06017_));
 sg13g2_nand3_1 _23300_ (.B(net4966),
    .C(_06019_),
    .A(net5803),
    .Y(_06020_));
 sg13g2_nand2_1 _23301_ (.Y(_00997_),
    .A(_06015_),
    .B(_06020_));
 sg13g2_nand2_1 _23302_ (.Y(_06021_),
    .A(net3262),
    .B(net5838));
 sg13g2_xnor2_1 _23303_ (.Y(_06022_),
    .A(_00103_),
    .B(_06018_));
 sg13g2_nand3_1 _23304_ (.B(net4965),
    .C(_06022_),
    .A(net5803),
    .Y(_06023_));
 sg13g2_nand2_1 _23305_ (.Y(_00998_),
    .A(_06021_),
    .B(_06023_));
 sg13g2_nand2_1 _23306_ (.Y(_06024_),
    .A(net3828),
    .B(net5838));
 sg13g2_nand3_1 _23307_ (.B(net3137),
    .C(_06017_),
    .A(net3262),
    .Y(_06025_));
 sg13g2_inv_1 _23308_ (.Y(_06026_),
    .A(_06025_));
 sg13g2_nor2_1 _23309_ (.A(_00104_),
    .B(_06025_),
    .Y(_06027_));
 sg13g2_xor2_1 _23310_ (.B(_06025_),
    .A(_00104_),
    .X(_06028_));
 sg13g2_nand3_1 _23311_ (.B(net4965),
    .C(_06028_),
    .A(net5803),
    .Y(_06029_));
 sg13g2_nand2_1 _23312_ (.Y(_00999_),
    .A(_06024_),
    .B(_06029_));
 sg13g2_nand2_1 _23313_ (.Y(_06030_),
    .A(net3118),
    .B(net5839));
 sg13g2_xnor2_1 _23314_ (.Y(_06031_),
    .A(_00105_),
    .B(_06027_));
 sg13g2_nand3_1 _23315_ (.B(net4966),
    .C(_06031_),
    .A(net5804),
    .Y(_06032_));
 sg13g2_nand2_1 _23316_ (.Y(_01000_),
    .A(_06030_),
    .B(_06032_));
 sg13g2_nand2_1 _23317_ (.Y(_06033_),
    .A(net3777),
    .B(net5839));
 sg13g2_and3_1 _23318_ (.X(_06034_),
    .A(\atari2600.tia.audio_left_counter[9] ),
    .B(\atari2600.tia.audio_left_counter[8] ),
    .C(_06026_));
 sg13g2_nor2b_1 _23319_ (.A(_00106_),
    .B_N(_06034_),
    .Y(_06035_));
 sg13g2_xnor2_1 _23320_ (.Y(_06036_),
    .A(_00106_),
    .B(_06034_));
 sg13g2_nand3_1 _23321_ (.B(net4966),
    .C(_06036_),
    .A(net5804),
    .Y(_06037_));
 sg13g2_nand2_1 _23322_ (.Y(_01001_),
    .A(_06033_),
    .B(_06037_));
 sg13g2_nand2_1 _23323_ (.Y(_06038_),
    .A(net2986),
    .B(net5839));
 sg13g2_xnor2_1 _23324_ (.Y(_06039_),
    .A(_00107_),
    .B(_06035_));
 sg13g2_nand3_1 _23325_ (.B(net4966),
    .C(_06039_),
    .A(net5803),
    .Y(_06040_));
 sg13g2_nand2_1 _23326_ (.Y(_01002_),
    .A(_06038_),
    .B(_06040_));
 sg13g2_nand2_1 _23327_ (.Y(_06041_),
    .A(net3605),
    .B(net5839));
 sg13g2_nand3_1 _23328_ (.B(\atari2600.tia.audio_left_counter[10] ),
    .C(_06034_),
    .A(net2986),
    .Y(_06042_));
 sg13g2_inv_1 _23329_ (.Y(_06043_),
    .A(_06042_));
 sg13g2_nor2_1 _23330_ (.A(_00108_),
    .B(_06042_),
    .Y(_06044_));
 sg13g2_xor2_1 _23331_ (.B(_06042_),
    .A(_00108_),
    .X(_06045_));
 sg13g2_nand3_1 _23332_ (.B(net4965),
    .C(_06045_),
    .A(net5804),
    .Y(_06046_));
 sg13g2_nand2_1 _23333_ (.Y(_01003_),
    .A(_06041_),
    .B(_06046_));
 sg13g2_nand2_1 _23334_ (.Y(_06047_),
    .A(net3212),
    .B(net5839));
 sg13g2_xnor2_1 _23335_ (.Y(_06048_),
    .A(_00109_),
    .B(_06044_));
 sg13g2_nand3_1 _23336_ (.B(net4966),
    .C(_06048_),
    .A(net5804),
    .Y(_06049_));
 sg13g2_nand2_1 _23337_ (.Y(_01004_),
    .A(_06047_),
    .B(_06049_));
 sg13g2_nand2_1 _23338_ (.Y(_06050_),
    .A(net2965),
    .B(net5839));
 sg13g2_nand3_1 _23339_ (.B(\atari2600.tia.audio_left_counter[12] ),
    .C(_06043_),
    .A(\atari2600.tia.audio_left_counter[13] ),
    .Y(_06051_));
 sg13g2_nor2_1 _23340_ (.A(_00110_),
    .B(_06051_),
    .Y(_06052_));
 sg13g2_xor2_1 _23341_ (.B(_06051_),
    .A(_00110_),
    .X(_06053_));
 sg13g2_nand3_1 _23342_ (.B(net4966),
    .C(_06053_),
    .A(net5804),
    .Y(_06054_));
 sg13g2_nand2_1 _23343_ (.Y(_01005_),
    .A(_06050_),
    .B(_06054_));
 sg13g2_nand2_1 _23344_ (.Y(_06055_),
    .A(net2952),
    .B(net5839));
 sg13g2_xnor2_1 _23345_ (.Y(_06056_),
    .A(_00111_),
    .B(_06052_));
 sg13g2_nand3_1 _23346_ (.B(net4966),
    .C(_06056_),
    .A(net5804),
    .Y(_06057_));
 sg13g2_nand2_1 _23347_ (.Y(_01006_),
    .A(_06055_),
    .B(_06057_));
 sg13g2_nor2_2 _23348_ (.A(_08507_),
    .B(\atari2600.tia.audc1[0] ),
    .Y(_06058_));
 sg13g2_nand2_2 _23349_ (.Y(_06059_),
    .A(\atari2600.tia.audc1[1] ),
    .B(_08508_));
 sg13g2_nand2_1 _23350_ (.Y(_06060_),
    .A(\atari2600.tia.audc1[3] ),
    .B(_08506_));
 sg13g2_nand2_1 _23351_ (.Y(_06061_),
    .A(_08505_),
    .B(_08506_));
 sg13g2_nor2_2 _23352_ (.A(\atari2600.tia.audc1[1] ),
    .B(_06061_),
    .Y(_06062_));
 sg13g2_nor3_1 _23353_ (.A(_08507_),
    .B(_08508_),
    .C(_06060_),
    .Y(_06063_));
 sg13g2_a21oi_2 _23354_ (.B1(_06063_),
    .Y(_06064_),
    .A2(_06062_),
    .A1(_08508_));
 sg13g2_inv_1 _23355_ (.Y(_06065_),
    .A(_06064_));
 sg13g2_xnor2_1 _23356_ (.Y(_06066_),
    .A(\atari2600.tia.audf1[1] ),
    .B(\atari2600.tia.audf1[0] ));
 sg13g2_nor2_2 _23357_ (.A(_08501_),
    .B(_06066_),
    .Y(_06067_));
 sg13g2_mux2_1 _23358_ (.A0(\atari2600.tia.audf1[1] ),
    .A1(_06066_),
    .S(\atari2600.tia.audf1[2] ),
    .X(_06068_));
 sg13g2_xnor2_1 _23359_ (.Y(_06069_),
    .A(\atari2600.tia.audf1[3] ),
    .B(_06068_));
 sg13g2_inv_1 _23360_ (.Y(_06070_),
    .A(_06069_));
 sg13g2_nor2_2 _23361_ (.A(_08505_),
    .B(_08506_),
    .Y(_06071_));
 sg13g2_nand2_1 _23362_ (.Y(_06072_),
    .A(\atari2600.tia.audc1[3] ),
    .B(\atari2600.tia.audc1[2] ));
 sg13g2_nand3_1 _23363_ (.B(\atari2600.tia.audf1[1] ),
    .C(\atari2600.tia.audf1[0] ),
    .A(\atari2600.tia.audf1[2] ),
    .Y(_06073_));
 sg13g2_a21oi_1 _23364_ (.A1(\atari2600.tia.audf1[1] ),
    .A2(\atari2600.tia.audf1[0] ),
    .Y(_06074_),
    .B1(\atari2600.tia.audf1[2] ));
 sg13g2_nor2b_1 _23365_ (.A(_06074_),
    .B_N(_06073_),
    .Y(_06075_));
 sg13g2_nand2_1 _23366_ (.Y(_06076_),
    .A(\atari2600.tia.audf1[3] ),
    .B(_06075_));
 sg13g2_nand4_1 _23367_ (.B(\atari2600.tia.audf1[2] ),
    .C(\atari2600.tia.audf1[1] ),
    .A(\atari2600.tia.audf1[3] ),
    .Y(_06077_),
    .D(\atari2600.tia.audf1[0] ));
 sg13g2_nor2_1 _23368_ (.A(_00128_),
    .B(_06077_),
    .Y(_06078_));
 sg13g2_xor2_1 _23369_ (.B(_06077_),
    .A(_00128_),
    .X(_06079_));
 sg13g2_xnor2_1 _23370_ (.Y(_06080_),
    .A(_00128_),
    .B(_06077_));
 sg13g2_xnor2_1 _23371_ (.Y(_06081_),
    .A(\atari2600.tia.audf1[3] ),
    .B(_06073_));
 sg13g2_nand2_1 _23372_ (.Y(_06082_),
    .A(net6259),
    .B(_06081_));
 sg13g2_xnor2_1 _23373_ (.Y(_06083_),
    .A(net6259),
    .B(_06081_));
 sg13g2_nor2_1 _23374_ (.A(_06080_),
    .B(_06083_),
    .Y(_06084_));
 sg13g2_xnor2_1 _23375_ (.Y(_06085_),
    .A(_06080_),
    .B(_06083_));
 sg13g2_nor2_1 _23376_ (.A(_06076_),
    .B(_06085_),
    .Y(_06086_));
 sg13g2_xor2_1 _23377_ (.B(_06085_),
    .A(_06076_),
    .X(_06087_));
 sg13g2_nand2_1 _23378_ (.Y(_06088_),
    .A(_08501_),
    .B(\atari2600.tia.audf1[1] ));
 sg13g2_o21ai_1 _23379_ (.B1(\atari2600.tia.audf1[3] ),
    .Y(_06089_),
    .A1(\atari2600.tia.audf1[0] ),
    .A2(_06088_));
 sg13g2_o21ai_1 _23380_ (.B1(_06089_),
    .Y(_06090_),
    .A1(\atari2600.tia.audf1[3] ),
    .A2(_06067_));
 sg13g2_inv_1 _23381_ (.Y(_06091_),
    .A(_06090_));
 sg13g2_a21o_1 _23382_ (.A2(_06091_),
    .A1(_06087_),
    .B1(_06086_),
    .X(_06092_));
 sg13g2_nor2_1 _23383_ (.A(_06066_),
    .B(_06080_),
    .Y(_06093_));
 sg13g2_xnor2_1 _23384_ (.Y(_06094_),
    .A(_06066_),
    .B(_06079_));
 sg13g2_nor2b_1 _23385_ (.A(_06082_),
    .B_N(_06094_),
    .Y(_06095_));
 sg13g2_inv_1 _23386_ (.Y(_06096_),
    .A(_06095_));
 sg13g2_xnor2_1 _23387_ (.Y(_06097_),
    .A(_06082_),
    .B(_06094_));
 sg13g2_nor2_1 _23388_ (.A(_06078_),
    .B(_06097_),
    .Y(_06098_));
 sg13g2_nor2b_1 _23389_ (.A(_06098_),
    .B_N(_06084_),
    .Y(_06099_));
 sg13g2_xnor2_1 _23390_ (.Y(_06100_),
    .A(_06084_),
    .B(_06098_));
 sg13g2_xor2_1 _23391_ (.B(_06100_),
    .A(_06092_),
    .X(_06101_));
 sg13g2_xnor2_1 _23392_ (.Y(_06102_),
    .A(_06092_),
    .B(_06100_));
 sg13g2_nand2_1 _23393_ (.Y(_06103_),
    .A(net6006),
    .B(_06101_));
 sg13g2_nor2_2 _23394_ (.A(net6042),
    .B(_06103_),
    .Y(_06104_));
 sg13g2_nor2_2 _23395_ (.A(_06059_),
    .B(_06069_),
    .Y(_06105_));
 sg13g2_nand2_1 _23396_ (.Y(_06106_),
    .A(_06070_),
    .B(_06104_));
 sg13g2_xnor2_1 _23397_ (.Y(_06107_),
    .A(_06087_),
    .B(_06090_));
 sg13g2_xnor2_1 _23398_ (.Y(_06108_),
    .A(_06087_),
    .B(_06091_));
 sg13g2_a21o_1 _23399_ (.A2(_06100_),
    .A1(_06092_),
    .B1(_06099_),
    .X(_06109_));
 sg13g2_nor3_1 _23400_ (.A(_06075_),
    .B(_06078_),
    .C(_06093_),
    .Y(_06110_));
 sg13g2_a21o_1 _23401_ (.A2(_06079_),
    .A1(_06067_),
    .B1(_06110_),
    .X(_06111_));
 sg13g2_nor2_1 _23402_ (.A(_06096_),
    .B(_06111_),
    .Y(_06112_));
 sg13g2_xnor2_1 _23403_ (.Y(_06113_),
    .A(_06096_),
    .B(_06111_));
 sg13g2_inv_1 _23404_ (.Y(_06114_),
    .A(_06113_));
 sg13g2_nand2_1 _23405_ (.Y(_06115_),
    .A(_06109_),
    .B(_06114_));
 sg13g2_xnor2_1 _23406_ (.Y(_06116_),
    .A(_06109_),
    .B(_06113_));
 sg13g2_xnor2_1 _23407_ (.Y(_06117_),
    .A(_06109_),
    .B(_06114_));
 sg13g2_nor2_1 _23408_ (.A(_06059_),
    .B(_06117_),
    .Y(_06118_));
 sg13g2_nor3_1 _23409_ (.A(_06059_),
    .B(net6042),
    .C(_06117_),
    .Y(_06119_));
 sg13g2_nand2_2 _23410_ (.Y(_06120_),
    .A(net6006),
    .B(_06107_));
 sg13g2_nor2_1 _23411_ (.A(net6042),
    .B(_06120_),
    .Y(_06121_));
 sg13g2_and2_1 _23412_ (.A(_06116_),
    .B(_06121_),
    .X(_06122_));
 sg13g2_and2_1 _23413_ (.A(net6006),
    .B(_06061_),
    .X(_06123_));
 sg13g2_a21oi_1 _23414_ (.A1(_06116_),
    .A2(_06123_),
    .Y(_06124_),
    .B1(_06121_));
 sg13g2_or2_1 _23415_ (.X(_06125_),
    .B(_06124_),
    .A(_06122_));
 sg13g2_nor2_1 _23416_ (.A(_06106_),
    .B(_06125_),
    .Y(_06126_));
 sg13g2_a21oi_1 _23417_ (.A1(_06067_),
    .A2(_06079_),
    .Y(_06127_),
    .B1(_06081_));
 sg13g2_and3_1 _23418_ (.X(_06128_),
    .A(_06067_),
    .B(_06079_),
    .C(_06081_));
 sg13g2_nor2_1 _23419_ (.A(_06112_),
    .B(_06128_),
    .Y(_06129_));
 sg13g2_o21ai_1 _23420_ (.B1(_06129_),
    .Y(_06130_),
    .A1(_06115_),
    .A2(_06127_));
 sg13g2_a21o_2 _23421_ (.A2(_06130_),
    .A1(_06079_),
    .B1(_06078_),
    .X(_06131_));
 sg13g2_nand2_1 _23422_ (.Y(_06132_),
    .A(net6006),
    .B(net6042));
 sg13g2_nand2_1 _23423_ (.Y(_06133_),
    .A(_08505_),
    .B(\atari2600.tia.audc1[1] ));
 sg13g2_nand3_1 _23424_ (.B(_06059_),
    .C(_06133_),
    .A(\atari2600.tia.audc1[2] ),
    .Y(_06134_));
 sg13g2_and2_1 _23425_ (.A(_06132_),
    .B(net5971),
    .X(_06135_));
 sg13g2_nand2_1 _23426_ (.Y(_06136_),
    .A(_06132_),
    .B(net5972));
 sg13g2_xnor2_1 _23427_ (.Y(_06137_),
    .A(_06080_),
    .B(_06130_));
 sg13g2_nor2_1 _23428_ (.A(_06127_),
    .B(_06128_),
    .Y(_06138_));
 sg13g2_a21oi_1 _23429_ (.A1(_06109_),
    .A2(_06114_),
    .Y(_06139_),
    .B1(_06112_));
 sg13g2_xnor2_1 _23430_ (.Y(_06140_),
    .A(_06138_),
    .B(_06139_));
 sg13g2_and2_2 _23431_ (.A(_06058_),
    .B(_06140_),
    .X(_06141_));
 sg13g2_nand2_1 _23432_ (.Y(_06142_),
    .A(_06058_),
    .B(net5757));
 sg13g2_nand2_1 _23433_ (.Y(_06143_),
    .A(net5756),
    .B(_06141_));
 sg13g2_nor2_1 _23434_ (.A(net6006),
    .B(_06071_),
    .Y(_06144_));
 sg13g2_nand2_1 _23435_ (.Y(_06145_),
    .A(_06059_),
    .B(net6042));
 sg13g2_o21ai_1 _23436_ (.B1(_06145_),
    .Y(_06146_),
    .A1(net5756),
    .A2(_06141_));
 sg13g2_a21oi_1 _23437_ (.A1(net5756),
    .A2(_06141_),
    .Y(_06147_),
    .B1(_06146_));
 sg13g2_a21o_1 _23438_ (.A2(net5943),
    .A1(_06131_),
    .B1(_06147_),
    .X(_06148_));
 sg13g2_xor2_1 _23439_ (.B(_06125_),
    .A(_06106_),
    .X(_06149_));
 sg13g2_a21oi_2 _23440_ (.B1(_06126_),
    .Y(_06150_),
    .A2(_06149_),
    .A1(_06148_));
 sg13g2_and2_1 _23441_ (.A(_06104_),
    .B(_06140_),
    .X(_06151_));
 sg13g2_a21oi_1 _23442_ (.A1(net5973),
    .A2(_06140_),
    .Y(_06152_),
    .B1(_06104_));
 sg13g2_nor2_1 _23443_ (.A(_06151_),
    .B(_06152_),
    .Y(_06153_));
 sg13g2_and2_1 _23444_ (.A(_06122_),
    .B(_06153_),
    .X(_06154_));
 sg13g2_xor2_1 _23445_ (.B(_06153_),
    .A(_06122_),
    .X(_06155_));
 sg13g2_nand2_1 _23446_ (.Y(_06156_),
    .A(_06131_),
    .B(_06145_));
 sg13g2_nand2_1 _23447_ (.Y(_06157_),
    .A(_06142_),
    .B(_06156_));
 sg13g2_and2_1 _23448_ (.A(_06155_),
    .B(_06157_),
    .X(_06158_));
 sg13g2_xnor2_1 _23449_ (.Y(_06159_),
    .A(_06155_),
    .B(_06157_));
 sg13g2_nor2_1 _23450_ (.A(_06150_),
    .B(_06159_),
    .Y(_06160_));
 sg13g2_xor2_1 _23451_ (.B(_06159_),
    .A(_06150_),
    .X(_06161_));
 sg13g2_nor2b_1 _23452_ (.A(_06143_),
    .B_N(_06161_),
    .Y(_06162_));
 sg13g2_nor2_1 _23453_ (.A(_06160_),
    .B(_06162_),
    .Y(_06163_));
 sg13g2_nand2_1 _23454_ (.Y(_06164_),
    .A(_06058_),
    .B(_06131_));
 sg13g2_nor2_1 _23455_ (.A(_06072_),
    .B(_06142_),
    .Y(_06165_));
 sg13g2_nand2_1 _23456_ (.Y(_06166_),
    .A(_06119_),
    .B(net5756));
 sg13g2_a21oi_1 _23457_ (.A1(net5973),
    .A2(net5756),
    .Y(_06167_),
    .B1(_06119_));
 sg13g2_a21oi_1 _23458_ (.A1(_06119_),
    .A2(net5756),
    .Y(_06168_),
    .B1(_06167_));
 sg13g2_nand2_1 _23459_ (.Y(_06169_),
    .A(_06151_),
    .B(_06168_));
 sg13g2_xor2_1 _23460_ (.B(_06168_),
    .A(_06151_),
    .X(_06170_));
 sg13g2_nand2b_1 _23461_ (.Y(_06171_),
    .B(_06170_),
    .A_N(_06164_));
 sg13g2_xnor2_1 _23462_ (.Y(_06172_),
    .A(_06164_),
    .B(_06170_));
 sg13g2_nor3_1 _23463_ (.A(_06154_),
    .B(_06158_),
    .C(_06172_),
    .Y(_06173_));
 sg13g2_o21ai_1 _23464_ (.B1(_06172_),
    .Y(_06174_),
    .A1(_06154_),
    .A2(_06158_));
 sg13g2_nor2b_1 _23465_ (.A(_06173_),
    .B_N(_06174_),
    .Y(_06175_));
 sg13g2_o21ai_1 _23466_ (.B1(_06175_),
    .Y(_06176_),
    .A1(_06160_),
    .A2(_06162_));
 sg13g2_a22oi_1 _23467_ (.Y(_06177_),
    .B1(_06141_),
    .B2(_06071_),
    .A2(_06131_),
    .A1(net5973));
 sg13g2_nand2_1 _23468_ (.Y(_06178_),
    .A(_06166_),
    .B(_06177_));
 sg13g2_or2_1 _23469_ (.X(_06179_),
    .B(_06177_),
    .A(_06166_));
 sg13g2_nand4_1 _23470_ (.B(_06171_),
    .C(_06178_),
    .A(_06169_),
    .Y(_06180_),
    .D(_06179_));
 sg13g2_or2_1 _23471_ (.X(_06181_),
    .B(_06180_),
    .A(_06176_));
 sg13g2_xnor2_1 _23472_ (.Y(_06182_),
    .A(_06143_),
    .B(_06161_));
 sg13g2_xor2_1 _23473_ (.B(\atari2600.tia.audf1[0] ),
    .A(\atari2600.tia.audf1[2] ),
    .X(_06183_));
 sg13g2_nand2_1 _23474_ (.Y(_06184_),
    .A(net6006),
    .B(_06183_));
 sg13g2_nor2_1 _23475_ (.A(net6042),
    .B(_06184_),
    .Y(_06185_));
 sg13g2_nand2_1 _23476_ (.Y(_06186_),
    .A(_06107_),
    .B(_06185_));
 sg13g2_a22oi_1 _23477_ (.Y(_06187_),
    .B1(_06123_),
    .B2(_06101_),
    .A2(_06105_),
    .A1(_06071_));
 sg13g2_a21oi_1 _23478_ (.A1(_06070_),
    .A2(_06104_),
    .Y(_06188_),
    .B1(_06187_));
 sg13g2_inv_1 _23479_ (.Y(_06189_),
    .A(_06188_));
 sg13g2_xor2_1 _23480_ (.B(_06188_),
    .A(_06186_),
    .X(_06190_));
 sg13g2_xor2_1 _23481_ (.B(_06140_),
    .A(_06118_),
    .X(_06191_));
 sg13g2_and4_1 _23482_ (.A(net5943),
    .B(net5756),
    .C(_06145_),
    .D(_06191_),
    .X(_06192_));
 sg13g2_a22oi_1 _23483_ (.Y(_06193_),
    .B1(net5970),
    .B2(_06191_),
    .A2(net5756),
    .A1(net5943));
 sg13g2_or3_1 _23484_ (.A(_06190_),
    .B(_06192_),
    .C(_06193_),
    .X(_06194_));
 sg13g2_o21ai_1 _23485_ (.B1(_06194_),
    .Y(_06195_),
    .A1(_06186_),
    .A2(_06189_));
 sg13g2_xnor2_1 _23486_ (.Y(_06196_),
    .A(_06148_),
    .B(_06149_));
 sg13g2_nor2b_1 _23487_ (.A(_06196_),
    .B_N(_06195_),
    .Y(_06197_));
 sg13g2_a21o_1 _23488_ (.A2(_06141_),
    .A1(_06116_),
    .B1(_06192_),
    .X(_06198_));
 sg13g2_xnor2_1 _23489_ (.Y(_06199_),
    .A(_06195_),
    .B(_06196_));
 sg13g2_a21oi_2 _23490_ (.B1(_06197_),
    .Y(_06200_),
    .A2(_06199_),
    .A1(_06198_));
 sg13g2_nand2b_1 _23491_ (.Y(_06201_),
    .B(_06182_),
    .A_N(_06200_));
 sg13g2_xnor2_1 _23492_ (.Y(_06202_),
    .A(_06163_),
    .B(_06175_));
 sg13g2_nor2b_1 _23493_ (.A(_06201_),
    .B_N(_06202_),
    .Y(_06203_));
 sg13g2_xnor2_1 _23494_ (.Y(_06204_),
    .A(_06182_),
    .B(_06200_));
 sg13g2_xnor2_1 _23495_ (.Y(_06205_),
    .A(_06198_),
    .B(_06199_));
 sg13g2_xor2_1 _23496_ (.B(_06066_),
    .A(net6258),
    .X(_06206_));
 sg13g2_xnor2_1 _23497_ (.Y(_06207_),
    .A(net6259),
    .B(_06066_));
 sg13g2_nor2_1 _23498_ (.A(_06059_),
    .B(_06206_),
    .Y(_06208_));
 sg13g2_nor4_2 _23499_ (.A(_06059_),
    .B(_06069_),
    .C(net6042),
    .Y(_06209_),
    .D(_06206_));
 sg13g2_a21oi_1 _23500_ (.A1(_06107_),
    .A2(_06123_),
    .Y(_06210_),
    .B1(_06185_));
 sg13g2_a21oi_1 _23501_ (.A1(_06107_),
    .A2(_06185_),
    .Y(_06211_),
    .B1(_06210_));
 sg13g2_nand2_1 _23502_ (.Y(_06212_),
    .A(_06209_),
    .B(_06211_));
 sg13g2_xnor2_1 _23503_ (.Y(_06213_),
    .A(_06209_),
    .B(_06211_));
 sg13g2_nand2b_1 _23504_ (.Y(_06214_),
    .B(_06116_),
    .A_N(_06103_));
 sg13g2_a21oi_1 _23505_ (.A1(_06103_),
    .A2(_06117_),
    .Y(_06215_),
    .B1(_06144_));
 sg13g2_and4_1 _23506_ (.A(net5943),
    .B(_06140_),
    .C(_06214_),
    .D(_06215_),
    .X(_06216_));
 sg13g2_a22oi_1 _23507_ (.Y(_06217_),
    .B1(_06214_),
    .B2(_06215_),
    .A2(_06140_),
    .A1(net5943));
 sg13g2_or3_1 _23508_ (.A(_06213_),
    .B(_06216_),
    .C(_06217_),
    .X(_06218_));
 sg13g2_nand2_1 _23509_ (.Y(_06219_),
    .A(_06212_),
    .B(_06218_));
 sg13g2_o21ai_1 _23510_ (.B1(_06190_),
    .Y(_06220_),
    .A1(_06192_),
    .A2(_06193_));
 sg13g2_nand3_1 _23511_ (.B(_06219_),
    .C(_06220_),
    .A(_06194_),
    .Y(_06221_));
 sg13g2_a21o_1 _23512_ (.A2(_06118_),
    .A1(_06101_),
    .B1(_06216_),
    .X(_06222_));
 sg13g2_a21o_1 _23513_ (.A2(_06220_),
    .A1(_06194_),
    .B1(_06219_),
    .X(_06223_));
 sg13g2_nand3_1 _23514_ (.B(_06222_),
    .C(_06223_),
    .A(_06221_),
    .Y(_06224_));
 sg13g2_and2_1 _23515_ (.A(_06221_),
    .B(_06224_),
    .X(_06225_));
 sg13g2_or2_1 _23516_ (.X(_06226_),
    .B(_06225_),
    .A(_06205_));
 sg13g2_inv_1 _23517_ (.Y(_06227_),
    .A(_06226_));
 sg13g2_nand2_1 _23518_ (.Y(_06228_),
    .A(_06204_),
    .B(_06227_));
 sg13g2_xor2_1 _23519_ (.B(_06225_),
    .A(_06205_),
    .X(_06229_));
 sg13g2_nand3_1 _23520_ (.B(net6006),
    .C(_06071_),
    .A(net6258),
    .Y(_06230_));
 sg13g2_and2_1 _23521_ (.A(net6259),
    .B(_06185_),
    .X(_06231_));
 sg13g2_inv_1 _23522_ (.Y(_06232_),
    .A(_06231_));
 sg13g2_a22oi_1 _23523_ (.Y(_06233_),
    .B1(_06208_),
    .B2(_06071_),
    .A2(net5973),
    .A1(_06070_));
 sg13g2_or2_1 _23524_ (.X(_06234_),
    .B(_06233_),
    .A(_06209_));
 sg13g2_xnor2_1 _23525_ (.Y(_06235_),
    .A(_06232_),
    .B(_06234_));
 sg13g2_nor2_1 _23526_ (.A(_06102_),
    .B(_06120_),
    .Y(_06236_));
 sg13g2_or2_1 _23527_ (.X(_06237_),
    .B(_06120_),
    .A(_06102_));
 sg13g2_a21oi_1 _23528_ (.A1(_06102_),
    .A2(_06120_),
    .Y(_06238_),
    .B1(_06144_));
 sg13g2_and4_1 _23529_ (.A(_06116_),
    .B(net5942),
    .C(_06237_),
    .D(_06238_),
    .X(_06239_));
 sg13g2_a22oi_1 _23530_ (.Y(_06240_),
    .B1(_06237_),
    .B2(_06238_),
    .A2(net5943),
    .A1(_06116_));
 sg13g2_or3_1 _23531_ (.A(_06235_),
    .B(_06239_),
    .C(_06240_),
    .X(_06241_));
 sg13g2_o21ai_1 _23532_ (.B1(_06241_),
    .Y(_06242_),
    .A1(_06232_),
    .A2(_06234_));
 sg13g2_o21ai_1 _23533_ (.B1(_06213_),
    .Y(_06243_),
    .A1(_06216_),
    .A2(_06217_));
 sg13g2_nand3_1 _23534_ (.B(_06242_),
    .C(_06243_),
    .A(_06218_),
    .Y(_06244_));
 sg13g2_or2_1 _23535_ (.X(_06245_),
    .B(_06239_),
    .A(_06236_));
 sg13g2_a21o_1 _23536_ (.A2(_06243_),
    .A1(_06218_),
    .B1(_06242_),
    .X(_06246_));
 sg13g2_nand3_1 _23537_ (.B(_06245_),
    .C(_06246_),
    .A(_06244_),
    .Y(_06247_));
 sg13g2_nand2_1 _23538_ (.Y(_06248_),
    .A(_06244_),
    .B(_06247_));
 sg13g2_a21o_1 _23539_ (.A2(_06223_),
    .A1(_06221_),
    .B1(_06222_),
    .X(_06249_));
 sg13g2_nand3_1 _23540_ (.B(_06248_),
    .C(_06249_),
    .A(_06224_),
    .Y(_06250_));
 sg13g2_nand2_1 _23541_ (.Y(_06251_),
    .A(_06131_),
    .B(_06134_));
 sg13g2_inv_1 _23542_ (.Y(_06252_),
    .A(_06251_));
 sg13g2_a21o_1 _23543_ (.A2(_06249_),
    .A1(_06224_),
    .B1(_06248_),
    .X(_06253_));
 sg13g2_nand3_1 _23544_ (.B(_06252_),
    .C(_06253_),
    .A(_06250_),
    .Y(_06254_));
 sg13g2_nand2_1 _23545_ (.Y(_06255_),
    .A(_06250_),
    .B(_06254_));
 sg13g2_and2_1 _23546_ (.A(_06229_),
    .B(_06255_),
    .X(_06256_));
 sg13g2_nand2_1 _23547_ (.Y(_06257_),
    .A(net5973),
    .B(_06183_));
 sg13g2_a21oi_1 _23548_ (.A1(_06230_),
    .A2(_06257_),
    .Y(_06258_),
    .B1(_06231_));
 sg13g2_inv_1 _23549_ (.Y(_06259_),
    .A(_06258_));
 sg13g2_xnor2_1 _23550_ (.Y(_06260_),
    .A(_06105_),
    .B(_06108_));
 sg13g2_a22oi_1 _23551_ (.Y(_06261_),
    .B1(net5970),
    .B2(_06260_),
    .A2(net5942),
    .A1(_06101_));
 sg13g2_and4_1 _23552_ (.A(_06101_),
    .B(net5942),
    .C(net5970),
    .D(_06260_),
    .X(_06262_));
 sg13g2_nand4_1 _23553_ (.B(net5942),
    .C(net5970),
    .A(_06101_),
    .Y(_06263_),
    .D(_06260_));
 sg13g2_nand3b_1 _23554_ (.B(_06263_),
    .C(_06258_),
    .Y(_06264_),
    .A_N(_06261_));
 sg13g2_inv_1 _23555_ (.Y(_06265_),
    .A(_06264_));
 sg13g2_o21ai_1 _23556_ (.B1(_06235_),
    .Y(_06266_),
    .A1(_06239_),
    .A2(_06240_));
 sg13g2_nand3_1 _23557_ (.B(_06265_),
    .C(_06266_),
    .A(_06241_),
    .Y(_06267_));
 sg13g2_o21ai_1 _23558_ (.B1(_06263_),
    .Y(_06268_),
    .A1(_06069_),
    .A2(_06120_));
 sg13g2_a21o_1 _23559_ (.A2(_06266_),
    .A1(_06241_),
    .B1(_06265_),
    .X(_06269_));
 sg13g2_nand3_1 _23560_ (.B(_06268_),
    .C(_06269_),
    .A(_06267_),
    .Y(_06270_));
 sg13g2_nand2_1 _23561_ (.Y(_06271_),
    .A(_06267_),
    .B(_06270_));
 sg13g2_a21o_1 _23562_ (.A2(_06246_),
    .A1(_06244_),
    .B1(_06245_),
    .X(_06272_));
 sg13g2_nand3_1 _23563_ (.B(_06271_),
    .C(_06272_),
    .A(_06247_),
    .Y(_06273_));
 sg13g2_nand2_1 _23564_ (.Y(_06274_),
    .A(net5971),
    .B(net5757));
 sg13g2_a21oi_1 _23565_ (.A1(_06247_),
    .A2(_06272_),
    .Y(_06275_),
    .B1(_06271_));
 sg13g2_a21o_1 _23566_ (.A2(_06272_),
    .A1(_06247_),
    .B1(_06271_),
    .X(_06276_));
 sg13g2_and4_1 _23567_ (.A(net5971),
    .B(net5757),
    .C(_06273_),
    .D(_06276_),
    .X(_06277_));
 sg13g2_o21ai_1 _23568_ (.B1(_06273_),
    .Y(_06278_),
    .A1(_06274_),
    .A2(_06275_));
 sg13g2_a21o_1 _23569_ (.A2(_06253_),
    .A1(_06250_),
    .B1(_06252_),
    .X(_06279_));
 sg13g2_and3_1 _23570_ (.X(_06280_),
    .A(_06254_),
    .B(_06278_),
    .C(_06279_));
 sg13g2_nand3_1 _23571_ (.B(_06278_),
    .C(_06279_),
    .A(_06254_),
    .Y(_06281_));
 sg13g2_nand2_1 _23572_ (.Y(_06282_),
    .A(_06105_),
    .B(_06183_));
 sg13g2_o21ai_1 _23573_ (.B1(_06184_),
    .Y(_06283_),
    .A1(_06069_),
    .A2(_06144_));
 sg13g2_nand2_1 _23574_ (.Y(_06284_),
    .A(_06282_),
    .B(_06283_));
 sg13g2_o21ai_1 _23575_ (.B1(_06284_),
    .Y(_06285_),
    .A1(_06108_),
    .A2(_06135_));
 sg13g2_nand4_1 _23576_ (.B(net5942),
    .C(_06282_),
    .A(_06107_),
    .Y(_06286_),
    .D(_06283_));
 sg13g2_and4_1 _23577_ (.A(net5973),
    .B(_06207_),
    .C(_06285_),
    .D(_06286_),
    .X(_06287_));
 sg13g2_o21ai_1 _23578_ (.B1(_06259_),
    .Y(_06288_),
    .A1(_06261_),
    .A2(_06262_));
 sg13g2_nand3_1 _23579_ (.B(_06287_),
    .C(_06288_),
    .A(_06264_),
    .Y(_06289_));
 sg13g2_nand2_1 _23580_ (.Y(_06290_),
    .A(_06282_),
    .B(_06286_));
 sg13g2_a21o_1 _23581_ (.A2(_06288_),
    .A1(_06264_),
    .B1(_06287_),
    .X(_06291_));
 sg13g2_nand3_1 _23582_ (.B(_06290_),
    .C(_06291_),
    .A(_06289_),
    .Y(_06292_));
 sg13g2_nand2_1 _23583_ (.Y(_06293_),
    .A(_06289_),
    .B(_06292_));
 sg13g2_a21o_1 _23584_ (.A2(_06269_),
    .A1(_06267_),
    .B1(_06268_),
    .X(_06294_));
 sg13g2_nand3_1 _23585_ (.B(_06293_),
    .C(_06294_),
    .A(_06270_),
    .Y(_06295_));
 sg13g2_and2_1 _23586_ (.A(net5971),
    .B(_06140_),
    .X(_06296_));
 sg13g2_a21o_1 _23587_ (.A2(_06294_),
    .A1(_06270_),
    .B1(_06293_),
    .X(_06297_));
 sg13g2_nand3_1 _23588_ (.B(_06296_),
    .C(_06297_),
    .A(_06295_),
    .Y(_06298_));
 sg13g2_and2_1 _23589_ (.A(_06295_),
    .B(_06298_),
    .X(_06299_));
 sg13g2_a22oi_1 _23590_ (.Y(_06300_),
    .B1(_06273_),
    .B2(_06276_),
    .A2(net5757),
    .A1(net5971));
 sg13g2_nor3_1 _23591_ (.A(_06277_),
    .B(_06299_),
    .C(_06300_),
    .Y(_06301_));
 sg13g2_nand2_1 _23592_ (.Y(_06302_),
    .A(net6258),
    .B(net5973));
 sg13g2_nor2_1 _23593_ (.A(_06184_),
    .B(_06206_),
    .Y(_06303_));
 sg13g2_a21oi_1 _23594_ (.A1(net5970),
    .A2(_06183_),
    .Y(_06304_),
    .B1(_06208_));
 sg13g2_nor2_1 _23595_ (.A(_06303_),
    .B(_06304_),
    .Y(_06305_));
 sg13g2_nor2_1 _23596_ (.A(_06069_),
    .B(_06135_),
    .Y(_06306_));
 sg13g2_xor2_1 _23597_ (.B(_06306_),
    .A(_06305_),
    .X(_06307_));
 sg13g2_nand2b_1 _23598_ (.Y(_06308_),
    .B(_06307_),
    .A_N(_06302_));
 sg13g2_a22oi_1 _23599_ (.Y(_06309_),
    .B1(_06285_),
    .B2(_06286_),
    .A2(_06207_),
    .A1(net5973));
 sg13g2_or3_1 _23600_ (.A(_06287_),
    .B(_06308_),
    .C(_06309_),
    .X(_06310_));
 sg13g2_a21o_1 _23601_ (.A2(_06306_),
    .A1(_06305_),
    .B1(_06303_),
    .X(_06311_));
 sg13g2_o21ai_1 _23602_ (.B1(_06308_),
    .Y(_06312_),
    .A1(_06287_),
    .A2(_06309_));
 sg13g2_nand3_1 _23603_ (.B(_06311_),
    .C(_06312_),
    .A(_06310_),
    .Y(_06313_));
 sg13g2_nand2_1 _23604_ (.Y(_06314_),
    .A(_06310_),
    .B(_06313_));
 sg13g2_a21o_1 _23605_ (.A2(_06291_),
    .A1(_06289_),
    .B1(_06290_),
    .X(_06315_));
 sg13g2_and2_1 _23606_ (.A(_06292_),
    .B(_06315_),
    .X(_06316_));
 sg13g2_nand3_1 _23607_ (.B(_06314_),
    .C(_06315_),
    .A(_06292_),
    .Y(_06317_));
 sg13g2_a21o_1 _23608_ (.A2(_06315_),
    .A1(_06292_),
    .B1(_06314_),
    .X(_06318_));
 sg13g2_and4_1 _23609_ (.A(_06116_),
    .B(net5971),
    .C(_06317_),
    .D(_06318_),
    .X(_06319_));
 sg13g2_a21o_1 _23610_ (.A2(_06316_),
    .A1(_06314_),
    .B1(_06319_),
    .X(_06320_));
 sg13g2_a21o_1 _23611_ (.A2(_06297_),
    .A1(_06295_),
    .B1(_06296_),
    .X(_06321_));
 sg13g2_nand3_1 _23612_ (.B(_06320_),
    .C(_06321_),
    .A(_06298_),
    .Y(_06322_));
 sg13g2_xnor2_1 _23613_ (.Y(_06323_),
    .A(_06302_),
    .B(_06307_));
 sg13g2_nor2_1 _23614_ (.A(\atari2600.tia.audf1[0] ),
    .B(_06059_),
    .Y(_06324_));
 sg13g2_nand2_1 _23615_ (.Y(_06325_),
    .A(_06207_),
    .B(_06324_));
 sg13g2_a21oi_1 _23616_ (.A1(net5970),
    .A2(_06207_),
    .Y(_06326_),
    .B1(_06324_));
 sg13g2_a21oi_1 _23617_ (.A1(_06207_),
    .A2(_06324_),
    .Y(_06327_),
    .B1(_06326_));
 sg13g2_nand2_1 _23618_ (.Y(_06328_),
    .A(net5942),
    .B(_06183_));
 sg13g2_o21ai_1 _23619_ (.B1(_06325_),
    .Y(_06329_),
    .A1(_06326_),
    .A2(_06328_));
 sg13g2_nand2_1 _23620_ (.Y(_06330_),
    .A(_06323_),
    .B(_06329_));
 sg13g2_inv_1 _23621_ (.Y(_06331_),
    .A(_06330_));
 sg13g2_a21o_1 _23622_ (.A2(_06312_),
    .A1(_06310_),
    .B1(_06311_),
    .X(_06332_));
 sg13g2_nand3_1 _23623_ (.B(_06331_),
    .C(_06332_),
    .A(_06313_),
    .Y(_06333_));
 sg13g2_and2_1 _23624_ (.A(_06101_),
    .B(net5971),
    .X(_06334_));
 sg13g2_a21o_1 _23625_ (.A2(_06332_),
    .A1(_06313_),
    .B1(_06331_),
    .X(_06335_));
 sg13g2_nand3_1 _23626_ (.B(_06334_),
    .C(_06335_),
    .A(_06333_),
    .Y(_06336_));
 sg13g2_and2_1 _23627_ (.A(_06333_),
    .B(_06336_),
    .X(_06337_));
 sg13g2_a22oi_1 _23628_ (.Y(_06338_),
    .B1(_06317_),
    .B2(_06318_),
    .A2(net5971),
    .A1(_06116_));
 sg13g2_nor3_1 _23629_ (.A(_06319_),
    .B(_06337_),
    .C(_06338_),
    .Y(_06339_));
 sg13g2_nand2_1 _23630_ (.Y(_06340_),
    .A(net6258),
    .B(net5970));
 sg13g2_nand4_1 _23631_ (.B(net5942),
    .C(net5970),
    .A(net6258),
    .Y(_06341_),
    .D(_06207_));
 sg13g2_xor2_1 _23632_ (.B(_06328_),
    .A(_06327_),
    .X(_06342_));
 sg13g2_or2_1 _23633_ (.X(_06343_),
    .B(_06342_),
    .A(_06341_));
 sg13g2_inv_1 _23634_ (.Y(_06344_),
    .A(_06343_));
 sg13g2_xor2_1 _23635_ (.B(_06329_),
    .A(_06323_),
    .X(_06345_));
 sg13g2_nand2_1 _23636_ (.Y(_06346_),
    .A(_06107_),
    .B(net5972));
 sg13g2_xnor2_1 _23637_ (.Y(_06347_),
    .A(_06343_),
    .B(_06345_));
 sg13g2_nor2b_1 _23638_ (.A(_06346_),
    .B_N(_06347_),
    .Y(_06348_));
 sg13g2_a21oi_1 _23639_ (.A1(_06344_),
    .A2(_06345_),
    .Y(_06349_),
    .B1(_06348_));
 sg13g2_inv_1 _23640_ (.Y(_06350_),
    .A(_06349_));
 sg13g2_a21o_1 _23641_ (.A2(_06335_),
    .A1(_06333_),
    .B1(_06334_),
    .X(_06351_));
 sg13g2_nand2_1 _23642_ (.Y(_06352_),
    .A(_06336_),
    .B(_06351_));
 sg13g2_nand3_1 _23643_ (.B(_06350_),
    .C(_06351_),
    .A(_06336_),
    .Y(_06353_));
 sg13g2_xnor2_1 _23644_ (.Y(_06354_),
    .A(_06341_),
    .B(_06342_));
 sg13g2_nor2b_1 _23645_ (.A(_06069_),
    .B_N(net5972),
    .Y(_06355_));
 sg13g2_nor2b_1 _23646_ (.A(_06354_),
    .B_N(_06355_),
    .Y(_06356_));
 sg13g2_xnor2_1 _23647_ (.Y(_06357_),
    .A(_06346_),
    .B(_06347_));
 sg13g2_xnor2_1 _23648_ (.Y(_06358_),
    .A(_06354_),
    .B(_06355_));
 sg13g2_o21ai_1 _23649_ (.B1(_06340_),
    .Y(_06359_),
    .A1(_06135_),
    .A2(_06206_));
 sg13g2_and4_1 _23650_ (.A(net5972),
    .B(_06183_),
    .C(_06341_),
    .D(_06359_),
    .X(_06360_));
 sg13g2_nand4_1 _23651_ (.B(net6006),
    .C(_06066_),
    .A(net6258),
    .Y(_06361_),
    .D(net6042));
 sg13g2_a22oi_1 _23652_ (.Y(_06362_),
    .B1(_06341_),
    .B2(_06359_),
    .A2(_06183_),
    .A1(net5972));
 sg13g2_nor2_1 _23653_ (.A(_06360_),
    .B(_06362_),
    .Y(_06363_));
 sg13g2_nor3_1 _23654_ (.A(_06360_),
    .B(_06361_),
    .C(_06362_),
    .Y(_06364_));
 sg13g2_o21ai_1 _23655_ (.B1(_06358_),
    .Y(_06365_),
    .A1(_06360_),
    .A2(_06364_));
 sg13g2_xnor2_1 _23656_ (.Y(_06366_),
    .A(_06356_),
    .B(_06357_));
 sg13g2_nor2_1 _23657_ (.A(_06365_),
    .B(_06366_),
    .Y(_06367_));
 sg13g2_a21oi_1 _23658_ (.A1(_06356_),
    .A2(_06357_),
    .Y(_06368_),
    .B1(_06367_));
 sg13g2_a21o_1 _23659_ (.A2(_06357_),
    .A1(_06356_),
    .B1(_06367_),
    .X(_06369_));
 sg13g2_a21oi_1 _23660_ (.A1(_06336_),
    .A2(_06351_),
    .Y(_06370_),
    .B1(_06350_));
 sg13g2_xnor2_1 _23661_ (.Y(_06371_),
    .A(_06350_),
    .B(_06352_));
 sg13g2_o21ai_1 _23662_ (.B1(_06353_),
    .Y(_06372_),
    .A1(_06368_),
    .A2(_06370_));
 sg13g2_o21ai_1 _23663_ (.B1(_06337_),
    .Y(_06373_),
    .A1(_06319_),
    .A2(_06338_));
 sg13g2_nand2b_1 _23664_ (.Y(_06374_),
    .B(_06373_),
    .A_N(_06339_));
 sg13g2_a21oi_1 _23665_ (.A1(_06372_),
    .A2(_06373_),
    .Y(_06375_),
    .B1(_06339_));
 sg13g2_a21oi_1 _23666_ (.A1(_06298_),
    .A2(_06321_),
    .Y(_06376_),
    .B1(_06320_));
 sg13g2_a21o_1 _23667_ (.A2(_06321_),
    .A1(_06298_),
    .B1(_06320_),
    .X(_06377_));
 sg13g2_nand2_1 _23668_ (.Y(_06378_),
    .A(_06322_),
    .B(_06377_));
 sg13g2_o21ai_1 _23669_ (.B1(_06322_),
    .Y(_06379_),
    .A1(_06375_),
    .A2(_06376_));
 sg13g2_o21ai_1 _23670_ (.B1(_06299_),
    .Y(_06380_),
    .A1(_06277_),
    .A2(_06300_));
 sg13g2_nor2b_1 _23671_ (.A(_06301_),
    .B_N(_06380_),
    .Y(_06381_));
 sg13g2_a21oi_2 _23672_ (.B1(_06301_),
    .Y(_06382_),
    .A2(_06380_),
    .A1(_06379_));
 sg13g2_a21oi_1 _23673_ (.A1(_06254_),
    .A2(_06279_),
    .Y(_06383_),
    .B1(_06278_));
 sg13g2_nor3_1 _23674_ (.A(_06280_),
    .B(_06382_),
    .C(_06383_),
    .Y(_06384_));
 sg13g2_o21ai_1 _23675_ (.B1(_06281_),
    .Y(_06385_),
    .A1(_06382_),
    .A2(_06383_));
 sg13g2_xor2_1 _23676_ (.B(_06255_),
    .A(_06229_),
    .X(_06386_));
 sg13g2_a21oi_1 _23677_ (.A1(_06385_),
    .A2(_06386_),
    .Y(_06387_),
    .B1(_06256_));
 sg13g2_nor2_1 _23678_ (.A(_06204_),
    .B(_06227_),
    .Y(_06388_));
 sg13g2_xnor2_1 _23679_ (.Y(_06389_),
    .A(_06204_),
    .B(_06226_));
 sg13g2_o21ai_1 _23680_ (.B1(_06228_),
    .Y(_06390_),
    .A1(_06387_),
    .A2(_06388_));
 sg13g2_xnor2_1 _23681_ (.Y(_06391_),
    .A(_06201_),
    .B(_06202_));
 sg13g2_a21oi_1 _23682_ (.A1(_06390_),
    .A2(_06391_),
    .Y(_06392_),
    .B1(_06203_));
 sg13g2_nand2_1 _23683_ (.Y(_06393_),
    .A(_06174_),
    .B(_06176_));
 sg13g2_xor2_1 _23684_ (.B(_06393_),
    .A(_06180_),
    .X(_06394_));
 sg13g2_o21ai_1 _23685_ (.B1(_06181_),
    .Y(_06395_),
    .A1(_06392_),
    .A2(_06394_));
 sg13g2_a21o_1 _23686_ (.A2(_06177_),
    .A1(_06166_),
    .B1(_06174_),
    .X(_06396_));
 sg13g2_nand4_1 _23687_ (.B(_06171_),
    .C(_06179_),
    .A(_06169_),
    .Y(_06397_),
    .D(_06396_));
 sg13g2_xnor2_1 _23688_ (.Y(_06398_),
    .A(_06165_),
    .B(_06397_));
 sg13g2_xnor2_1 _23689_ (.Y(_06399_),
    .A(_06395_),
    .B(_06398_));
 sg13g2_nand2_1 _23690_ (.Y(_06400_),
    .A(_00126_),
    .B(_06399_));
 sg13g2_xor2_1 _23691_ (.B(_06394_),
    .A(_06392_),
    .X(_06401_));
 sg13g2_xnor2_1 _23692_ (.Y(_06402_),
    .A(_00125_),
    .B(_06401_));
 sg13g2_xor2_1 _23693_ (.B(_06391_),
    .A(_06390_),
    .X(_06403_));
 sg13g2_nand2_1 _23694_ (.Y(_06404_),
    .A(_00124_),
    .B(_06403_));
 sg13g2_xnor2_1 _23695_ (.Y(_06405_),
    .A(_06387_),
    .B(_06389_));
 sg13g2_xnor2_1 _23696_ (.Y(_06406_),
    .A(_00123_),
    .B(_06405_));
 sg13g2_xor2_1 _23697_ (.B(_06386_),
    .A(_06385_),
    .X(_06407_));
 sg13g2_nor2_1 _23698_ (.A(_00122_),
    .B(_06407_),
    .Y(_06408_));
 sg13g2_xnor2_1 _23699_ (.Y(_06409_),
    .A(_06379_),
    .B(_06381_));
 sg13g2_nand2_1 _23700_ (.Y(_06410_),
    .A(_08623_),
    .B(_06409_));
 sg13g2_nor2_1 _23701_ (.A(_08623_),
    .B(_06409_),
    .Y(_06411_));
 sg13g2_xnor2_1 _23702_ (.Y(_06412_),
    .A(_06375_),
    .B(_06378_));
 sg13g2_xnor2_1 _23703_ (.Y(_06413_),
    .A(_00119_),
    .B(_06412_));
 sg13g2_xor2_1 _23704_ (.B(_06374_),
    .A(_06372_),
    .X(_06414_));
 sg13g2_xnor2_1 _23705_ (.Y(_06415_),
    .A(_06369_),
    .B(_06371_));
 sg13g2_nor3_1 _23706_ (.A(_06358_),
    .B(_06360_),
    .C(_06364_),
    .Y(_06416_));
 sg13g2_nand2b_1 _23707_ (.Y(_06417_),
    .B(_06365_),
    .A_N(_06416_));
 sg13g2_a22oi_1 _23708_ (.Y(_06418_),
    .B1(_06207_),
    .B2(net5972),
    .A2(net5942),
    .A1(net6258));
 sg13g2_inv_1 _23709_ (.Y(_06419_),
    .A(_06418_));
 sg13g2_nand2_1 _23710_ (.Y(_06420_),
    .A(_06361_),
    .B(_06419_));
 sg13g2_nand3b_1 _23711_ (.B(net6258),
    .C(net5972),
    .Y(_06421_),
    .A_N(\atari2600.tia.audio_right_counter[1] ));
 sg13g2_xnor2_1 _23712_ (.Y(_06422_),
    .A(_00113_),
    .B(_06420_));
 sg13g2_a22oi_1 _23713_ (.Y(_06423_),
    .B1(_06421_),
    .B2(_06422_),
    .A2(_06420_),
    .A1(\atari2600.tia.audio_right_counter[2] ));
 sg13g2_nor2_1 _23714_ (.A(_00114_),
    .B(_06423_),
    .Y(_06424_));
 sg13g2_xnor2_1 _23715_ (.Y(_06425_),
    .A(_06361_),
    .B(_06363_));
 sg13g2_a21oi_1 _23716_ (.A1(_00114_),
    .A2(_06423_),
    .Y(_06426_),
    .B1(_06425_));
 sg13g2_or2_1 _23717_ (.X(_06427_),
    .B(_06426_),
    .A(_06424_));
 sg13g2_xor2_1 _23718_ (.B(_06366_),
    .A(_06365_),
    .X(_06428_));
 sg13g2_xnor2_1 _23719_ (.Y(_06429_),
    .A(_00115_),
    .B(_06417_));
 sg13g2_nor2_1 _23720_ (.A(_00116_),
    .B(_06428_),
    .Y(_06430_));
 sg13g2_a221oi_1 _23721_ (.B2(_06429_),
    .C1(_06430_),
    .B1(_06427_),
    .A1(\atari2600.tia.audio_right_counter[4] ),
    .Y(_06431_),
    .A2(_06417_));
 sg13g2_a21oi_1 _23722_ (.A1(_00116_),
    .A2(_06428_),
    .Y(_06432_),
    .B1(_06431_));
 sg13g2_xnor2_1 _23723_ (.Y(_06433_),
    .A(_00117_),
    .B(_06415_));
 sg13g2_a22oi_1 _23724_ (.Y(_06434_),
    .B1(_06432_),
    .B2(_06433_),
    .A2(_06415_),
    .A1(\atari2600.tia.audio_right_counter[6] ));
 sg13g2_nand2_1 _23725_ (.Y(_06435_),
    .A(_08622_),
    .B(_06414_));
 sg13g2_nor2_1 _23726_ (.A(_08622_),
    .B(_06414_),
    .Y(_06436_));
 sg13g2_a21oi_1 _23727_ (.A1(_06434_),
    .A2(_06435_),
    .Y(_06437_),
    .B1(_06436_));
 sg13g2_a22oi_1 _23728_ (.Y(_06438_),
    .B1(_06413_),
    .B2(_06437_),
    .A2(_06412_),
    .A1(\atari2600.tia.audio_right_counter[8] ));
 sg13g2_o21ai_1 _23729_ (.B1(_06410_),
    .Y(_06439_),
    .A1(_06411_),
    .A2(_06438_));
 sg13g2_o21ai_1 _23730_ (.B1(_06382_),
    .Y(_06440_),
    .A1(_06280_),
    .A2(_06383_));
 sg13g2_nand2b_1 _23731_ (.Y(_06441_),
    .B(_06440_),
    .A_N(_06384_));
 sg13g2_xnor2_1 _23732_ (.Y(_06442_),
    .A(_00121_),
    .B(_06441_));
 sg13g2_nand2_1 _23733_ (.Y(_06443_),
    .A(_06439_),
    .B(_06442_));
 sg13g2_a21oi_1 _23734_ (.A1(\atari2600.tia.audio_right_counter[10] ),
    .A2(_06441_),
    .Y(_06444_),
    .B1(_06408_));
 sg13g2_a221oi_1 _23735_ (.B2(_06444_),
    .C1(_06406_),
    .B1(_06443_),
    .A1(_00122_),
    .Y(_06445_),
    .A2(_06407_));
 sg13g2_nand2b_1 _23736_ (.Y(_06446_),
    .B(\atari2600.tia.audio_right_counter[12] ),
    .A_N(_06405_));
 sg13g2_o21ai_1 _23737_ (.B1(_06446_),
    .Y(_06447_),
    .A1(_00124_),
    .A2(_06403_));
 sg13g2_o21ai_1 _23738_ (.B1(_06404_),
    .Y(_06448_),
    .A1(_06445_),
    .A2(_06447_));
 sg13g2_nor2_1 _23739_ (.A(_00126_),
    .B(_06399_),
    .Y(_06449_));
 sg13g2_nand2b_1 _23740_ (.Y(_06450_),
    .B(\atari2600.tia.audio_right_counter[14] ),
    .A_N(_06401_));
 sg13g2_o21ai_1 _23741_ (.B1(_06450_),
    .Y(_06451_),
    .A1(_06402_),
    .A2(_06448_));
 sg13g2_a21oi_2 _23742_ (.B1(_06449_),
    .Y(_06452_),
    .A2(_06451_),
    .A1(_06400_));
 sg13g2_nand3b_1 _23743_ (.B(_06064_),
    .C(_06452_),
    .Y(_06453_),
    .A_N(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_nand2_1 _23744_ (.Y(_06454_),
    .A(net7351),
    .B(_06065_));
 sg13g2_a21oi_1 _23745_ (.A1(_06453_),
    .A2(_06454_),
    .Y(_06455_),
    .B1(_05366_));
 sg13g2_a21o_1 _23746_ (.A2(net5841),
    .A1(\atari2600.tia.audio_right_counter[0] ),
    .B1(_06455_),
    .X(_01007_));
 sg13g2_nand2_1 _23747_ (.Y(_06456_),
    .A(net7309),
    .B(net5841));
 sg13g2_nand2b_1 _23748_ (.Y(_06457_),
    .B(_06064_),
    .A_N(_06452_));
 sg13g2_nand2_1 _23749_ (.Y(_06458_),
    .A(\atari2600.tia.audio_right_counter[1] ),
    .B(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_or2_1 _23750_ (.X(_06459_),
    .B(\atari2600.tia.audio_right_counter[0] ),
    .A(net7309));
 sg13g2_nand4_1 _23751_ (.B(net4963),
    .C(_06458_),
    .A(net5805),
    .Y(_06460_),
    .D(_06459_));
 sg13g2_nand2_1 _23752_ (.Y(_01008_),
    .A(_06456_),
    .B(_06460_));
 sg13g2_nand2_1 _23753_ (.Y(_06461_),
    .A(net4210),
    .B(net5841));
 sg13g2_nor2_1 _23754_ (.A(_00113_),
    .B(_06458_),
    .Y(_06462_));
 sg13g2_xor2_1 _23755_ (.B(_06458_),
    .A(_00113_),
    .X(_06463_));
 sg13g2_nand3_1 _23756_ (.B(net4963),
    .C(_06463_),
    .A(net5806),
    .Y(_06464_));
 sg13g2_nand2_1 _23757_ (.Y(_01009_),
    .A(_06461_),
    .B(_06464_));
 sg13g2_nand2_1 _23758_ (.Y(_06465_),
    .A(net3091),
    .B(net5843));
 sg13g2_xnor2_1 _23759_ (.Y(_06466_),
    .A(_00114_),
    .B(_06462_));
 sg13g2_nand3_1 _23760_ (.B(net4963),
    .C(_06466_),
    .A(net5806),
    .Y(_06467_));
 sg13g2_nand2_1 _23761_ (.Y(_01010_),
    .A(_06465_),
    .B(_06467_));
 sg13g2_nand2_1 _23762_ (.Y(_06468_),
    .A(net3363),
    .B(net5843));
 sg13g2_nand4_1 _23763_ (.B(\atari2600.tia.audio_right_counter[2] ),
    .C(\atari2600.tia.audio_right_counter[1] ),
    .A(net3091),
    .Y(_06469_),
    .D(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_nor2_1 _23764_ (.A(_00115_),
    .B(_06469_),
    .Y(_06470_));
 sg13g2_xnor2_1 _23765_ (.Y(_06471_),
    .A(_08620_),
    .B(_06469_));
 sg13g2_nand3_1 _23766_ (.B(net4963),
    .C(_06471_),
    .A(net5806),
    .Y(_06472_));
 sg13g2_nand2_1 _23767_ (.Y(_01011_),
    .A(_06468_),
    .B(_06472_));
 sg13g2_nand2_1 _23768_ (.Y(_06473_),
    .A(net3027),
    .B(net5843));
 sg13g2_xnor2_1 _23769_ (.Y(_06474_),
    .A(_00116_),
    .B(_06470_));
 sg13g2_nand3_1 _23770_ (.B(net4963),
    .C(_06474_),
    .A(net5806),
    .Y(_06475_));
 sg13g2_nand2_1 _23771_ (.Y(_01012_),
    .A(_06473_),
    .B(_06475_));
 sg13g2_nand2_1 _23772_ (.Y(_06476_),
    .A(net3799),
    .B(net5841));
 sg13g2_nand2_1 _23773_ (.Y(_06477_),
    .A(\atari2600.tia.audio_right_counter[5] ),
    .B(\atari2600.tia.audio_right_counter[4] ));
 sg13g2_nor2_1 _23774_ (.A(_06469_),
    .B(_06477_),
    .Y(_06478_));
 sg13g2_nor3_1 _23775_ (.A(_00117_),
    .B(_06469_),
    .C(_06477_),
    .Y(_06479_));
 sg13g2_xnor2_1 _23776_ (.Y(_06480_),
    .A(_00117_),
    .B(_06478_));
 sg13g2_nand3_1 _23777_ (.B(net4963),
    .C(_06480_),
    .A(net5805),
    .Y(_06481_));
 sg13g2_nand2_1 _23778_ (.Y(_01013_),
    .A(_06476_),
    .B(_06481_));
 sg13g2_nand2_1 _23779_ (.Y(_06482_),
    .A(net2957),
    .B(net5840));
 sg13g2_xnor2_1 _23780_ (.Y(_06483_),
    .A(_00118_),
    .B(_06479_));
 sg13g2_nand3_1 _23781_ (.B(net4963),
    .C(_06483_),
    .A(net5805),
    .Y(_06484_));
 sg13g2_nand2_1 _23782_ (.Y(_01014_),
    .A(_06482_),
    .B(_06484_));
 sg13g2_nand2_1 _23783_ (.Y(_06485_),
    .A(net3043),
    .B(net5841));
 sg13g2_and2_1 _23784_ (.A(\atari2600.tia.audio_right_counter[7] ),
    .B(\atari2600.tia.audio_right_counter[6] ),
    .X(_06486_));
 sg13g2_nand2_1 _23785_ (.Y(_06487_),
    .A(_06478_),
    .B(_06486_));
 sg13g2_nor2_1 _23786_ (.A(_00119_),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_xor2_1 _23787_ (.B(_06487_),
    .A(_00119_),
    .X(_06489_));
 sg13g2_nand3_1 _23788_ (.B(net4964),
    .C(_06489_),
    .A(net5805),
    .Y(_06490_));
 sg13g2_nand2_1 _23789_ (.Y(_01015_),
    .A(_06485_),
    .B(_06490_));
 sg13g2_nand2_1 _23790_ (.Y(_06491_),
    .A(net2996),
    .B(net5840));
 sg13g2_xnor2_1 _23791_ (.Y(_06492_),
    .A(_00120_),
    .B(_06488_));
 sg13g2_nand3_1 _23792_ (.B(net4964),
    .C(_06492_),
    .A(net5805),
    .Y(_06493_));
 sg13g2_nand2_1 _23793_ (.Y(_01016_),
    .A(_06491_),
    .B(_06493_));
 sg13g2_nand2_1 _23794_ (.Y(_06494_),
    .A(net3843),
    .B(net5842));
 sg13g2_nand4_1 _23795_ (.B(net3043),
    .C(_06478_),
    .A(net2996),
    .Y(_06495_),
    .D(_06486_));
 sg13g2_inv_1 _23796_ (.Y(_06496_),
    .A(_06495_));
 sg13g2_nor2_1 _23797_ (.A(_00121_),
    .B(_06495_),
    .Y(_06497_));
 sg13g2_xor2_1 _23798_ (.B(_06495_),
    .A(_00121_),
    .X(_06498_));
 sg13g2_nand3_1 _23799_ (.B(net4964),
    .C(_06498_),
    .A(net5806),
    .Y(_06499_));
 sg13g2_nand2_1 _23800_ (.Y(_01017_),
    .A(_06494_),
    .B(_06499_));
 sg13g2_nand2_1 _23801_ (.Y(_06500_),
    .A(net3002),
    .B(net5842));
 sg13g2_xnor2_1 _23802_ (.Y(_06501_),
    .A(_00122_),
    .B(_06497_));
 sg13g2_nand3_1 _23803_ (.B(net4964),
    .C(_06501_),
    .A(net5805),
    .Y(_06502_));
 sg13g2_nand2_1 _23804_ (.Y(_01018_),
    .A(_06500_),
    .B(_06502_));
 sg13g2_nand2_1 _23805_ (.Y(_06503_),
    .A(net3175),
    .B(net5841));
 sg13g2_nand3_1 _23806_ (.B(\atari2600.tia.audio_right_counter[10] ),
    .C(_06496_),
    .A(net3002),
    .Y(_06504_));
 sg13g2_inv_1 _23807_ (.Y(_06505_),
    .A(_06504_));
 sg13g2_nor2_1 _23808_ (.A(_00123_),
    .B(_06504_),
    .Y(_06506_));
 sg13g2_xor2_1 _23809_ (.B(_06504_),
    .A(_00123_),
    .X(_06507_));
 sg13g2_nand3_1 _23810_ (.B(net4964),
    .C(_06507_),
    .A(net5805),
    .Y(_06508_));
 sg13g2_nand2_1 _23811_ (.Y(_01019_),
    .A(_06503_),
    .B(_06508_));
 sg13g2_nand2_1 _23812_ (.Y(_06509_),
    .A(net2974),
    .B(net5841));
 sg13g2_xnor2_1 _23813_ (.Y(_06510_),
    .A(_00124_),
    .B(_06506_));
 sg13g2_nand3_1 _23814_ (.B(net4964),
    .C(_06510_),
    .A(net5806),
    .Y(_06511_));
 sg13g2_nand2_1 _23815_ (.Y(_01020_),
    .A(_06509_),
    .B(_06511_));
 sg13g2_nand2_1 _23816_ (.Y(_06512_),
    .A(net3011),
    .B(net5841));
 sg13g2_nand3_1 _23817_ (.B(\atari2600.tia.audio_right_counter[12] ),
    .C(_06505_),
    .A(net2974),
    .Y(_06513_));
 sg13g2_nor2_1 _23818_ (.A(_00125_),
    .B(_06513_),
    .Y(_06514_));
 sg13g2_xnor2_1 _23819_ (.Y(_06515_),
    .A(_08624_),
    .B(_06513_));
 sg13g2_nand3_1 _23820_ (.B(net4964),
    .C(_06515_),
    .A(net5805),
    .Y(_06516_));
 sg13g2_nand2_1 _23821_ (.Y(_01021_),
    .A(_06512_),
    .B(_06516_));
 sg13g2_nand2_1 _23822_ (.Y(_06517_),
    .A(net2943),
    .B(net5842));
 sg13g2_xnor2_1 _23823_ (.Y(_06518_),
    .A(_00126_),
    .B(_06514_));
 sg13g2_nand3_1 _23824_ (.B(net4963),
    .C(_06518_),
    .A(net5806),
    .Y(_06519_));
 sg13g2_nand2_1 _23825_ (.Y(_01022_),
    .A(_06517_),
    .B(_06519_));
 sg13g2_o21ai_1 _23826_ (.B1(net5913),
    .Y(_06520_),
    .A1(_05988_),
    .A2(_05992_));
 sg13g2_nor4_1 _23827_ (.A(net6262),
    .B(net6263),
    .C(\atari2600.tia.audc0[1] ),
    .D(_08510_),
    .Y(_06521_));
 sg13g2_a21oi_1 _23828_ (.A1(\atari2600.tia.p4_l ),
    .A2(_06521_),
    .Y(_06522_),
    .B1(_05992_));
 sg13g2_nor2_1 _23829_ (.A(\atari2600.tia.audc0[1] ),
    .B(_05990_),
    .Y(_06523_));
 sg13g2_nor3_1 _23830_ (.A(net6262),
    .B(_08509_),
    .C(_08510_),
    .Y(_06524_));
 sg13g2_a22oi_1 _23831_ (.Y(_06525_),
    .B1(_06524_),
    .B2(net6263),
    .A2(_06523_),
    .A1(\atari2600.tia.audc0[0] ));
 sg13g2_nor3_1 _23832_ (.A(\atari2600.tia.audc0[1] ),
    .B(\atari2600.tia.audc0[0] ),
    .C(_05990_),
    .Y(_06526_));
 sg13g2_a221oi_1 _23833_ (.B2(net6263),
    .C1(_00155_),
    .B1(_06524_),
    .A1(_08509_),
    .Y(_06527_),
    .A2(_05989_));
 sg13g2_a21oi_1 _23834_ (.A1(_08497_),
    .A2(_06526_),
    .Y(_06528_),
    .B1(_06521_));
 sg13g2_o21ai_1 _23835_ (.B1(_06528_),
    .Y(_06529_),
    .A1(\atari2600.tia.p5_l ),
    .A2(_06525_));
 sg13g2_o21ai_1 _23836_ (.B1(_06522_),
    .Y(_06530_),
    .A1(_06527_),
    .A2(_06529_));
 sg13g2_o21ai_1 _23837_ (.B1(net6576),
    .Y(_06531_),
    .A1(_06520_),
    .A2(_06530_));
 sg13g2_a21oi_1 _23838_ (.A1(_08557_),
    .A2(_06520_),
    .Y(_01023_),
    .B1(_06531_));
 sg13g2_a21oi_1 _23839_ (.A1(_06064_),
    .A2(_06452_),
    .Y(_06532_),
    .B1(_08712_));
 sg13g2_nand3_1 _23840_ (.B(\atari2600.tia.audc1[0] ),
    .C(_06062_),
    .A(net7325),
    .Y(_06533_));
 sg13g2_nor2_1 _23841_ (.A(\atari2600.tia.audc1[1] ),
    .B(_06060_),
    .Y(_06534_));
 sg13g2_nor2_1 _23842_ (.A(_08506_),
    .B(_06133_),
    .Y(_06535_));
 sg13g2_o21ai_1 _23843_ (.B1(\atari2600.tia.audc1[0] ),
    .Y(_06536_),
    .A1(_06534_),
    .A2(_06535_));
 sg13g2_nor3_1 _23844_ (.A(\atari2600.tia.audc1[1] ),
    .B(\atari2600.tia.audc1[0] ),
    .C(_06060_),
    .Y(_06537_));
 sg13g2_nor2_1 _23845_ (.A(_00154_),
    .B(_06537_),
    .Y(_06538_));
 sg13g2_and2_1 _23846_ (.A(_06536_),
    .B(_06538_),
    .X(_06539_));
 sg13g2_a22oi_1 _23847_ (.Y(_06540_),
    .B1(_06537_),
    .B2(_08492_),
    .A2(_06062_),
    .A1(\atari2600.tia.audc1[0] ));
 sg13g2_o21ai_1 _23848_ (.B1(_06540_),
    .Y(_06541_),
    .A1(\atari2600.tia.p5_r ),
    .A2(_06536_));
 sg13g2_o21ai_1 _23849_ (.B1(_06533_),
    .Y(_06542_),
    .A1(_06539_),
    .A2(_06541_));
 sg13g2_nor2_1 _23850_ (.A(_06065_),
    .B(_06542_),
    .Y(_06543_));
 sg13g2_o21ai_1 _23851_ (.B1(net6576),
    .Y(_06544_),
    .A1(net6509),
    .A2(_06532_));
 sg13g2_a21oi_1 _23852_ (.A1(_06532_),
    .A2(_06543_),
    .Y(_01024_),
    .B1(_06544_));
 sg13g2_o21ai_1 _23853_ (.B1(net2931),
    .Y(_06545_),
    .A1(net5246),
    .A2(_10064_));
 sg13g2_a21oi_1 _23854_ (.A1(_10065_),
    .A2(_06545_),
    .Y(_01025_),
    .B1(net6541));
 sg13g2_and2_1 _23855_ (.A(_09127_),
    .B(_05374_),
    .X(_06546_));
 sg13g2_o21ai_1 _23856_ (.B1(net6573),
    .Y(_06547_),
    .A1(net7169),
    .A2(_06546_));
 sg13g2_a21oi_1 _23857_ (.A1(net5799),
    .A2(_06546_),
    .Y(_01026_),
    .B1(_06547_));
 sg13g2_a21oi_1 _23858_ (.A1(_09127_),
    .A2(_09444_),
    .Y(_06548_),
    .B1(net7584));
 sg13g2_nor2_2 _23859_ (.A(net6504),
    .B(net6507),
    .Y(_06549_));
 sg13g2_nor2b_2 _23860_ (.A(_10069_),
    .B_N(_06549_),
    .Y(_06550_));
 sg13g2_and3_2 _23861_ (.X(_06551_),
    .A(_10012_),
    .B(_10025_),
    .C(net5969));
 sg13g2_nor3_1 _23862_ (.A(net6531),
    .B(_06548_),
    .C(_06551_),
    .Y(_01027_));
 sg13g2_nor3_2 _23863_ (.A(net5203),
    .B(_09437_),
    .C(_05465_),
    .Y(_06552_));
 sg13g2_nor2_1 _23864_ (.A(net4191),
    .B(_06552_),
    .Y(_06553_));
 sg13g2_a21oi_1 _23865_ (.A1(net5712),
    .A2(_06552_),
    .Y(_01028_),
    .B1(_06553_));
 sg13g2_nor2_1 _23866_ (.A(net3199),
    .B(_06552_),
    .Y(_06554_));
 sg13g2_a21oi_1 _23867_ (.A1(net5668),
    .A2(_06552_),
    .Y(_01029_),
    .B1(_06554_));
 sg13g2_nor2_1 _23868_ (.A(net3888),
    .B(_06552_),
    .Y(_06555_));
 sg13g2_a21oi_1 _23869_ (.A1(net5591),
    .A2(_06552_),
    .Y(_01030_),
    .B1(_06555_));
 sg13g2_nor2_1 _23870_ (.A(net5246),
    .B(_09404_),
    .Y(_06556_));
 sg13g2_o21ai_1 _23871_ (.B1(net6568),
    .Y(_06557_),
    .A1(net7038),
    .A2(net5123));
 sg13g2_a21oi_1 _23872_ (.A1(net5798),
    .A2(net5123),
    .Y(_01031_),
    .B1(_06557_));
 sg13g2_o21ai_1 _23873_ (.B1(net6567),
    .Y(_06558_),
    .A1(net7172),
    .A2(net5124));
 sg13g2_a21oi_1 _23874_ (.A1(net5727),
    .A2(net5124),
    .Y(_01032_),
    .B1(_06558_));
 sg13g2_o21ai_1 _23875_ (.B1(net6567),
    .Y(_06559_),
    .A1(net7286),
    .A2(net5124));
 sg13g2_a21oi_1 _23876_ (.A1(net5704),
    .A2(net5124),
    .Y(_01033_),
    .B1(_06559_));
 sg13g2_o21ai_1 _23877_ (.B1(net6568),
    .Y(_06560_),
    .A1(net7287),
    .A2(net5124));
 sg13g2_a21oi_1 _23878_ (.A1(net5683),
    .A2(net5124),
    .Y(_01034_),
    .B1(_06560_));
 sg13g2_o21ai_1 _23879_ (.B1(net6558),
    .Y(_06561_),
    .A1(net7264),
    .A2(net5123));
 sg13g2_a21oi_1 _23880_ (.A1(net5602),
    .A2(net5123),
    .Y(_01035_),
    .B1(_06561_));
 sg13g2_o21ai_1 _23881_ (.B1(net6568),
    .Y(_06562_),
    .A1(net7222),
    .A2(net5123));
 sg13g2_a21oi_1 _23882_ (.A1(net5664),
    .A2(net5123),
    .Y(_01036_),
    .B1(_06562_));
 sg13g2_o21ai_1 _23883_ (.B1(net6567),
    .Y(_06563_),
    .A1(net7210),
    .A2(net5123));
 sg13g2_a21oi_1 _23884_ (.A1(net5638),
    .A2(net5123),
    .Y(_01037_),
    .B1(_06563_));
 sg13g2_nor2_1 _23885_ (.A(net5246),
    .B(_09307_),
    .Y(_06564_));
 sg13g2_o21ai_1 _23886_ (.B1(net6558),
    .Y(_06565_),
    .A1(net7443),
    .A2(net5121));
 sg13g2_a21oi_1 _23887_ (.A1(net5796),
    .A2(net5121),
    .Y(_01038_),
    .B1(_06565_));
 sg13g2_o21ai_1 _23888_ (.B1(net6569),
    .Y(_06566_),
    .A1(net7439),
    .A2(net5122));
 sg13g2_a21oi_1 _23889_ (.A1(net5727),
    .A2(net5122),
    .Y(_01039_),
    .B1(_06566_));
 sg13g2_o21ai_1 _23890_ (.B1(net6569),
    .Y(_06567_),
    .A1(net7385),
    .A2(net5122));
 sg13g2_a21oi_1 _23891_ (.A1(net5704),
    .A2(net5122),
    .Y(_01040_),
    .B1(_06567_));
 sg13g2_o21ai_1 _23892_ (.B1(net6568),
    .Y(_06568_),
    .A1(net7435),
    .A2(net5121));
 sg13g2_a21oi_1 _23893_ (.A1(net5684),
    .A2(net5121),
    .Y(_01041_),
    .B1(_06568_));
 sg13g2_o21ai_1 _23894_ (.B1(net6558),
    .Y(_06569_),
    .A1(net7389),
    .A2(net5121));
 sg13g2_a21oi_1 _23895_ (.A1(net5602),
    .A2(net5121),
    .Y(_01042_),
    .B1(_06569_));
 sg13g2_o21ai_1 _23896_ (.B1(net6568),
    .Y(_06570_),
    .A1(net7457),
    .A2(net5121));
 sg13g2_a21oi_1 _23897_ (.A1(net5664),
    .A2(net5121),
    .Y(_01043_),
    .B1(_06570_));
 sg13g2_o21ai_1 _23898_ (.B1(net6569),
    .Y(_06571_),
    .A1(net7453),
    .A2(net5122));
 sg13g2_a21oi_1 _23899_ (.A1(net5638),
    .A2(net5122),
    .Y(_01044_),
    .B1(_06571_));
 sg13g2_nor2_2 _23900_ (.A(net5524),
    .B(net5339),
    .Y(_06572_));
 sg13g2_and2_1 _23901_ (.A(_09127_),
    .B(_06572_),
    .X(_06573_));
 sg13g2_o21ai_1 _23902_ (.B1(net6568),
    .Y(_06574_),
    .A1(net7293),
    .A2(net5119));
 sg13g2_a21oi_1 _23903_ (.A1(net5798),
    .A2(net5119),
    .Y(_01045_),
    .B1(_06574_));
 sg13g2_o21ai_1 _23904_ (.B1(net6567),
    .Y(_06575_),
    .A1(net7355),
    .A2(net5119));
 sg13g2_a21oi_1 _23905_ (.A1(net5727),
    .A2(net5119),
    .Y(_01046_),
    .B1(_06575_));
 sg13g2_o21ai_1 _23906_ (.B1(net6574),
    .Y(_06576_),
    .A1(net7363),
    .A2(net5120));
 sg13g2_a21oi_1 _23907_ (.A1(net5704),
    .A2(net5120),
    .Y(_01047_),
    .B1(_06576_));
 sg13g2_o21ai_1 _23908_ (.B1(net6573),
    .Y(_06577_),
    .A1(net7436),
    .A2(net5120));
 sg13g2_a21oi_1 _23909_ (.A1(net5684),
    .A2(net5120),
    .Y(_01048_),
    .B1(_06577_));
 sg13g2_o21ai_1 _23910_ (.B1(net6573),
    .Y(_06578_),
    .A1(net7288),
    .A2(net5120));
 sg13g2_a21oi_1 _23911_ (.A1(net5603),
    .A2(net5120),
    .Y(_01049_),
    .B1(_06578_));
 sg13g2_o21ai_1 _23912_ (.B1(net6568),
    .Y(_06579_),
    .A1(net7380),
    .A2(net5119));
 sg13g2_a21oi_1 _23913_ (.A1(net5663),
    .A2(net5119),
    .Y(_01050_),
    .B1(_06579_));
 sg13g2_o21ai_1 _23914_ (.B1(net6568),
    .Y(_06580_),
    .A1(net7334),
    .A2(net5119));
 sg13g2_a21oi_1 _23915_ (.A1(net5638),
    .A2(net5119),
    .Y(_01051_),
    .B1(_06580_));
 sg13g2_nor2_1 _23916_ (.A(net5246),
    .B(_09343_),
    .Y(_06581_));
 sg13g2_o21ai_1 _23917_ (.B1(net6573),
    .Y(_06582_),
    .A1(net7302),
    .A2(net5117));
 sg13g2_a21oi_1 _23918_ (.A1(net5798),
    .A2(net5117),
    .Y(_01052_),
    .B1(_06582_));
 sg13g2_o21ai_1 _23919_ (.B1(net6573),
    .Y(_06583_),
    .A1(net7174),
    .A2(net5118));
 sg13g2_a21oi_1 _23920_ (.A1(net5727),
    .A2(net5118),
    .Y(_01053_),
    .B1(_06583_));
 sg13g2_o21ai_1 _23921_ (.B1(net6574),
    .Y(_06584_),
    .A1(net7220),
    .A2(net5118));
 sg13g2_a21oi_1 _23922_ (.A1(net5704),
    .A2(net5118),
    .Y(_01054_),
    .B1(_06584_));
 sg13g2_o21ai_1 _23923_ (.B1(net6573),
    .Y(_06585_),
    .A1(net7341),
    .A2(net5117));
 sg13g2_a21oi_1 _23924_ (.A1(net5684),
    .A2(net5117),
    .Y(_01055_),
    .B1(_06585_));
 sg13g2_o21ai_1 _23925_ (.B1(net6573),
    .Y(_06586_),
    .A1(net7387),
    .A2(net5117));
 sg13g2_a21oi_1 _23926_ (.A1(net5603),
    .A2(net5117),
    .Y(_01056_),
    .B1(_06586_));
 sg13g2_o21ai_1 _23927_ (.B1(net6573),
    .Y(_06587_),
    .A1(net7319),
    .A2(net5117));
 sg13g2_a21oi_1 _23928_ (.A1(net5663),
    .A2(net5117),
    .Y(_01057_),
    .B1(_06587_));
 sg13g2_o21ai_1 _23929_ (.B1(net6574),
    .Y(_06588_),
    .A1(net7049),
    .A2(net5118));
 sg13g2_a21oi_1 _23930_ (.A1(net5638),
    .A2(net5118),
    .Y(_01058_),
    .B1(_06588_));
 sg13g2_nor3_1 _23931_ (.A(net5432),
    .B(net5497),
    .C(net5217),
    .Y(_06589_));
 sg13g2_o21ai_1 _23932_ (.B1(net6558),
    .Y(_06590_),
    .A1(net7408),
    .A2(_06589_));
 sg13g2_a21oi_1 _23933_ (.A1(net5796),
    .A2(_06589_),
    .Y(_01059_),
    .B1(_06590_));
 sg13g2_and2_1 _23934_ (.A(_09398_),
    .B(net5218),
    .X(_06591_));
 sg13g2_o21ai_1 _23935_ (.B1(net6558),
    .Y(_06592_),
    .A1(net7483),
    .A2(_06591_));
 sg13g2_a21oi_1 _23936_ (.A1(net5796),
    .A2(_06591_),
    .Y(_01060_),
    .B1(_06592_));
 sg13g2_nor3_2 _23937_ (.A(net5339),
    .B(net5499),
    .C(net5217),
    .Y(_06593_));
 sg13g2_o21ai_1 _23938_ (.B1(net6565),
    .Y(_06594_),
    .A1(net7315),
    .A2(_06593_));
 sg13g2_a21oi_1 _23939_ (.A1(net5797),
    .A2(_06593_),
    .Y(_01061_),
    .B1(_06594_));
 sg13g2_nor2_1 _23940_ (.A(net5533),
    .B(net5269),
    .Y(_06595_));
 sg13g2_nand2b_2 _23941_ (.Y(_06596_),
    .B(_09301_),
    .A_N(net5533));
 sg13g2_and2_1 _23942_ (.A(_09172_),
    .B(_06595_),
    .X(_06597_));
 sg13g2_o21ai_1 _23943_ (.B1(net6555),
    .Y(_06598_),
    .A1(net7553),
    .A2(_06597_));
 sg13g2_a21oi_1 _23944_ (.A1(net5772),
    .A2(_06597_),
    .Y(_01062_),
    .B1(_06598_));
 sg13g2_nor2_2 _23945_ (.A(_09307_),
    .B(_06596_),
    .Y(_06599_));
 sg13g2_o21ai_1 _23946_ (.B1(net6561),
    .Y(_06600_),
    .A1(net7571),
    .A2(_06599_));
 sg13g2_a21oi_1 _23947_ (.A1(net5776),
    .A2(_06599_),
    .Y(_01063_),
    .B1(_06600_));
 sg13g2_nor2_1 _23948_ (.A(net5246),
    .B(_05506_),
    .Y(_06601_));
 sg13g2_o21ai_1 _23949_ (.B1(net6552),
    .Y(_06602_),
    .A1(net6668),
    .A2(_06601_));
 sg13g2_a21oi_1 _23950_ (.A1(net5703),
    .A2(_06601_),
    .Y(_01064_),
    .B1(_06602_));
 sg13g2_nor3_2 _23951_ (.A(net5246),
    .B(net5384),
    .C(net5497),
    .Y(_06603_));
 sg13g2_o21ai_1 _23952_ (.B1(net6550),
    .Y(_06604_),
    .A1(net7081),
    .A2(_06603_));
 sg13g2_a21oi_1 _23953_ (.A1(net5703),
    .A2(_06603_),
    .Y(_01065_),
    .B1(_06604_));
 sg13g2_nand2_1 _23954_ (.Y(_06605_),
    .A(net5776),
    .B(net5125));
 sg13g2_o21ai_1 _23955_ (.B1(_06605_),
    .Y(_06606_),
    .A1(net7589),
    .A2(net5126));
 sg13g2_nor2_1 _23956_ (.A(net6534),
    .B(_06606_),
    .Y(_01066_));
 sg13g2_o21ai_1 _23957_ (.B1(net6558),
    .Y(_06607_),
    .A1(net6479),
    .A2(net5126));
 sg13g2_a21oi_1 _23958_ (.A1(net5796),
    .A2(net5126),
    .Y(_01067_),
    .B1(_06607_));
 sg13g2_o21ai_1 _23959_ (.B1(net6566),
    .Y(_06608_),
    .A1(net7539),
    .A2(net5126));
 sg13g2_a21oi_1 _23960_ (.A1(net5727),
    .A2(net5126),
    .Y(_01068_),
    .B1(_06608_));
 sg13g2_o21ai_1 _23961_ (.B1(net6555),
    .Y(_06609_),
    .A1(net7364),
    .A2(net5128));
 sg13g2_a21oi_1 _23962_ (.A1(net5772),
    .A2(_05507_),
    .Y(_01069_),
    .B1(_06609_));
 sg13g2_nand2_1 _23963_ (.Y(_06610_),
    .A(net5792),
    .B(net5128));
 sg13g2_o21ai_1 _23964_ (.B1(_06610_),
    .Y(_06611_),
    .A1(net7371),
    .A2(net5128));
 sg13g2_nor2_1 _23965_ (.A(net6528),
    .B(_06611_),
    .Y(_01070_));
 sg13g2_o21ai_1 _23966_ (.B1(net6555),
    .Y(_06612_),
    .A1(net7360),
    .A2(_05507_));
 sg13g2_a21oi_1 _23967_ (.A1(net5722),
    .A2(net5128),
    .Y(_01071_),
    .B1(_06612_));
 sg13g2_o21ai_1 _23968_ (.B1(net6555),
    .Y(_06613_),
    .A1(net7390),
    .A2(net5128));
 sg13g2_a21oi_1 _23969_ (.A1(net5698),
    .A2(net5128),
    .Y(_01072_),
    .B1(_06613_));
 sg13g2_o21ai_1 _23970_ (.B1(net6555),
    .Y(_06614_),
    .A1(net7382),
    .A2(net5127));
 sg13g2_a21oi_1 _23971_ (.A1(net5683),
    .A2(net5127),
    .Y(_01073_),
    .B1(_06614_));
 sg13g2_o21ai_1 _23972_ (.B1(net6555),
    .Y(_06615_),
    .A1(net7320),
    .A2(net5127));
 sg13g2_a21oi_1 _23973_ (.A1(net5598),
    .A2(net5127),
    .Y(_01074_),
    .B1(_06615_));
 sg13g2_o21ai_1 _23974_ (.B1(net6555),
    .Y(_06616_),
    .A1(net7301),
    .A2(net5127));
 sg13g2_a21oi_1 _23975_ (.A1(net5661),
    .A2(net5127),
    .Y(_01075_),
    .B1(_06616_));
 sg13g2_o21ai_1 _23976_ (.B1(net6555),
    .Y(_06617_),
    .A1(net7370),
    .A2(net5128));
 sg13g2_a21oi_1 _23977_ (.A1(net5632),
    .A2(net5127),
    .Y(_01076_),
    .B1(_06617_));
 sg13g2_nor3_1 _23978_ (.A(net5384),
    .B(net5497),
    .C(net5217),
    .Y(_06618_));
 sg13g2_nand2_1 _23979_ (.Y(_06619_),
    .A(net5776),
    .B(net5115));
 sg13g2_o21ai_1 _23980_ (.B1(_06619_),
    .Y(_06620_),
    .A1(net7332),
    .A2(net5115));
 sg13g2_nor2_1 _23981_ (.A(net6535),
    .B(_06620_),
    .Y(_01077_));
 sg13g2_o21ai_1 _23982_ (.B1(net6563),
    .Y(_06621_),
    .A1(net6764),
    .A2(net5114));
 sg13g2_a21oi_1 _23983_ (.A1(net5797),
    .A2(net5115),
    .Y(_01078_),
    .B1(_06621_));
 sg13g2_o21ai_1 _23984_ (.B1(net6563),
    .Y(_06622_),
    .A1(net7289),
    .A2(net5115));
 sg13g2_a21oi_1 _23985_ (.A1(net5726),
    .A2(net5115),
    .Y(_01079_),
    .B1(_06622_));
 sg13g2_o21ai_1 _23986_ (.B1(net6563),
    .Y(_06623_),
    .A1(net7149),
    .A2(net5115));
 sg13g2_a21oi_1 _23987_ (.A1(net5703),
    .A2(net5114),
    .Y(_01080_),
    .B1(_06623_));
 sg13g2_o21ai_1 _23988_ (.B1(net6561),
    .Y(_06624_),
    .A1(net7263),
    .A2(net5114));
 sg13g2_a21oi_1 _23989_ (.A1(net5683),
    .A2(net5114),
    .Y(_01081_),
    .B1(_06624_));
 sg13g2_o21ai_1 _23990_ (.B1(net6561),
    .Y(_06625_),
    .A1(net4346),
    .A2(net5114));
 sg13g2_a21oi_1 _23991_ (.A1(net5598),
    .A2(net5114),
    .Y(_01082_),
    .B1(_06625_));
 sg13g2_nand2_1 _23992_ (.Y(_06626_),
    .A(net5662),
    .B(net5114));
 sg13g2_o21ai_1 _23993_ (.B1(_06626_),
    .Y(_06627_),
    .A1(net4704),
    .A2(net5114));
 sg13g2_nor2_1 _23994_ (.A(net6533),
    .B(_06627_),
    .Y(_01083_));
 sg13g2_nand2_1 _23995_ (.Y(_06628_),
    .A(net5632),
    .B(net5116));
 sg13g2_o21ai_1 _23996_ (.B1(_06628_),
    .Y(_06629_),
    .A1(net4574),
    .A2(net5116));
 sg13g2_nor2_1 _23997_ (.A(net6533),
    .B(_06629_),
    .Y(_01084_));
 sg13g2_a21oi_1 _23998_ (.A1(\atari2600.tia.vid_ypos[2] ),
    .A2(\atari2600.tia.vid_ypos[1] ),
    .Y(_06630_),
    .B1(\atari2600.tia.vid_ypos[3] ));
 sg13g2_nand2b_1 _23999_ (.Y(_06631_),
    .B(\atari2600.tia.vid_ypos[4] ),
    .A_N(_06630_));
 sg13g2_nand4_1 _24000_ (.B(_00130_),
    .C(_08701_),
    .A(_08570_),
    .Y(_06632_),
    .D(_06631_));
 sg13g2_nand3_1 _24001_ (.B(net6071),
    .C(_06632_),
    .A(net5758),
    .Y(_06633_));
 sg13g2_nand2_1 _24002_ (.Y(_06634_),
    .A(net6452),
    .B(_06633_));
 sg13g2_and2_1 _24003_ (.A(\atari2600.tia.pf_priority ),
    .B(net5707),
    .X(_06635_));
 sg13g2_nor2b_1 _24004_ (.A(net6070),
    .B_N(\atari2600.tia.colup1[0] ),
    .Y(_06636_));
 sg13g2_a21oi_1 _24005_ (.A1(\atari2600.tia.colup0[0] ),
    .A2(net6070),
    .Y(_06637_),
    .B1(_06636_));
 sg13g2_nor2_1 _24006_ (.A(net6479),
    .B(\atari2600.tia.colupf[0] ),
    .Y(_06638_));
 sg13g2_a21oi_1 _24007_ (.A1(net6479),
    .A2(_06637_),
    .Y(_06639_),
    .B1(_06638_));
 sg13g2_mux2_1 _24008_ (.A0(\atari2600.tia.colubk[0] ),
    .A1(_06639_),
    .S(net5707),
    .X(_06640_));
 sg13g2_mux2_1 _24009_ (.A0(\atari2600.tia.colup1[0] ),
    .A1(_06640_),
    .S(net5260),
    .X(_06641_));
 sg13g2_mux2_1 _24010_ (.A0(_06641_),
    .A1(\atari2600.tia.colup0[0] ),
    .S(net5290),
    .X(_06642_));
 sg13g2_mux2_1 _24011_ (.A0(_06642_),
    .A1(_06639_),
    .S(net5573),
    .X(_06643_));
 sg13g2_nand2b_1 _24012_ (.Y(_06644_),
    .B(net5284),
    .A_N(\atari2600.tia.colup1[0] ));
 sg13g2_and2_1 _24013_ (.A(net5287),
    .B(_06644_),
    .X(_06645_));
 sg13g2_o21ai_1 _24014_ (.B1(_06645_),
    .Y(_06646_),
    .A1(net5284),
    .A2(_06643_));
 sg13g2_nand4_1 _24015_ (.B(\atari2600.tia.colup0[0] ),
    .C(_09862_),
    .A(\atari2600.tia.enam0 ),
    .Y(_06647_),
    .D(_09876_));
 sg13g2_nand3_1 _24016_ (.B(_06646_),
    .C(_06647_),
    .A(net5537),
    .Y(_06648_));
 sg13g2_o21ai_1 _24017_ (.B1(_06648_),
    .Y(_06649_),
    .A1(net7302),
    .A2(net5537));
 sg13g2_o21ai_1 _24018_ (.B1(_06634_),
    .Y(_01085_),
    .A1(_06633_),
    .A2(_06649_));
 sg13g2_nor2b_1 _24019_ (.A(\atari2600.tia.colup0[1] ),
    .B_N(net5291),
    .Y(_06650_));
 sg13g2_nor3_1 _24020_ (.A(net5261),
    .B(net5574),
    .C(_06650_),
    .Y(_06651_));
 sg13g2_o21ai_1 _24021_ (.B1(\atari2600.tia.colup1[1] ),
    .Y(_06652_),
    .A1(net5285),
    .A2(_06651_));
 sg13g2_nand2b_1 _24022_ (.Y(_06653_),
    .B(\atari2600.tia.colup1[1] ),
    .A_N(net6068));
 sg13g2_a21oi_1 _24023_ (.A1(\atari2600.tia.colup0[1] ),
    .A2(net6069),
    .Y(_06654_),
    .B1(_08541_));
 sg13g2_a22oi_1 _24024_ (.Y(_06655_),
    .B1(_06653_),
    .B2(_06654_),
    .A2(_08547_),
    .A1(_08541_));
 sg13g2_nand2_1 _24025_ (.Y(_06656_),
    .A(net5708),
    .B(_06655_));
 sg13g2_inv_1 _24026_ (.Y(_06657_),
    .A(_06656_));
 sg13g2_o21ai_1 _24027_ (.B1(_06656_),
    .Y(_06658_),
    .A1(_08556_),
    .A2(net5708));
 sg13g2_a21oi_1 _24028_ (.A1(net5261),
    .A2(_06658_),
    .Y(_06659_),
    .B1(net5291));
 sg13g2_nor3_1 _24029_ (.A(net5573),
    .B(_06650_),
    .C(_06659_),
    .Y(_06660_));
 sg13g2_a21oi_1 _24030_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06657_),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_and2_1 _24031_ (.A(net5288),
    .B(_06652_),
    .X(_06662_));
 sg13g2_o21ai_1 _24032_ (.B1(_06662_),
    .Y(_06663_),
    .A1(net5285),
    .A2(_06661_));
 sg13g2_o21ai_1 _24033_ (.B1(net5538),
    .Y(_06664_),
    .A1(\atari2600.tia.colup0[1] ),
    .A2(net5288));
 sg13g2_nand2b_1 _24034_ (.Y(_06665_),
    .B(_06663_),
    .A_N(_06664_));
 sg13g2_o21ai_1 _24035_ (.B1(_06665_),
    .Y(_06666_),
    .A1(_08547_),
    .A2(net5538));
 sg13g2_mux2_1 _24036_ (.A0(_06666_),
    .A1(net6431),
    .S(_06633_),
    .X(_01086_));
 sg13g2_nor2b_1 _24037_ (.A(\atari2600.tia.colup0[2] ),
    .B_N(net5291),
    .Y(_06667_));
 sg13g2_nor3_1 _24038_ (.A(net5261),
    .B(net5574),
    .C(_06667_),
    .Y(_06668_));
 sg13g2_o21ai_1 _24039_ (.B1(\atari2600.tia.colup1[2] ),
    .Y(_06669_),
    .A1(net5285),
    .A2(_06668_));
 sg13g2_nand2b_1 _24040_ (.Y(_06670_),
    .B(\atari2600.tia.colup1[2] ),
    .A_N(net6069));
 sg13g2_a21oi_1 _24041_ (.A1(\atari2600.tia.colup0[2] ),
    .A2(net6069),
    .Y(_06671_),
    .B1(_08541_));
 sg13g2_a22oi_1 _24042_ (.Y(_06672_),
    .B1(_06670_),
    .B2(_06671_),
    .A2(_08546_),
    .A1(_08541_));
 sg13g2_nand2_1 _24043_ (.Y(_06673_),
    .A(net5707),
    .B(_06672_));
 sg13g2_inv_1 _24044_ (.Y(_06674_),
    .A(_06673_));
 sg13g2_o21ai_1 _24045_ (.B1(_06673_),
    .Y(_06675_),
    .A1(_08555_),
    .A2(net5708));
 sg13g2_a21oi_1 _24046_ (.A1(net5261),
    .A2(_06675_),
    .Y(_06676_),
    .B1(net5290));
 sg13g2_nor3_1 _24047_ (.A(net5573),
    .B(_06667_),
    .C(_06676_),
    .Y(_06677_));
 sg13g2_a21oi_1 _24048_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06674_),
    .Y(_06678_),
    .B1(_06677_));
 sg13g2_and2_1 _24049_ (.A(net5288),
    .B(_06669_),
    .X(_06679_));
 sg13g2_o21ai_1 _24050_ (.B1(_06679_),
    .Y(_06680_),
    .A1(net5285),
    .A2(_06678_));
 sg13g2_o21ai_1 _24051_ (.B1(net5538),
    .Y(_06681_),
    .A1(\atari2600.tia.colup0[2] ),
    .A2(net5288));
 sg13g2_nand2b_1 _24052_ (.Y(_06682_),
    .B(_06680_),
    .A_N(_06681_));
 sg13g2_o21ai_1 _24053_ (.B1(_06682_),
    .Y(_06683_),
    .A1(_08546_),
    .A2(net5538));
 sg13g2_mux2_1 _24054_ (.A0(_06683_),
    .A1(net6401),
    .S(_06633_),
    .X(_01087_));
 sg13g2_nor2b_1 _24055_ (.A(\atari2600.tia.colup0[3] ),
    .B_N(net5290),
    .Y(_06684_));
 sg13g2_nor3_1 _24056_ (.A(net5260),
    .B(net5573),
    .C(_06684_),
    .Y(_06685_));
 sg13g2_o21ai_1 _24057_ (.B1(\atari2600.tia.colup1[3] ),
    .Y(_06686_),
    .A1(net5284),
    .A2(_06685_));
 sg13g2_o21ai_1 _24058_ (.B1(\atari2600.tia.scorepf ),
    .Y(_06687_),
    .A1(_08550_),
    .A2(net6068));
 sg13g2_a21oi_1 _24059_ (.A1(\atari2600.tia.colup0[3] ),
    .A2(net6068),
    .Y(_06688_),
    .B1(_06687_));
 sg13g2_nor3_1 _24060_ (.A(_10041_),
    .B(_10045_),
    .C(_06688_),
    .Y(_06689_));
 sg13g2_o21ai_1 _24061_ (.B1(_06689_),
    .Y(_06690_),
    .A1(net6479),
    .A2(\atari2600.tia.colupf[3] ));
 sg13g2_inv_1 _24062_ (.Y(_06691_),
    .A(_06690_));
 sg13g2_o21ai_1 _24063_ (.B1(_06690_),
    .Y(_06692_),
    .A1(_08554_),
    .A2(net5707));
 sg13g2_a21oi_1 _24064_ (.A1(net5260),
    .A2(_06692_),
    .Y(_06693_),
    .B1(net5291));
 sg13g2_nor3_1 _24065_ (.A(net5574),
    .B(_06684_),
    .C(_06693_),
    .Y(_06694_));
 sg13g2_a21oi_1 _24066_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06691_),
    .Y(_06695_),
    .B1(_06694_));
 sg13g2_and2_1 _24067_ (.A(net5287),
    .B(_06686_),
    .X(_06696_));
 sg13g2_o21ai_1 _24068_ (.B1(_06696_),
    .Y(_06697_),
    .A1(net5284),
    .A2(_06695_));
 sg13g2_o21ai_1 _24069_ (.B1(net5537),
    .Y(_06698_),
    .A1(\atari2600.tia.colup0[3] ),
    .A2(net5287));
 sg13g2_nand2b_1 _24070_ (.Y(_06699_),
    .B(_06697_),
    .A_N(_06698_));
 sg13g2_o21ai_1 _24071_ (.B1(_06699_),
    .Y(_06700_),
    .A1(_08545_),
    .A2(net5538));
 sg13g2_mux2_1 _24072_ (.A0(_06700_),
    .A1(net6373),
    .S(_06633_),
    .X(_01088_));
 sg13g2_nor2b_1 _24073_ (.A(\atari2600.tia.colup0[4] ),
    .B_N(net5290),
    .Y(_06701_));
 sg13g2_nor3_1 _24074_ (.A(net5260),
    .B(net5573),
    .C(_06701_),
    .Y(_06702_));
 sg13g2_o21ai_1 _24075_ (.B1(\atari2600.tia.colup1[4] ),
    .Y(_06703_),
    .A1(net5284),
    .A2(_06702_));
 sg13g2_o21ai_1 _24076_ (.B1(net6479),
    .Y(_06704_),
    .A1(_08549_),
    .A2(net6068));
 sg13g2_a21oi_1 _24077_ (.A1(\atari2600.tia.colup0[4] ),
    .A2(net6070),
    .Y(_06705_),
    .B1(_06704_));
 sg13g2_nor3_1 _24078_ (.A(_10041_),
    .B(_10045_),
    .C(_06705_),
    .Y(_06706_));
 sg13g2_o21ai_1 _24079_ (.B1(_06706_),
    .Y(_06707_),
    .A1(net6479),
    .A2(\atari2600.tia.colupf[4] ));
 sg13g2_inv_1 _24080_ (.Y(_06708_),
    .A(_06707_));
 sg13g2_o21ai_1 _24081_ (.B1(_06707_),
    .Y(_06709_),
    .A1(_08553_),
    .A2(net5707));
 sg13g2_a21oi_1 _24082_ (.A1(net5260),
    .A2(_06709_),
    .Y(_06710_),
    .B1(net5290));
 sg13g2_nor3_1 _24083_ (.A(net5573),
    .B(_06701_),
    .C(_06710_),
    .Y(_06711_));
 sg13g2_a21oi_1 _24084_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06708_),
    .Y(_06712_),
    .B1(_06711_));
 sg13g2_and2_1 _24085_ (.A(net5287),
    .B(_06703_),
    .X(_06713_));
 sg13g2_o21ai_1 _24086_ (.B1(_06713_),
    .Y(_06714_),
    .A1(net5284),
    .A2(_06712_));
 sg13g2_o21ai_1 _24087_ (.B1(net5537),
    .Y(_06715_),
    .A1(\atari2600.tia.colup0[4] ),
    .A2(net5287));
 sg13g2_nand2b_1 _24088_ (.Y(_06716_),
    .B(_06714_),
    .A_N(_06715_));
 sg13g2_o21ai_1 _24089_ (.B1(_06716_),
    .Y(_06717_),
    .A1(_08544_),
    .A2(net5537));
 sg13g2_mux2_1 _24090_ (.A0(_06717_),
    .A1(net6337),
    .S(_06633_),
    .X(_01089_));
 sg13g2_nor2b_1 _24091_ (.A(\atari2600.tia.colup0[5] ),
    .B_N(net5290),
    .Y(_06718_));
 sg13g2_nor3_1 _24092_ (.A(net5260),
    .B(net5573),
    .C(_06718_),
    .Y(_06719_));
 sg13g2_o21ai_1 _24093_ (.B1(\atari2600.tia.colup1[5] ),
    .Y(_06720_),
    .A1(net5284),
    .A2(_06719_));
 sg13g2_o21ai_1 _24094_ (.B1(net6479),
    .Y(_06721_),
    .A1(_08548_),
    .A2(net6068));
 sg13g2_a21oi_1 _24095_ (.A1(\atari2600.tia.colup0[5] ),
    .A2(net6068),
    .Y(_06722_),
    .B1(_06721_));
 sg13g2_nor3_1 _24096_ (.A(_10041_),
    .B(_10045_),
    .C(_06722_),
    .Y(_06723_));
 sg13g2_o21ai_1 _24097_ (.B1(_06723_),
    .Y(_06724_),
    .A1(net6479),
    .A2(\atari2600.tia.colupf[5] ));
 sg13g2_inv_1 _24098_ (.Y(_06725_),
    .A(_06724_));
 sg13g2_o21ai_1 _24099_ (.B1(_06724_),
    .Y(_06726_),
    .A1(_08552_),
    .A2(net5707));
 sg13g2_a21oi_1 _24100_ (.A1(net5260),
    .A2(_06726_),
    .Y(_06727_),
    .B1(net5290));
 sg13g2_nor3_1 _24101_ (.A(net5573),
    .B(_06718_),
    .C(_06727_),
    .Y(_06728_));
 sg13g2_a21oi_1 _24102_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06725_),
    .Y(_06729_),
    .B1(_06728_));
 sg13g2_and2_1 _24103_ (.A(net5287),
    .B(_06720_),
    .X(_06730_));
 sg13g2_o21ai_1 _24104_ (.B1(_06730_),
    .Y(_06731_),
    .A1(net5284),
    .A2(_06729_));
 sg13g2_o21ai_1 _24105_ (.B1(net5537),
    .Y(_06732_),
    .A1(\atari2600.tia.colup0[5] ),
    .A2(net5287));
 sg13g2_nand2b_1 _24106_ (.Y(_06733_),
    .B(_06731_),
    .A_N(_06732_));
 sg13g2_o21ai_1 _24107_ (.B1(_06733_),
    .Y(_06734_),
    .A1(_08543_),
    .A2(net5537));
 sg13g2_mux2_1 _24108_ (.A0(_06734_),
    .A1(net6313),
    .S(_06633_),
    .X(_01090_));
 sg13g2_nor2b_1 _24109_ (.A(\atari2600.tia.colup0[6] ),
    .B_N(net5291),
    .Y(_06735_));
 sg13g2_nor3_1 _24110_ (.A(net5261),
    .B(net5574),
    .C(_06735_),
    .Y(_06736_));
 sg13g2_o21ai_1 _24111_ (.B1(\atari2600.tia.colup1[6] ),
    .Y(_06737_),
    .A1(net5285),
    .A2(_06736_));
 sg13g2_nand2b_1 _24112_ (.Y(_06738_),
    .B(\atari2600.tia.colup1[6] ),
    .A_N(net6068));
 sg13g2_a21oi_1 _24113_ (.A1(\atari2600.tia.colup0[6] ),
    .A2(net6068),
    .Y(_06739_),
    .B1(_08541_));
 sg13g2_a22oi_1 _24114_ (.Y(_06740_),
    .B1(_06738_),
    .B2(_06739_),
    .A2(_08542_),
    .A1(_08541_));
 sg13g2_nand2_1 _24115_ (.Y(_06741_),
    .A(net5707),
    .B(_06740_));
 sg13g2_inv_1 _24116_ (.Y(_06742_),
    .A(_06741_));
 sg13g2_o21ai_1 _24117_ (.B1(_06741_),
    .Y(_06743_),
    .A1(_08551_),
    .A2(net5707));
 sg13g2_a21oi_1 _24118_ (.A1(net5260),
    .A2(_06743_),
    .Y(_06744_),
    .B1(net5290));
 sg13g2_nor3_1 _24119_ (.A(net5574),
    .B(_06735_),
    .C(_06744_),
    .Y(_06745_));
 sg13g2_a21oi_1 _24120_ (.A1(\atari2600.tia.pf_priority ),
    .A2(_06742_),
    .Y(_06746_),
    .B1(_06745_));
 sg13g2_and2_1 _24121_ (.A(net5288),
    .B(_06737_),
    .X(_06747_));
 sg13g2_o21ai_1 _24122_ (.B1(_06747_),
    .Y(_06748_),
    .A1(net5285),
    .A2(_06746_));
 sg13g2_o21ai_1 _24123_ (.B1(net5538),
    .Y(_06749_),
    .A1(\atari2600.tia.colup0[6] ),
    .A2(net5288));
 sg13g2_nand2b_1 _24124_ (.Y(_06750_),
    .B(_06748_),
    .A_N(_06749_));
 sg13g2_o21ai_1 _24125_ (.B1(_06750_),
    .Y(_06751_),
    .A1(_08542_),
    .A2(net5537));
 sg13g2_mux2_1 _24126_ (.A0(_06751_),
    .A1(net6282),
    .S(_06633_),
    .X(_01091_));
 sg13g2_and2_2 _24127_ (.A(net5808),
    .B(net5116),
    .X(_06752_));
 sg13g2_mux2_1 _24128_ (.A0(net3639),
    .A1(\atari2600.tia.diag[104] ),
    .S(_06752_),
    .X(_01092_));
 sg13g2_mux2_1 _24129_ (.A0(net3918),
    .A1(\atari2600.tia.diag[105] ),
    .S(_06752_),
    .X(_01093_));
 sg13g2_mux2_1 _24130_ (.A0(net3656),
    .A1(\atari2600.tia.diag[106] ),
    .S(_06752_),
    .X(_01094_));
 sg13g2_mux2_1 _24131_ (.A0(net3812),
    .A1(\atari2600.tia.diag[107] ),
    .S(_06752_),
    .X(_01095_));
 sg13g2_mux2_1 _24132_ (.A0(net3665),
    .A1(\atari2600.tia.diag[108] ),
    .S(_06752_),
    .X(_01096_));
 sg13g2_mux2_1 _24133_ (.A0(net4189),
    .A1(\atari2600.tia.diag[109] ),
    .S(_06752_),
    .X(_01097_));
 sg13g2_mux2_1 _24134_ (.A0(net3533),
    .A1(\atari2600.tia.diag[110] ),
    .S(_06752_),
    .X(_01098_));
 sg13g2_mux2_1 _24135_ (.A0(net3536),
    .A1(\atari2600.tia.diag[111] ),
    .S(_06752_),
    .X(_01099_));
 sg13g2_nor2_1 _24136_ (.A(net5533),
    .B(_09365_),
    .Y(_06753_));
 sg13g2_nand2b_1 _24137_ (.Y(_06754_),
    .B(net5240),
    .A_N(net5533));
 sg13g2_a21oi_2 _24138_ (.B1(_06753_),
    .Y(_06755_),
    .A2(net5218),
    .A1(_10063_));
 sg13g2_o21ai_1 _24139_ (.B1(_06754_),
    .Y(_06756_),
    .A1(_10064_),
    .A2(net5217));
 sg13g2_o21ai_1 _24140_ (.B1(net6557),
    .Y(_06757_),
    .A1(net7481),
    .A2(net5057));
 sg13g2_nand2_2 _24141_ (.Y(_06758_),
    .A(_09365_),
    .B(net6071));
 sg13g2_nor2_2 _24142_ (.A(net6506),
    .B(_06758_),
    .Y(_06759_));
 sg13g2_nand2_1 _24143_ (.Y(_06760_),
    .A(\atari2600.tia.hmp0[0] ),
    .B(_08540_));
 sg13g2_xor2_1 _24144_ (.B(\atari2600.tia.diag[64] ),
    .A(net7410),
    .X(_06761_));
 sg13g2_a21oi_1 _24145_ (.A1(net5242),
    .A2(_06761_),
    .Y(_06762_),
    .B1(_06759_));
 sg13g2_a21oi_1 _24146_ (.A1(net5057),
    .A2(_06762_),
    .Y(_01100_),
    .B1(_06757_));
 sg13g2_o21ai_1 _24147_ (.B1(net6557),
    .Y(_06763_),
    .A1(net7536),
    .A2(net5057));
 sg13g2_a21oi_2 _24148_ (.B1(_06758_),
    .Y(_06764_),
    .A2(_10126_),
    .A1(_10124_));
 sg13g2_nor2b_1 _24149_ (.A(\atari2600.tia.hmp0[1] ),
    .B_N(\atari2600.tia.diag[65] ),
    .Y(_06765_));
 sg13g2_xnor2_1 _24150_ (.Y(_06766_),
    .A(\atari2600.tia.hmp0[1] ),
    .B(\atari2600.tia.diag[65] ));
 sg13g2_xor2_1 _24151_ (.B(_06766_),
    .A(_06760_),
    .X(_06767_));
 sg13g2_a21oi_1 _24152_ (.A1(net5240),
    .A2(_06767_),
    .Y(_06768_),
    .B1(_06764_));
 sg13g2_a21oi_1 _24153_ (.A1(net5057),
    .A2(_06768_),
    .Y(_01101_),
    .B1(_06763_));
 sg13g2_o21ai_1 _24154_ (.B1(net6553),
    .Y(_06769_),
    .A1(net7527),
    .A2(net5056));
 sg13g2_nand2_1 _24155_ (.Y(_06770_),
    .A(net6124),
    .B(net6067));
 sg13g2_a21oi_2 _24156_ (.B1(_06758_),
    .Y(_06771_),
    .A2(_06770_),
    .A1(_10135_));
 sg13g2_xnor2_1 _24157_ (.Y(_06772_),
    .A(\atari2600.tia.hmp0[2] ),
    .B(\atari2600.tia.diag[66] ));
 sg13g2_a21oi_1 _24158_ (.A1(_06760_),
    .A2(_06766_),
    .Y(_06773_),
    .B1(_06765_));
 sg13g2_nor2b_1 _24159_ (.A(_06773_),
    .B_N(_06772_),
    .Y(_06774_));
 sg13g2_xnor2_1 _24160_ (.Y(_06775_),
    .A(_06772_),
    .B(_06773_));
 sg13g2_a21oi_1 _24161_ (.A1(net5240),
    .A2(_06775_),
    .Y(_06776_),
    .B1(_06771_));
 sg13g2_a21oi_1 _24162_ (.A1(net5056),
    .A2(_06776_),
    .Y(_01102_),
    .B1(_06769_));
 sg13g2_o21ai_1 _24163_ (.B1(net6553),
    .Y(_06777_),
    .A1(net6276),
    .A2(net5056));
 sg13g2_xnor2_1 _24164_ (.Y(_06778_),
    .A(net6500),
    .B(_10130_));
 sg13g2_nor2_2 _24165_ (.A(_06758_),
    .B(_06778_),
    .Y(_06779_));
 sg13g2_xnor2_1 _24166_ (.Y(_06780_),
    .A(\atari2600.tia.hmp0[3] ),
    .B(net6276));
 sg13g2_a21oi_1 _24167_ (.A1(_08518_),
    .A2(\atari2600.tia.diag[66] ),
    .Y(_06781_),
    .B1(_06774_));
 sg13g2_nor2b_1 _24168_ (.A(_06781_),
    .B_N(_06780_),
    .Y(_06782_));
 sg13g2_xor2_1 _24169_ (.B(_06781_),
    .A(_06780_),
    .X(_06783_));
 sg13g2_nor2_1 _24170_ (.A(_09365_),
    .B(_06783_),
    .Y(_06784_));
 sg13g2_nor3_1 _24171_ (.A(_06755_),
    .B(_06779_),
    .C(_06784_),
    .Y(_06785_));
 sg13g2_nor2_1 _24172_ (.A(_06777_),
    .B(_06785_),
    .Y(_01103_));
 sg13g2_and3_1 _24173_ (.X(_06786_),
    .A(net6500),
    .B(\atari2600.tia.vid_xpos[4] ),
    .C(_06770_));
 sg13g2_a21oi_1 _24174_ (.A1(net6500),
    .A2(_06770_),
    .Y(_06787_),
    .B1(\atari2600.tia.vid_xpos[4] ));
 sg13g2_nor3_2 _24175_ (.A(_06758_),
    .B(_06786_),
    .C(_06787_),
    .Y(_06788_));
 sg13g2_xnor2_1 _24176_ (.Y(_06789_),
    .A(net6267),
    .B(net6274));
 sg13g2_a21oi_1 _24177_ (.A1(_08517_),
    .A2(net6276),
    .Y(_06790_),
    .B1(_06782_));
 sg13g2_nor2b_1 _24178_ (.A(_06790_),
    .B_N(_06789_),
    .Y(_06791_));
 sg13g2_nor2b_1 _24179_ (.A(_06789_),
    .B_N(_06790_),
    .Y(_06792_));
 sg13g2_nor3_1 _24180_ (.A(_09365_),
    .B(_06791_),
    .C(_06792_),
    .Y(_06793_));
 sg13g2_nor3_1 _24181_ (.A(_06755_),
    .B(_06788_),
    .C(_06793_),
    .Y(_06794_));
 sg13g2_o21ai_1 _24182_ (.B1(net6553),
    .Y(_06795_),
    .A1(net6274),
    .A2(net5056));
 sg13g2_nor2_1 _24183_ (.A(_06794_),
    .B(_06795_),
    .Y(_01104_));
 sg13g2_o21ai_1 _24184_ (.B1(net6552),
    .Y(_06796_),
    .A1(net6273),
    .A2(net5056));
 sg13g2_xnor2_1 _24185_ (.Y(_06797_),
    .A(_08661_),
    .B(_06786_));
 sg13g2_nor2_2 _24186_ (.A(_06758_),
    .B(_06797_),
    .Y(_06798_));
 sg13g2_a21oi_2 _24187_ (.B1(_06791_),
    .Y(_06799_),
    .A2(net6274),
    .A1(_08517_));
 sg13g2_nand2_1 _24188_ (.Y(_06800_),
    .A(net6267),
    .B(_08538_));
 sg13g2_xor2_1 _24189_ (.B(net6273),
    .A(net6267),
    .X(_06801_));
 sg13g2_o21ai_1 _24190_ (.B1(net5241),
    .Y(_06802_),
    .A1(_06799_),
    .A2(_06801_));
 sg13g2_a21oi_1 _24191_ (.A1(_06799_),
    .A2(_06801_),
    .Y(_06803_),
    .B1(_06802_));
 sg13g2_nor3_1 _24192_ (.A(_06755_),
    .B(_06798_),
    .C(_06803_),
    .Y(_06804_));
 sg13g2_nor2_1 _24193_ (.A(_06796_),
    .B(_06804_),
    .Y(_01105_));
 sg13g2_nand2_1 _24194_ (.Y(_06805_),
    .A(net6491),
    .B(_06786_));
 sg13g2_xnor2_1 _24195_ (.Y(_06806_),
    .A(net6484),
    .B(_06805_));
 sg13g2_nor2_2 _24196_ (.A(_06758_),
    .B(_06806_),
    .Y(_06807_));
 sg13g2_xnor2_1 _24197_ (.Y(_06808_),
    .A(net6267),
    .B(\atari2600.tia.diag[70] ));
 sg13g2_o21ai_1 _24198_ (.B1(_06799_),
    .Y(_06809_),
    .A1(net6267),
    .A2(_08538_));
 sg13g2_nand3_1 _24199_ (.B(_06808_),
    .C(_06809_),
    .A(_06800_),
    .Y(_06810_));
 sg13g2_a21o_1 _24200_ (.A2(_06809_),
    .A1(_06800_),
    .B1(_06808_),
    .X(_06811_));
 sg13g2_and3_1 _24201_ (.X(_06812_),
    .A(net5241),
    .B(_06810_),
    .C(_06811_));
 sg13g2_nor3_1 _24202_ (.A(_06755_),
    .B(_06807_),
    .C(_06812_),
    .Y(_06813_));
 sg13g2_o21ai_1 _24203_ (.B1(net6553),
    .Y(_06814_),
    .A1(net7544),
    .A2(net5056));
 sg13g2_nor2_1 _24204_ (.A(_06813_),
    .B(_06814_),
    .Y(_01106_));
 sg13g2_o21ai_1 _24205_ (.B1(net6562),
    .Y(_06815_),
    .A1(net6272),
    .A2(net5056));
 sg13g2_nor3_1 _24206_ (.A(net6480),
    .B(net6484),
    .C(_06805_),
    .Y(_06816_));
 sg13g2_o21ai_1 _24207_ (.B1(net6480),
    .Y(_06817_),
    .A1(net6484),
    .A2(_06805_));
 sg13g2_nand2b_1 _24208_ (.Y(_06818_),
    .B(_06817_),
    .A_N(_06816_));
 sg13g2_nor2_2 _24209_ (.A(_06758_),
    .B(_06818_),
    .Y(_06819_));
 sg13g2_o21ai_1 _24210_ (.B1(_06810_),
    .Y(_06820_),
    .A1(net6267),
    .A2(_08537_));
 sg13g2_xor2_1 _24211_ (.B(\atari2600.tia.diag[71] ),
    .A(net6267),
    .X(_06821_));
 sg13g2_xnor2_1 _24212_ (.Y(_06822_),
    .A(_06820_),
    .B(_06821_));
 sg13g2_a21oi_1 _24213_ (.A1(net5241),
    .A2(_06822_),
    .Y(_06823_),
    .B1(_06819_));
 sg13g2_a21oi_1 _24214_ (.A1(net5056),
    .A2(_06823_),
    .Y(_01107_),
    .B1(_06815_));
 sg13g2_a21o_2 _24215_ (.A2(net5218),
    .A1(_05374_),
    .B1(_06753_),
    .X(_06824_));
 sg13g2_o21ai_1 _24216_ (.B1(net6557),
    .Y(_06825_),
    .A1(net7550),
    .A2(net5055));
 sg13g2_nand2b_1 _24217_ (.Y(_06826_),
    .B(\atari2600.tia.hmp1[0] ),
    .A_N(\atari2600.tia.diag[56] ));
 sg13g2_xor2_1 _24218_ (.B(\atari2600.tia.diag[56] ),
    .A(net7397),
    .X(_06827_));
 sg13g2_a21oi_1 _24219_ (.A1(net5240),
    .A2(_06827_),
    .Y(_06828_),
    .B1(_06759_));
 sg13g2_a21oi_1 _24220_ (.A1(net5055),
    .A2(_06828_),
    .Y(_01108_),
    .B1(_06825_));
 sg13g2_o21ai_1 _24221_ (.B1(net6553),
    .Y(_06829_),
    .A1(net7555),
    .A2(net5055));
 sg13g2_nor2_1 _24222_ (.A(\atari2600.tia.hmp1[1] ),
    .B(_08536_),
    .Y(_06830_));
 sg13g2_xnor2_1 _24223_ (.Y(_06831_),
    .A(\atari2600.tia.hmp1[1] ),
    .B(\atari2600.tia.diag[57] ));
 sg13g2_xor2_1 _24224_ (.B(_06831_),
    .A(_06826_),
    .X(_06832_));
 sg13g2_a21oi_1 _24225_ (.A1(net5240),
    .A2(_06832_),
    .Y(_06833_),
    .B1(_06764_));
 sg13g2_a21oi_1 _24226_ (.A1(net5055),
    .A2(_06833_),
    .Y(_01109_),
    .B1(_06829_));
 sg13g2_o21ai_1 _24227_ (.B1(net6552),
    .Y(_06834_),
    .A1(net7586),
    .A2(net5055));
 sg13g2_xnor2_1 _24228_ (.Y(_06835_),
    .A(\atari2600.tia.hmp1[2] ),
    .B(\atari2600.tia.diag[58] ));
 sg13g2_a21oi_1 _24229_ (.A1(_06826_),
    .A2(_06831_),
    .Y(_06836_),
    .B1(_06830_));
 sg13g2_nor2b_1 _24230_ (.A(_06836_),
    .B_N(_06835_),
    .Y(_06837_));
 sg13g2_xnor2_1 _24231_ (.Y(_06838_),
    .A(_06835_),
    .B(_06836_));
 sg13g2_a21oi_1 _24232_ (.A1(net5240),
    .A2(_06838_),
    .Y(_06839_),
    .B1(_06771_));
 sg13g2_a21oi_1 _24233_ (.A1(net5055),
    .A2(_06839_),
    .Y(_01110_),
    .B1(_06834_));
 sg13g2_o21ai_1 _24234_ (.B1(net6564),
    .Y(_06840_),
    .A1(net6271),
    .A2(net5054));
 sg13g2_xnor2_1 _24235_ (.Y(_06841_),
    .A(net6266),
    .B(net6271));
 sg13g2_a21oi_2 _24236_ (.B1(_06837_),
    .Y(_06842_),
    .A2(\atari2600.tia.diag[58] ),
    .A1(_08516_));
 sg13g2_nor2b_1 _24237_ (.A(_06842_),
    .B_N(_06841_),
    .Y(_06843_));
 sg13g2_xnor2_1 _24238_ (.Y(_06844_),
    .A(_06841_),
    .B(_06842_));
 sg13g2_a21oi_1 _24239_ (.A1(net5243),
    .A2(_06844_),
    .Y(_06845_),
    .B1(_06779_));
 sg13g2_a21oi_1 _24240_ (.A1(net5054),
    .A2(_06845_),
    .Y(_01111_),
    .B1(_06840_));
 sg13g2_o21ai_1 _24241_ (.B1(net6564),
    .Y(_06846_),
    .A1(net6270),
    .A2(_06824_));
 sg13g2_xnor2_1 _24242_ (.Y(_06847_),
    .A(\atari2600.tia.hmp1[3] ),
    .B(net6270));
 sg13g2_a21oi_1 _24243_ (.A1(_08515_),
    .A2(\atari2600.tia.diag[59] ),
    .Y(_06848_),
    .B1(_06843_));
 sg13g2_nor2b_1 _24244_ (.A(_06848_),
    .B_N(_06847_),
    .Y(_06849_));
 sg13g2_xnor2_1 _24245_ (.Y(_06850_),
    .A(_06847_),
    .B(_06848_));
 sg13g2_a21oi_1 _24246_ (.A1(net5244),
    .A2(_06850_),
    .Y(_06851_),
    .B1(_06788_));
 sg13g2_a21oi_1 _24247_ (.A1(net5055),
    .A2(_06851_),
    .Y(_01112_),
    .B1(_06846_));
 sg13g2_o21ai_1 _24248_ (.B1(net6563),
    .Y(_06852_),
    .A1(net7421),
    .A2(net5054));
 sg13g2_a21oi_1 _24249_ (.A1(_08515_),
    .A2(\atari2600.tia.diag[60] ),
    .Y(_06853_),
    .B1(_06849_));
 sg13g2_nand2_1 _24250_ (.Y(_06854_),
    .A(net6266),
    .B(_08532_));
 sg13g2_xnor2_1 _24251_ (.Y(_06855_),
    .A(net6266),
    .B(\atari2600.tia.diag[61] ));
 sg13g2_xnor2_1 _24252_ (.Y(_06856_),
    .A(_06853_),
    .B(_06855_));
 sg13g2_a21oi_1 _24253_ (.A1(net5243),
    .A2(_06856_),
    .Y(_06857_),
    .B1(_06798_));
 sg13g2_a21oi_1 _24254_ (.A1(net5054),
    .A2(_06857_),
    .Y(_01113_),
    .B1(_06852_));
 sg13g2_o21ai_1 _24255_ (.B1(net6563),
    .Y(_06858_),
    .A1(net7570),
    .A2(net5054));
 sg13g2_xnor2_1 _24256_ (.Y(_06859_),
    .A(net6266),
    .B(\atari2600.tia.diag[62] ));
 sg13g2_o21ai_1 _24257_ (.B1(_06853_),
    .Y(_06860_),
    .A1(net6266),
    .A2(_08532_));
 sg13g2_nand3_1 _24258_ (.B(_06859_),
    .C(_06860_),
    .A(_06854_),
    .Y(_06861_));
 sg13g2_a21oi_1 _24259_ (.A1(_06854_),
    .A2(_06860_),
    .Y(_06862_),
    .B1(_06859_));
 sg13g2_nor2_1 _24260_ (.A(_09365_),
    .B(_06862_),
    .Y(_06863_));
 sg13g2_a21oi_1 _24261_ (.A1(_06861_),
    .A2(_06863_),
    .Y(_06864_),
    .B1(_06807_));
 sg13g2_a21oi_1 _24262_ (.A1(net5054),
    .A2(_06864_),
    .Y(_01114_),
    .B1(_06858_));
 sg13g2_o21ai_1 _24263_ (.B1(net6563),
    .Y(_06865_),
    .A1(net7583),
    .A2(net5054));
 sg13g2_o21ai_1 _24264_ (.B1(_06861_),
    .Y(_06866_),
    .A1(net6266),
    .A2(_08531_));
 sg13g2_xor2_1 _24265_ (.B(\atari2600.tia.diag[63] ),
    .A(net6266),
    .X(_06867_));
 sg13g2_xnor2_1 _24266_ (.Y(_06868_),
    .A(_06866_),
    .B(_06867_));
 sg13g2_a21oi_1 _24267_ (.A1(net5243),
    .A2(_06868_),
    .Y(_06869_),
    .B1(_06819_));
 sg13g2_a21oi_1 _24268_ (.A1(net5054),
    .A2(_06869_),
    .Y(_01115_),
    .B1(_06865_));
 sg13g2_nor2_2 _24269_ (.A(net5269),
    .B(_09343_),
    .Y(_06870_));
 sg13g2_or2_1 _24270_ (.X(_06871_),
    .B(_09343_),
    .A(net5269));
 sg13g2_nand2_1 _24271_ (.Y(_06872_),
    .A(_06759_),
    .B(net5214));
 sg13g2_and2_1 _24272_ (.A(_09342_),
    .B(_06595_),
    .X(_06873_));
 sg13g2_a21oi_2 _24273_ (.B1(_06873_),
    .Y(_06874_),
    .A2(net5218),
    .A1(_09444_));
 sg13g2_a21o_2 _24274_ (.A2(net5218),
    .A1(_09444_),
    .B1(_06873_),
    .X(_06875_));
 sg13g2_nand2b_1 _24275_ (.Y(_06876_),
    .B(\atari2600.tia.hmm0[0] ),
    .A_N(\atari2600.tia.diag[48] ));
 sg13g2_xor2_1 _24276_ (.B(\atari2600.tia.diag[48] ),
    .A(net7118),
    .X(_06877_));
 sg13g2_a221oi_1 _24277_ (.B2(net5241),
    .C1(net5053),
    .B1(_06877_),
    .A1(net7481),
    .Y(_06878_),
    .A2(_06870_));
 sg13g2_o21ai_1 _24278_ (.B1(net6557),
    .Y(_06879_),
    .A1(net7499),
    .A2(_06875_));
 sg13g2_a21oi_1 _24279_ (.A1(_06872_),
    .A2(_06878_),
    .Y(_01116_),
    .B1(_06879_));
 sg13g2_nand2_1 _24280_ (.Y(_06880_),
    .A(_06764_),
    .B(_06871_));
 sg13g2_nor2b_1 _24281_ (.A(\atari2600.tia.hmm0[1] ),
    .B_N(\atari2600.tia.diag[49] ),
    .Y(_06881_));
 sg13g2_xnor2_1 _24282_ (.Y(_06882_),
    .A(\atari2600.tia.hmm0[1] ),
    .B(\atari2600.tia.diag[49] ));
 sg13g2_xor2_1 _24283_ (.B(_06882_),
    .A(_06876_),
    .X(_06883_));
 sg13g2_a221oi_1 _24284_ (.B2(net5242),
    .C1(net5053),
    .B1(_06883_),
    .A1(net7536),
    .Y(_06884_),
    .A2(_06870_));
 sg13g2_o21ai_1 _24285_ (.B1(net6558),
    .Y(_06885_),
    .A1(net7560),
    .A2(_06875_));
 sg13g2_a21oi_1 _24286_ (.A1(_06880_),
    .A2(_06884_),
    .Y(_01117_),
    .B1(_06885_));
 sg13g2_xor2_1 _24287_ (.B(\atari2600.tia.diag[50] ),
    .A(\atari2600.tia.hmm0[2] ),
    .X(_06886_));
 sg13g2_a21oi_1 _24288_ (.A1(_06876_),
    .A2(_06882_),
    .Y(_06887_),
    .B1(_06881_));
 sg13g2_nor2_1 _24289_ (.A(_06886_),
    .B(_06887_),
    .Y(_06888_));
 sg13g2_xor2_1 _24290_ (.B(_06887_),
    .A(_06886_),
    .X(_06889_));
 sg13g2_or2_1 _24291_ (.X(_06890_),
    .B(\atari2600.tia.p0_w[3] ),
    .A(\atari2600.tia.diag[66] ));
 sg13g2_nand2_1 _24292_ (.Y(_06891_),
    .A(\atari2600.tia.diag[66] ),
    .B(\atari2600.tia.p0_w[3] ));
 sg13g2_nand3_1 _24293_ (.B(_06890_),
    .C(_06891_),
    .A(_06870_),
    .Y(_06892_));
 sg13g2_a221oi_1 _24294_ (.B2(net5241),
    .C1(net5053),
    .B1(_06889_),
    .A1(_06771_),
    .Y(_06893_),
    .A2(net5214));
 sg13g2_a221oi_1 _24295_ (.B2(_06893_),
    .C1(net6534),
    .B1(_06892_),
    .A1(_08530_),
    .Y(_01118_),
    .A2(net5053));
 sg13g2_nand2_1 _24296_ (.Y(_06894_),
    .A(_06779_),
    .B(net5214));
 sg13g2_xor2_1 _24297_ (.B(\atari2600.tia.diag[51] ),
    .A(\atari2600.tia.hmm0[3] ),
    .X(_06895_));
 sg13g2_a21oi_1 _24298_ (.A1(_08514_),
    .A2(\atari2600.tia.diag[50] ),
    .Y(_06896_),
    .B1(_06888_));
 sg13g2_nor2_1 _24299_ (.A(_06895_),
    .B(_06896_),
    .Y(_06897_));
 sg13g2_xor2_1 _24300_ (.B(_06896_),
    .A(_06895_),
    .X(_06898_));
 sg13g2_nand2_1 _24301_ (.Y(_06899_),
    .A(\atari2600.tia.diag[67] ),
    .B(\atari2600.tia.p0_w[4] ));
 sg13g2_xor2_1 _24302_ (.B(\atari2600.tia.p0_w[4] ),
    .A(net6276),
    .X(_06900_));
 sg13g2_nand2b_1 _24303_ (.Y(_06901_),
    .B(_06900_),
    .A_N(_06891_));
 sg13g2_xnor2_1 _24304_ (.Y(_06902_),
    .A(_06891_),
    .B(_06900_));
 sg13g2_a221oi_1 _24305_ (.B2(_06870_),
    .C1(net5053),
    .B1(_06902_),
    .A1(net5241),
    .Y(_06903_),
    .A2(_06898_));
 sg13g2_a221oi_1 _24306_ (.B2(_06903_),
    .C1(net6534),
    .B1(_06894_),
    .A1(_08529_),
    .Y(_01119_),
    .A2(net5053));
 sg13g2_nand2_1 _24307_ (.Y(_06904_),
    .A(_06788_),
    .B(net5214));
 sg13g2_nand2_1 _24308_ (.Y(_06905_),
    .A(net6274),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_xnor2_1 _24309_ (.Y(_06906_),
    .A(net6274),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_nand3_1 _24310_ (.B(_06901_),
    .C(_06906_),
    .A(_06899_),
    .Y(_06907_));
 sg13g2_a21oi_2 _24311_ (.B1(_06906_),
    .Y(_06908_),
    .A2(_06901_),
    .A1(_06899_));
 sg13g2_nor2_1 _24312_ (.A(net5214),
    .B(_06908_),
    .Y(_06909_));
 sg13g2_xnor2_1 _24313_ (.Y(_06910_),
    .A(\atari2600.tia.hmm0[3] ),
    .B(\atari2600.tia.diag[52] ));
 sg13g2_a21oi_1 _24314_ (.A1(_08513_),
    .A2(\atari2600.tia.diag[51] ),
    .Y(_06911_),
    .B1(_06897_));
 sg13g2_nor2b_1 _24315_ (.A(_06911_),
    .B_N(_06910_),
    .Y(_06912_));
 sg13g2_xnor2_1 _24316_ (.Y(_06913_),
    .A(_06910_),
    .B(_06911_));
 sg13g2_a221oi_1 _24317_ (.B2(net5241),
    .C1(net5053),
    .B1(_06913_),
    .A1(_06907_),
    .Y(_06914_),
    .A2(_06909_));
 sg13g2_o21ai_1 _24318_ (.B1(net6565),
    .Y(_06915_),
    .A1(net7510),
    .A2(_06875_));
 sg13g2_a21oi_1 _24319_ (.A1(_06904_),
    .A2(_06914_),
    .Y(_01120_),
    .B1(_06915_));
 sg13g2_nand2_1 _24320_ (.Y(_06916_),
    .A(_06798_),
    .B(net5214));
 sg13g2_a21oi_1 _24321_ (.A1(_08513_),
    .A2(\atari2600.tia.diag[52] ),
    .Y(_06917_),
    .B1(_06912_));
 sg13g2_nand2_1 _24322_ (.Y(_06918_),
    .A(_08513_),
    .B(net6268));
 sg13g2_nor2_1 _24323_ (.A(_08513_),
    .B(net6268),
    .Y(_06919_));
 sg13g2_xnor2_1 _24324_ (.Y(_06920_),
    .A(\atari2600.tia.hmm0[3] ),
    .B(net6268));
 sg13g2_xnor2_1 _24325_ (.Y(_06921_),
    .A(_06917_),
    .B(_06920_));
 sg13g2_a21oi_1 _24326_ (.A1(net6274),
    .A2(\atari2600.tia.p0_w[5] ),
    .Y(_06922_),
    .B1(_06908_));
 sg13g2_xnor2_1 _24327_ (.Y(_06923_),
    .A(net6273),
    .B(_06922_));
 sg13g2_a221oi_1 _24328_ (.B2(_06870_),
    .C1(_06874_),
    .B1(_06923_),
    .A1(net5242),
    .Y(_06924_),
    .A2(_06921_));
 sg13g2_o21ai_1 _24329_ (.B1(net6566),
    .Y(_06925_),
    .A1(net6268),
    .A2(_06875_));
 sg13g2_a21oi_1 _24330_ (.A1(_06916_),
    .A2(_06924_),
    .Y(_01121_),
    .B1(_06925_));
 sg13g2_nand2_1 _24331_ (.Y(_06926_),
    .A(_06807_),
    .B(net5214));
 sg13g2_nand2_1 _24332_ (.Y(_06927_),
    .A(net6273),
    .B(_06908_));
 sg13g2_o21ai_1 _24333_ (.B1(_06927_),
    .Y(_06928_),
    .A1(_00150_),
    .A2(_06905_));
 sg13g2_xnor2_1 _24334_ (.Y(_06929_),
    .A(_08537_),
    .B(_06928_));
 sg13g2_nor2b_1 _24335_ (.A(\atari2600.tia.hmm0[3] ),
    .B_N(\atari2600.tia.diag[54] ),
    .Y(_06930_));
 sg13g2_xnor2_1 _24336_ (.Y(_06931_),
    .A(\atari2600.tia.hmm0[3] ),
    .B(\atari2600.tia.diag[54] ));
 sg13g2_a21oi_1 _24337_ (.A1(_06917_),
    .A2(_06918_),
    .Y(_06932_),
    .B1(_06919_));
 sg13g2_xor2_1 _24338_ (.B(_06932_),
    .A(_06931_),
    .X(_06933_));
 sg13g2_a221oi_1 _24339_ (.B2(net5242),
    .C1(_06874_),
    .B1(_06933_),
    .A1(_06870_),
    .Y(_06934_),
    .A2(_06929_));
 sg13g2_o21ai_1 _24340_ (.B1(net6566),
    .Y(_06935_),
    .A1(net7502),
    .A2(_06875_));
 sg13g2_a21oi_1 _24341_ (.A1(_06926_),
    .A2(_06934_),
    .Y(_01122_),
    .B1(_06935_));
 sg13g2_nand2_1 _24342_ (.Y(_06936_),
    .A(_06819_),
    .B(net5214));
 sg13g2_a21oi_1 _24343_ (.A1(_06931_),
    .A2(_06932_),
    .Y(_06937_),
    .B1(_06930_));
 sg13g2_xnor2_1 _24344_ (.Y(_06938_),
    .A(\atari2600.tia.hmm0[3] ),
    .B(\atari2600.tia.diag[55] ));
 sg13g2_xnor2_1 _24345_ (.Y(_06939_),
    .A(_06937_),
    .B(_06938_));
 sg13g2_nand2b_1 _24346_ (.Y(_06940_),
    .B(_06928_),
    .A_N(_00149_));
 sg13g2_xnor2_1 _24347_ (.Y(_06941_),
    .A(\atari2600.tia.diag[71] ),
    .B(_06940_));
 sg13g2_a221oi_1 _24348_ (.B2(_06870_),
    .C1(_06874_),
    .B1(_06941_),
    .A1(net5242),
    .Y(_06942_),
    .A2(_06939_));
 sg13g2_a221oi_1 _24349_ (.B2(_06942_),
    .C1(net6534),
    .B1(_06936_),
    .A1(_08528_),
    .Y(_01123_),
    .A2(net5053));
 sg13g2_nor2_2 _24350_ (.A(net5268),
    .B(_09404_),
    .Y(_06943_));
 sg13g2_nand2_2 _24351_ (.Y(_06944_),
    .A(_09301_),
    .B(_09403_));
 sg13g2_nand2_1 _24352_ (.Y(_06945_),
    .A(_06759_),
    .B(net5213));
 sg13g2_a221oi_1 _24353_ (.B2(_09403_),
    .C1(_06753_),
    .B1(_06595_),
    .A1(_09401_),
    .Y(_06946_),
    .A2(net5218));
 sg13g2_nand2b_1 _24354_ (.Y(_06947_),
    .B(\atari2600.tia.hmm1[0] ),
    .A_N(\atari2600.tia.diag[40] ));
 sg13g2_xor2_1 _24355_ (.B(\atari2600.tia.diag[40] ),
    .A(net7396),
    .X(_06948_));
 sg13g2_a221oi_1 _24356_ (.B2(net5240),
    .C1(net5052),
    .B1(_06948_),
    .A1(net7550),
    .Y(_06949_),
    .A2(_06943_));
 sg13g2_a21oi_1 _24357_ (.A1(_09365_),
    .A2(net5213),
    .Y(_06950_),
    .B1(net5533));
 sg13g2_a21o_1 _24358_ (.A2(net5218),
    .A1(_09401_),
    .B1(_06950_),
    .X(_06951_));
 sg13g2_o21ai_1 _24359_ (.B1(net6556),
    .Y(_06952_),
    .A1(net7551),
    .A2(_06951_));
 sg13g2_a21oi_1 _24360_ (.A1(_06945_),
    .A2(_06949_),
    .Y(_01124_),
    .B1(_06952_));
 sg13g2_o21ai_1 _24361_ (.B1(net6556),
    .Y(_06953_),
    .A1(net7572),
    .A2(_06951_));
 sg13g2_nand2_1 _24362_ (.Y(_06954_),
    .A(_06764_),
    .B(net5213));
 sg13g2_nor2b_1 _24363_ (.A(\atari2600.tia.hmm1[1] ),
    .B_N(\atari2600.tia.diag[41] ),
    .Y(_06955_));
 sg13g2_xnor2_1 _24364_ (.Y(_06956_),
    .A(\atari2600.tia.hmm1[1] ),
    .B(\atari2600.tia.diag[41] ));
 sg13g2_xor2_1 _24365_ (.B(_06956_),
    .A(_06947_),
    .X(_06957_));
 sg13g2_a221oi_1 _24366_ (.B2(net5240),
    .C1(net5052),
    .B1(_06957_),
    .A1(net7555),
    .Y(_06958_),
    .A2(_06943_));
 sg13g2_a21oi_1 _24367_ (.A1(_06954_),
    .A2(_06958_),
    .Y(_01125_),
    .B1(_06953_));
 sg13g2_nand2_1 _24368_ (.Y(_06959_),
    .A(_06771_),
    .B(net5213));
 sg13g2_nand2_1 _24369_ (.Y(_06960_),
    .A(\atari2600.tia.diag[58] ),
    .B(\atari2600.tia.p1_w[3] ));
 sg13g2_xor2_1 _24370_ (.B(\atari2600.tia.p1_w[3] ),
    .A(\atari2600.tia.diag[58] ),
    .X(_06961_));
 sg13g2_nand2b_1 _24371_ (.Y(_06962_),
    .B(\atari2600.tia.diag[42] ),
    .A_N(\atari2600.tia.hmm1[2] ));
 sg13g2_xor2_1 _24372_ (.B(\atari2600.tia.diag[42] ),
    .A(\atari2600.tia.hmm1[2] ),
    .X(_06963_));
 sg13g2_a21oi_2 _24373_ (.B1(_06955_),
    .Y(_06964_),
    .A2(_06956_),
    .A1(_06947_));
 sg13g2_xor2_1 _24374_ (.B(_06964_),
    .A(_06963_),
    .X(_06965_));
 sg13g2_a221oi_1 _24375_ (.B2(net5241),
    .C1(net5052),
    .B1(_06965_),
    .A1(_06943_),
    .Y(_06966_),
    .A2(_06961_));
 sg13g2_a221oi_1 _24376_ (.B2(_06966_),
    .C1(net6533),
    .B1(_06959_),
    .A1(_08527_),
    .Y(_01126_),
    .A2(net5052));
 sg13g2_nand2_1 _24377_ (.Y(_06967_),
    .A(_06779_),
    .B(_06944_));
 sg13g2_xor2_1 _24378_ (.B(\atari2600.tia.diag[43] ),
    .A(net6265),
    .X(_06968_));
 sg13g2_o21ai_1 _24379_ (.B1(_06962_),
    .Y(_06969_),
    .A1(_06963_),
    .A2(_06964_));
 sg13g2_nand2b_1 _24380_ (.Y(_06970_),
    .B(_06969_),
    .A_N(_06968_));
 sg13g2_xnor2_1 _24381_ (.Y(_06971_),
    .A(_06968_),
    .B(_06969_));
 sg13g2_nand2_1 _24382_ (.Y(_06972_),
    .A(net6271),
    .B(\atari2600.tia.p1_w[4] ));
 sg13g2_xor2_1 _24383_ (.B(\atari2600.tia.p1_w[4] ),
    .A(net6271),
    .X(_06973_));
 sg13g2_nand2b_1 _24384_ (.Y(_06974_),
    .B(_06973_),
    .A_N(_06960_));
 sg13g2_xnor2_1 _24385_ (.Y(_06975_),
    .A(_06960_),
    .B(_06973_));
 sg13g2_a221oi_1 _24386_ (.B2(_06943_),
    .C1(net5051),
    .B1(_06975_),
    .A1(net5243),
    .Y(_06976_),
    .A2(_06971_));
 sg13g2_a221oi_1 _24387_ (.B2(_06976_),
    .C1(net6533),
    .B1(_06967_),
    .A1(_08526_),
    .Y(_01127_),
    .A2(net5051));
 sg13g2_nand2_1 _24388_ (.Y(_06977_),
    .A(_06788_),
    .B(net5213));
 sg13g2_xor2_1 _24389_ (.B(\atari2600.tia.diag[44] ),
    .A(net6265),
    .X(_06978_));
 sg13g2_o21ai_1 _24390_ (.B1(_06970_),
    .Y(_06979_),
    .A1(net6265),
    .A2(_08526_));
 sg13g2_nand2b_1 _24391_ (.Y(_06980_),
    .B(_06979_),
    .A_N(_06978_));
 sg13g2_xnor2_1 _24392_ (.Y(_06981_),
    .A(_06978_),
    .B(_06979_));
 sg13g2_nand2_1 _24393_ (.Y(_06982_),
    .A(net6270),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_xnor2_1 _24394_ (.Y(_06983_),
    .A(net6270),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_and3_1 _24395_ (.X(_06984_),
    .A(_06972_),
    .B(_06974_),
    .C(_06983_));
 sg13g2_a21oi_1 _24396_ (.A1(_06972_),
    .A2(_06974_),
    .Y(_06985_),
    .B1(_06983_));
 sg13g2_nor2_1 _24397_ (.A(_06984_),
    .B(_06985_),
    .Y(_06986_));
 sg13g2_a221oi_1 _24398_ (.B2(_06943_),
    .C1(net5051),
    .B1(_06986_),
    .A1(net5243),
    .Y(_06987_),
    .A2(_06981_));
 sg13g2_a221oi_1 _24399_ (.B2(_06987_),
    .C1(net6535),
    .B1(_06977_),
    .A1(_08525_),
    .Y(_01128_),
    .A2(net5052));
 sg13g2_nand2_1 _24400_ (.Y(_06988_),
    .A(_06798_),
    .B(net5213));
 sg13g2_o21ai_1 _24401_ (.B1(_06980_),
    .Y(_06989_),
    .A1(net6265),
    .A2(_08525_));
 sg13g2_nor2_1 _24402_ (.A(net6265),
    .B(_08524_),
    .Y(_06990_));
 sg13g2_nand2_1 _24403_ (.Y(_06991_),
    .A(net6265),
    .B(_08524_));
 sg13g2_nand2b_1 _24404_ (.Y(_06992_),
    .B(_06991_),
    .A_N(_06990_));
 sg13g2_xnor2_1 _24405_ (.Y(_06993_),
    .A(_06989_),
    .B(_06992_));
 sg13g2_a21oi_1 _24406_ (.A1(net6270),
    .A2(\atari2600.tia.p1_w[5] ),
    .Y(_06994_),
    .B1(_06985_));
 sg13g2_xnor2_1 _24407_ (.Y(_06995_),
    .A(net6269),
    .B(_06994_));
 sg13g2_a221oi_1 _24408_ (.B2(_06943_),
    .C1(net5051),
    .B1(_06995_),
    .A1(net5243),
    .Y(_06996_),
    .A2(_06993_));
 sg13g2_a221oi_1 _24409_ (.B2(_06996_),
    .C1(net6535),
    .B1(_06988_),
    .A1(_08524_),
    .Y(_01129_),
    .A2(net5051));
 sg13g2_nand2_1 _24410_ (.Y(_06997_),
    .A(_06807_),
    .B(net5213));
 sg13g2_xnor2_1 _24411_ (.Y(_06998_),
    .A(net6265),
    .B(\atari2600.tia.diag[46] ));
 sg13g2_o21ai_1 _24412_ (.B1(_06991_),
    .Y(_06999_),
    .A1(_06989_),
    .A2(_06990_));
 sg13g2_nand2b_1 _24413_ (.Y(_07000_),
    .B(_06998_),
    .A_N(_06999_));
 sg13g2_xnor2_1 _24414_ (.Y(_07001_),
    .A(_06998_),
    .B(_06999_));
 sg13g2_nand2_1 _24415_ (.Y(_07002_),
    .A(net6269),
    .B(_06985_));
 sg13g2_o21ai_1 _24416_ (.B1(_07002_),
    .Y(_07003_),
    .A1(_00146_),
    .A2(_06982_));
 sg13g2_nand2_1 _24417_ (.Y(_07004_),
    .A(\atari2600.tia.diag[62] ),
    .B(_07003_));
 sg13g2_xnor2_1 _24418_ (.Y(_07005_),
    .A(_08531_),
    .B(_07003_));
 sg13g2_a221oi_1 _24419_ (.B2(_06943_),
    .C1(net5051),
    .B1(_07005_),
    .A1(net5243),
    .Y(_07006_),
    .A2(_07001_));
 sg13g2_a221oi_1 _24420_ (.B2(_07006_),
    .C1(net6535),
    .B1(_06997_),
    .A1(_08523_),
    .Y(_01130_),
    .A2(net5051));
 sg13g2_nand2_1 _24421_ (.Y(_07007_),
    .A(_06819_),
    .B(net5213));
 sg13g2_o21ai_1 _24422_ (.B1(_07000_),
    .Y(_07008_),
    .A1(net6265),
    .A2(_08523_));
 sg13g2_xor2_1 _24423_ (.B(\atari2600.tia.diag[47] ),
    .A(\atari2600.tia.hmm1[3] ),
    .X(_07009_));
 sg13g2_xnor2_1 _24424_ (.Y(_07010_),
    .A(_07008_),
    .B(_07009_));
 sg13g2_xor2_1 _24425_ (.B(_07004_),
    .A(_00147_),
    .X(_07011_));
 sg13g2_a221oi_1 _24426_ (.B2(_06943_),
    .C1(net5051),
    .B1(_07011_),
    .A1(net5243),
    .Y(_07012_),
    .A2(_07010_));
 sg13g2_a221oi_1 _24427_ (.B2(_07012_),
    .C1(net6535),
    .B1(_07007_),
    .A1(_08522_),
    .Y(_01131_),
    .A2(net5052));
 sg13g2_o21ai_1 _24428_ (.B1(_06754_),
    .Y(_07013_),
    .A1(_09212_),
    .A2(net5217));
 sg13g2_o21ai_1 _24429_ (.B1(net6559),
    .Y(_07014_),
    .A1(net7531),
    .A2(net5050));
 sg13g2_nand2b_1 _24430_ (.Y(_07015_),
    .B(\atari2600.tia.hmbl[0] ),
    .A_N(\atari2600.tia.diag[32] ));
 sg13g2_xor2_1 _24431_ (.B(\atari2600.tia.diag[32] ),
    .A(net7383),
    .X(_07016_));
 sg13g2_a21oi_1 _24432_ (.A1(net5245),
    .A2(_07016_),
    .Y(_07017_),
    .B1(_06759_));
 sg13g2_a21oi_1 _24433_ (.A1(net5050),
    .A2(_07017_),
    .Y(_01132_),
    .B1(_07014_));
 sg13g2_o21ai_1 _24434_ (.B1(net6559),
    .Y(_07018_),
    .A1(net7567),
    .A2(net5050));
 sg13g2_nor2b_1 _24435_ (.A(\atari2600.tia.hmbl[1] ),
    .B_N(\atari2600.tia.diag[33] ),
    .Y(_07019_));
 sg13g2_xnor2_1 _24436_ (.Y(_07020_),
    .A(\atari2600.tia.hmbl[1] ),
    .B(\atari2600.tia.diag[33] ));
 sg13g2_xor2_1 _24437_ (.B(_07020_),
    .A(_07015_),
    .X(_07021_));
 sg13g2_a21oi_1 _24438_ (.A1(net5245),
    .A2(_07021_),
    .Y(_07022_),
    .B1(_06764_));
 sg13g2_a21oi_1 _24439_ (.A1(net5050),
    .A2(_07022_),
    .Y(_01133_),
    .B1(_07018_));
 sg13g2_o21ai_1 _24440_ (.B1(net6565),
    .Y(_07023_),
    .A1(net7519),
    .A2(net5050));
 sg13g2_xnor2_1 _24441_ (.Y(_07024_),
    .A(\atari2600.tia.hmbl[2] ),
    .B(\atari2600.tia.diag[34] ));
 sg13g2_a21oi_2 _24442_ (.B1(_07019_),
    .Y(_07025_),
    .A2(_07020_),
    .A1(_07015_));
 sg13g2_nor2b_1 _24443_ (.A(_07025_),
    .B_N(_07024_),
    .Y(_07026_));
 sg13g2_xnor2_1 _24444_ (.Y(_07027_),
    .A(_07024_),
    .B(_07025_));
 sg13g2_a21oi_1 _24445_ (.A1(net5242),
    .A2(_07027_),
    .Y(_07028_),
    .B1(_06771_));
 sg13g2_a21oi_1 _24446_ (.A1(net5050),
    .A2(_07028_),
    .Y(_01134_),
    .B1(_07023_));
 sg13g2_o21ai_1 _24447_ (.B1(net6565),
    .Y(_07029_),
    .A1(net7538),
    .A2(net5049));
 sg13g2_xnor2_1 _24448_ (.Y(_07030_),
    .A(net6264),
    .B(\atari2600.tia.diag[35] ));
 sg13g2_a21oi_1 _24449_ (.A1(_08512_),
    .A2(\atari2600.tia.diag[34] ),
    .Y(_07031_),
    .B1(_07026_));
 sg13g2_nor2b_1 _24450_ (.A(_07031_),
    .B_N(_07030_),
    .Y(_07032_));
 sg13g2_xnor2_1 _24451_ (.Y(_07033_),
    .A(_07030_),
    .B(_07031_));
 sg13g2_a21oi_1 _24452_ (.A1(net5242),
    .A2(_07033_),
    .Y(_07034_),
    .B1(_06779_));
 sg13g2_a21oi_1 _24453_ (.A1(net5049),
    .A2(_07034_),
    .Y(_01135_),
    .B1(_07029_));
 sg13g2_o21ai_1 _24454_ (.B1(net6566),
    .Y(_07035_),
    .A1(net7522),
    .A2(net5050));
 sg13g2_xnor2_1 _24455_ (.Y(_07036_),
    .A(net6264),
    .B(\atari2600.tia.diag[36] ));
 sg13g2_a21oi_1 _24456_ (.A1(_08511_),
    .A2(\atari2600.tia.diag[35] ),
    .Y(_07037_),
    .B1(_07032_));
 sg13g2_nor2b_1 _24457_ (.A(_07037_),
    .B_N(_07036_),
    .Y(_07038_));
 sg13g2_xnor2_1 _24458_ (.Y(_07039_),
    .A(_07036_),
    .B(_07037_));
 sg13g2_a21oi_1 _24459_ (.A1(net5244),
    .A2(_07039_),
    .Y(_07040_),
    .B1(_06788_));
 sg13g2_a21oi_1 _24460_ (.A1(_07013_),
    .A2(_07040_),
    .Y(_01136_),
    .B1(_07035_));
 sg13g2_o21ai_1 _24461_ (.B1(net6566),
    .Y(_07041_),
    .A1(net7530),
    .A2(net5049));
 sg13g2_a21oi_2 _24462_ (.B1(_07038_),
    .Y(_07042_),
    .A2(\atari2600.tia.diag[36] ),
    .A1(_08511_));
 sg13g2_nand2_1 _24463_ (.Y(_07043_),
    .A(net6264),
    .B(_08520_));
 sg13g2_xnor2_1 _24464_ (.Y(_07044_),
    .A(net6264),
    .B(\atari2600.tia.diag[37] ));
 sg13g2_xnor2_1 _24465_ (.Y(_07045_),
    .A(_07042_),
    .B(_07044_));
 sg13g2_a21oi_1 _24466_ (.A1(net5244),
    .A2(_07045_),
    .Y(_07046_),
    .B1(_06798_));
 sg13g2_a21oi_1 _24467_ (.A1(net5049),
    .A2(_07046_),
    .Y(_01137_),
    .B1(_07041_));
 sg13g2_o21ai_1 _24468_ (.B1(net6566),
    .Y(_07047_),
    .A1(net7485),
    .A2(net5049));
 sg13g2_xnor2_1 _24469_ (.Y(_07048_),
    .A(net6264),
    .B(\atari2600.tia.diag[38] ));
 sg13g2_o21ai_1 _24470_ (.B1(_07042_),
    .Y(_07049_),
    .A1(net6264),
    .A2(_08520_));
 sg13g2_nand3_1 _24471_ (.B(_07048_),
    .C(_07049_),
    .A(_07043_),
    .Y(_07050_));
 sg13g2_a21oi_1 _24472_ (.A1(_07043_),
    .A2(_07049_),
    .Y(_07051_),
    .B1(_07048_));
 sg13g2_nor2_1 _24473_ (.A(_09365_),
    .B(_07051_),
    .Y(_07052_));
 sg13g2_a21oi_1 _24474_ (.A1(_07050_),
    .A2(_07052_),
    .Y(_07053_),
    .B1(_06807_));
 sg13g2_a21oi_1 _24475_ (.A1(net5049),
    .A2(_07053_),
    .Y(_01138_),
    .B1(_07047_));
 sg13g2_o21ai_1 _24476_ (.B1(net6566),
    .Y(_07054_),
    .A1(net7466),
    .A2(net5049));
 sg13g2_o21ai_1 _24477_ (.B1(_07050_),
    .Y(_07055_),
    .A1(net6264),
    .A2(_08519_));
 sg13g2_xor2_1 _24478_ (.B(\atari2600.tia.diag[39] ),
    .A(net6264),
    .X(_07056_));
 sg13g2_xnor2_1 _24479_ (.Y(_07057_),
    .A(_07055_),
    .B(_07056_));
 sg13g2_a21oi_1 _24480_ (.A1(net5244),
    .A2(_07057_),
    .Y(_07058_),
    .B1(_06819_));
 sg13g2_a21oi_1 _24481_ (.A1(net5049),
    .A2(_07058_),
    .Y(_01139_),
    .B1(_07054_));
 sg13g2_nor3_2 _24482_ (.A(net5246),
    .B(net5339),
    .C(net5497),
    .Y(_07059_));
 sg13g2_o21ai_1 _24483_ (.B1(net6550),
    .Y(_07060_),
    .A1(net7032),
    .A2(net5113));
 sg13g2_a21oi_1 _24484_ (.A1(net5776),
    .A2(net5112),
    .Y(_01140_),
    .B1(_07060_));
 sg13g2_o21ai_1 _24485_ (.B1(net6550),
    .Y(_07061_),
    .A1(net7229),
    .A2(net5113));
 sg13g2_a21oi_1 _24486_ (.A1(net5796),
    .A2(net5112),
    .Y(_01141_),
    .B1(_07061_));
 sg13g2_o21ai_1 _24487_ (.B1(net6550),
    .Y(_07062_),
    .A1(net7156),
    .A2(net5112));
 sg13g2_a21oi_1 _24488_ (.A1(net5726),
    .A2(net5112),
    .Y(_01142_),
    .B1(_07062_));
 sg13g2_o21ai_1 _24489_ (.B1(net6550),
    .Y(_07063_),
    .A1(net7173),
    .A2(net5112));
 sg13g2_a21oi_1 _24490_ (.A1(net5703),
    .A2(net5112),
    .Y(_01143_),
    .B1(_07063_));
 sg13g2_o21ai_1 _24491_ (.B1(net6554),
    .Y(_07064_),
    .A1(net7265),
    .A2(net5113));
 sg13g2_a21oi_1 _24492_ (.A1(net5683),
    .A2(_07059_),
    .Y(_01144_),
    .B1(_07064_));
 sg13g2_o21ai_1 _24493_ (.B1(net6550),
    .Y(_07065_),
    .A1(net7160),
    .A2(net5113));
 sg13g2_a21oi_1 _24494_ (.A1(net5598),
    .A2(net5113),
    .Y(_01145_),
    .B1(_07065_));
 sg13g2_o21ai_1 _24495_ (.B1(net6550),
    .Y(_07066_),
    .A1(net7190),
    .A2(net5112));
 sg13g2_a21oi_1 _24496_ (.A1(net5662),
    .A2(net5112),
    .Y(_01146_),
    .B1(_07066_));
 sg13g2_o21ai_1 _24497_ (.B1(net6551),
    .Y(_07067_),
    .A1(net7273),
    .A2(net5113));
 sg13g2_a21oi_1 _24498_ (.A1(net5632),
    .A2(net5113),
    .Y(_01147_),
    .B1(_07067_));
 sg13g2_a21oi_2 _24499_ (.B1(_06596_),
    .Y(_07068_),
    .A2(_05506_),
    .A1(_10064_));
 sg13g2_nand2_2 _24500_ (.Y(_07069_),
    .A(_09301_),
    .B(_05505_));
 sg13g2_nand2_2 _24501_ (.Y(_07070_),
    .A(net5610),
    .B(_07069_));
 sg13g2_o21ai_1 _24502_ (.B1(net6556),
    .Y(_07071_),
    .A1(net7410),
    .A2(_07068_));
 sg13g2_a21oi_1 _24503_ (.A1(_07068_),
    .A2(_07070_),
    .Y(_01148_),
    .B1(_07071_));
 sg13g2_nand2_2 _24504_ (.Y(_07072_),
    .A(net5584),
    .B(_07069_));
 sg13g2_o21ai_1 _24505_ (.B1(net6556),
    .Y(_07073_),
    .A1(net7449),
    .A2(_07068_));
 sg13g2_a21oi_1 _24506_ (.A1(_07068_),
    .A2(_07072_),
    .Y(_01149_),
    .B1(_07073_));
 sg13g2_nand2_2 _24507_ (.Y(_07074_),
    .A(net5577),
    .B(_07069_));
 sg13g2_o21ai_1 _24508_ (.B1(net6556),
    .Y(_07075_),
    .A1(net7427),
    .A2(_07068_));
 sg13g2_a21oi_1 _24509_ (.A1(_07068_),
    .A2(_07074_),
    .Y(_01150_),
    .B1(_07075_));
 sg13g2_nand2_2 _24510_ (.Y(_07076_),
    .A(net5643),
    .B(_07069_));
 sg13g2_o21ai_1 _24511_ (.B1(net6552),
    .Y(_07077_),
    .A1(net7432),
    .A2(_07068_));
 sg13g2_a21oi_1 _24512_ (.A1(_07068_),
    .A2(_07076_),
    .Y(_01151_),
    .B1(_07077_));
 sg13g2_nor2_1 _24513_ (.A(_05374_),
    .B(_05505_),
    .Y(_07078_));
 sg13g2_nor2_2 _24514_ (.A(_06596_),
    .B(_07078_),
    .Y(_07079_));
 sg13g2_o21ai_1 _24515_ (.B1(net6556),
    .Y(_07080_),
    .A1(net7397),
    .A2(_07079_));
 sg13g2_a21oi_1 _24516_ (.A1(_07070_),
    .A2(_07079_),
    .Y(_01152_),
    .B1(_07080_));
 sg13g2_o21ai_1 _24517_ (.B1(net6552),
    .Y(_07081_),
    .A1(net7417),
    .A2(_07079_));
 sg13g2_a21oi_1 _24518_ (.A1(_07072_),
    .A2(_07079_),
    .Y(_01153_),
    .B1(_07081_));
 sg13g2_o21ai_1 _24519_ (.B1(net6552),
    .Y(_07082_),
    .A1(net7441),
    .A2(_07079_));
 sg13g2_a21oi_1 _24520_ (.A1(_07074_),
    .A2(_07079_),
    .Y(_01154_),
    .B1(_07082_));
 sg13g2_o21ai_1 _24521_ (.B1(net6552),
    .Y(_07083_),
    .A1(net7488),
    .A2(_07079_));
 sg13g2_a21oi_1 _24522_ (.A1(_07076_),
    .A2(_07079_),
    .Y(_01155_),
    .B1(_07083_));
 sg13g2_nor3_2 _24523_ (.A(_09355_),
    .B(_09358_),
    .C(_06596_),
    .Y(_07084_));
 sg13g2_nor2_1 _24524_ (.A(net7118),
    .B(_07084_),
    .Y(_07085_));
 sg13g2_a21oi_1 _24525_ (.A1(_07070_),
    .A2(_07084_),
    .Y(_07086_),
    .B1(net6528));
 sg13g2_nor2b_1 _24526_ (.A(_07085_),
    .B_N(_07086_),
    .Y(_01156_));
 sg13g2_nor2_1 _24527_ (.A(net7148),
    .B(_07084_),
    .Y(_07087_));
 sg13g2_a21oi_1 _24528_ (.A1(_07072_),
    .A2(_07084_),
    .Y(_07088_),
    .B1(net6529));
 sg13g2_nor2b_1 _24529_ (.A(_07087_),
    .B_N(_07088_),
    .Y(_01157_));
 sg13g2_nor2_1 _24530_ (.A(net7295),
    .B(_07084_),
    .Y(_07089_));
 sg13g2_a21oi_1 _24531_ (.A1(_07074_),
    .A2(_07084_),
    .Y(_07090_),
    .B1(net6529));
 sg13g2_nor2b_1 _24532_ (.A(_07089_),
    .B_N(_07090_),
    .Y(_01158_));
 sg13g2_o21ai_1 _24533_ (.B1(net6557),
    .Y(_07091_),
    .A1(net7578),
    .A2(_07084_));
 sg13g2_a21oi_1 _24534_ (.A1(_07076_),
    .A2(_07084_),
    .Y(_01159_),
    .B1(_07091_));
 sg13g2_nor2_2 _24535_ (.A(_09437_),
    .B(_06596_),
    .Y(_07092_));
 sg13g2_nor3_2 _24536_ (.A(net5530),
    .B(_09355_),
    .C(_06596_),
    .Y(_07093_));
 sg13g2_o21ai_1 _24537_ (.B1(net6557),
    .Y(_07094_),
    .A1(net7396),
    .A2(_07093_));
 sg13g2_a21oi_1 _24538_ (.A1(_07070_),
    .A2(_07092_),
    .Y(_01160_),
    .B1(_07094_));
 sg13g2_o21ai_1 _24539_ (.B1(net6556),
    .Y(_07095_),
    .A1(net7377),
    .A2(_07093_));
 sg13g2_a21oi_1 _24540_ (.A1(_07072_),
    .A2(_07092_),
    .Y(_01161_),
    .B1(_07095_));
 sg13g2_o21ai_1 _24541_ (.B1(net6556),
    .Y(_07096_),
    .A1(net7445),
    .A2(_07093_));
 sg13g2_a21oi_1 _24542_ (.A1(_07074_),
    .A2(_07092_),
    .Y(_01162_),
    .B1(_07096_));
 sg13g2_o21ai_1 _24543_ (.B1(net6560),
    .Y(_07097_),
    .A1(net7506),
    .A2(_07093_));
 sg13g2_a21oi_1 _24544_ (.A1(_07076_),
    .A2(_07092_),
    .Y(_01163_),
    .B1(_07097_));
 sg13g2_a21oi_2 _24545_ (.B1(_06596_),
    .Y(_07098_),
    .A2(_05506_),
    .A1(_09212_));
 sg13g2_o21ai_1 _24546_ (.B1(net6558),
    .Y(_07099_),
    .A1(net7383),
    .A2(_07098_));
 sg13g2_a21oi_1 _24547_ (.A1(_07070_),
    .A2(_07098_),
    .Y(_01164_),
    .B1(_07099_));
 sg13g2_nor2_1 _24548_ (.A(net7152),
    .B(_07098_),
    .Y(_07100_));
 sg13g2_a21oi_1 _24549_ (.A1(_07072_),
    .A2(_07098_),
    .Y(_07101_),
    .B1(net6529));
 sg13g2_nor2b_1 _24550_ (.A(_07100_),
    .B_N(_07101_),
    .Y(_01165_));
 sg13g2_nor2_1 _24551_ (.A(net7284),
    .B(_07098_),
    .Y(_07102_));
 sg13g2_a21oi_1 _24552_ (.A1(_07074_),
    .A2(_07098_),
    .Y(_07103_),
    .B1(net6529));
 sg13g2_nor2b_1 _24553_ (.A(_07102_),
    .B_N(_07103_),
    .Y(_01166_));
 sg13g2_nand2_1 _24554_ (.Y(_07104_),
    .A(_07076_),
    .B(_07098_));
 sg13g2_o21ai_1 _24555_ (.B1(_07104_),
    .Y(_07105_),
    .A1(net7419),
    .A2(_07098_));
 sg13g2_nor2_1 _24556_ (.A(net6529),
    .B(_07105_),
    .Y(_01167_));
 sg13g2_nand2_1 _24557_ (.Y(_07106_),
    .A(net3358),
    .B(_05613_));
 sg13g2_nand3_1 _24558_ (.B(net5402),
    .C(_09314_),
    .A(net6549),
    .Y(_07107_));
 sg13g2_o21ai_1 _24559_ (.B1(_07106_),
    .Y(_01168_),
    .A1(_06596_),
    .A2(_07107_));
 sg13g2_and2_2 _24560_ (.A(_09172_),
    .B(_05503_),
    .X(_07108_));
 sg13g2_nand2_1 _24561_ (.Y(_07109_),
    .A(net5777),
    .B(_07108_));
 sg13g2_o21ai_1 _24562_ (.B1(_07109_),
    .Y(_07110_),
    .A1(net7426),
    .A2(_07108_));
 sg13g2_nor2_1 _24563_ (.A(net6541),
    .B(_07110_),
    .Y(_01169_));
 sg13g2_o21ai_1 _24564_ (.B1(net6567),
    .Y(_07111_),
    .A1(net7532),
    .A2(_07108_));
 sg13g2_a21oi_1 _24565_ (.A1(net5798),
    .A2(_07108_),
    .Y(_01170_),
    .B1(_07111_));
 sg13g2_o21ai_1 _24566_ (.B1(net6567),
    .Y(_07112_),
    .A1(net6263),
    .A2(_07108_));
 sg13g2_a21oi_1 _24567_ (.A1(net5727),
    .A2(_07108_),
    .Y(_01171_),
    .B1(_07112_));
 sg13g2_o21ai_1 _24568_ (.B1(net6567),
    .Y(_07113_),
    .A1(net6262),
    .A2(_07108_));
 sg13g2_a21oi_1 _24569_ (.A1(net5704),
    .A2(_07108_),
    .Y(_01172_),
    .B1(_07113_));
 sg13g2_nor2_2 _24570_ (.A(_09307_),
    .B(net5217),
    .Y(_07114_));
 sg13g2_nand2_1 _24571_ (.Y(_07115_),
    .A(net5777),
    .B(_07114_));
 sg13g2_o21ai_1 _24572_ (.B1(_07115_),
    .Y(_07116_),
    .A1(net7525),
    .A2(_07114_));
 sg13g2_nor2_1 _24573_ (.A(net6538),
    .B(_07116_),
    .Y(_01173_));
 sg13g2_nand2_1 _24574_ (.Y(_07117_),
    .A(net5798),
    .B(_07114_));
 sg13g2_o21ai_1 _24575_ (.B1(_07117_),
    .Y(_07118_),
    .A1(net7529),
    .A2(_07114_));
 sg13g2_nor2_1 _24576_ (.A(net6538),
    .B(_07118_),
    .Y(_01174_));
 sg13g2_o21ai_1 _24577_ (.B1(net6574),
    .Y(_07119_),
    .A1(net7463),
    .A2(_07114_));
 sg13g2_a21oi_1 _24578_ (.A1(net5728),
    .A2(_07114_),
    .Y(_01175_),
    .B1(_07119_));
 sg13g2_nand2_1 _24579_ (.Y(_07120_),
    .A(net5703),
    .B(_07114_));
 sg13g2_o21ai_1 _24580_ (.B1(_07120_),
    .Y(_07121_),
    .A1(net7472),
    .A2(_07114_));
 sg13g2_nor2_1 _24581_ (.A(net6540),
    .B(_07121_),
    .Y(_01176_));
 sg13g2_nor2_2 _24582_ (.A(_09404_),
    .B(_05504_),
    .Y(_07122_));
 sg13g2_nand2_1 _24583_ (.Y(_07123_),
    .A(net5775),
    .B(_07122_));
 sg13g2_o21ai_1 _24584_ (.B1(_07123_),
    .Y(_07124_),
    .A1(net7279),
    .A2(_07122_));
 sg13g2_nor2_1 _24585_ (.A(net6530),
    .B(_07124_),
    .Y(_01177_));
 sg13g2_o21ai_1 _24586_ (.B1(net6571),
    .Y(_07125_),
    .A1(net7111),
    .A2(_07122_));
 sg13g2_a21oi_1 _24587_ (.A1(net5795),
    .A2(_07122_),
    .Y(_01178_),
    .B1(_07125_));
 sg13g2_nand2_1 _24588_ (.Y(_07126_),
    .A(net5725),
    .B(_07122_));
 sg13g2_o21ai_1 _24589_ (.B1(_07126_),
    .Y(_07127_),
    .A1(net7112),
    .A2(_07122_));
 sg13g2_nor2_1 _24590_ (.A(net6530),
    .B(_07127_),
    .Y(_01179_));
 sg13g2_o21ai_1 _24591_ (.B1(net6570),
    .Y(_07128_),
    .A1(net7333),
    .A2(_07122_));
 sg13g2_a21oi_1 _24592_ (.A1(net5702),
    .A2(_07122_),
    .Y(_01180_),
    .B1(_07128_));
 sg13g2_nor2_2 _24593_ (.A(_09363_),
    .B(_05504_),
    .Y(_07129_));
 sg13g2_o21ai_1 _24594_ (.B1(net6572),
    .Y(_07130_),
    .A1(net7331),
    .A2(_07129_));
 sg13g2_a21oi_1 _24595_ (.A1(net5777),
    .A2(_07129_),
    .Y(_01181_),
    .B1(_07130_));
 sg13g2_nand2_1 _24596_ (.Y(_07131_),
    .A(net5798),
    .B(_07129_));
 sg13g2_o21ai_1 _24597_ (.B1(_07131_),
    .Y(_07132_),
    .A1(net7378),
    .A2(_07129_));
 sg13g2_nor2_1 _24598_ (.A(net6530),
    .B(_07132_),
    .Y(_01182_));
 sg13g2_o21ai_1 _24599_ (.B1(net6572),
    .Y(_07133_),
    .A1(net7388),
    .A2(_07129_));
 sg13g2_a21oi_1 _24600_ (.A1(net5727),
    .A2(_07129_),
    .Y(_01183_),
    .B1(_07133_));
 sg13g2_nand2_1 _24601_ (.Y(_07134_),
    .A(net5702),
    .B(_07129_));
 sg13g2_o21ai_1 _24602_ (.B1(_07134_),
    .Y(_07135_),
    .A1(net7342),
    .A2(_07129_));
 sg13g2_nor2_1 _24603_ (.A(net6530),
    .B(_07135_),
    .Y(_01184_));
 sg13g2_and2_2 _24604_ (.A(net5218),
    .B(_06572_),
    .X(_07136_));
 sg13g2_nand2_1 _24605_ (.Y(_07137_),
    .A(net5777),
    .B(net5111));
 sg13g2_o21ai_1 _24606_ (.B1(_07137_),
    .Y(_07138_),
    .A1(net6261),
    .A2(net5111));
 sg13g2_nor2_1 _24607_ (.A(net6531),
    .B(_07138_),
    .Y(_01185_));
 sg13g2_nand2_1 _24608_ (.Y(_07139_),
    .A(net5798),
    .B(net5111));
 sg13g2_o21ai_1 _24609_ (.B1(_07139_),
    .Y(_07140_),
    .A1(net7503),
    .A2(net5111));
 sg13g2_nor2_1 _24610_ (.A(net6530),
    .B(_07140_),
    .Y(_01186_));
 sg13g2_nand2_1 _24611_ (.Y(_07141_),
    .A(net5727),
    .B(net5111));
 sg13g2_o21ai_1 _24612_ (.B1(_07141_),
    .Y(_07142_),
    .A1(net6260),
    .A2(net5111));
 sg13g2_nor2_1 _24613_ (.A(net6530),
    .B(_07142_),
    .Y(_01187_));
 sg13g2_o21ai_1 _24614_ (.B1(net6572),
    .Y(_07143_),
    .A1(net7467),
    .A2(net5111));
 sg13g2_a21oi_1 _24615_ (.A1(net5703),
    .A2(net5111),
    .Y(_01188_),
    .B1(_07143_));
 sg13g2_o21ai_1 _24616_ (.B1(net6572),
    .Y(_07144_),
    .A1(net7193),
    .A2(_07136_));
 sg13g2_a21oi_1 _24617_ (.A1(net5684),
    .A2(_07136_),
    .Y(_01189_),
    .B1(_07144_));
 sg13g2_nor3_2 _24618_ (.A(net5533),
    .B(net5267),
    .C(_09343_),
    .Y(_07145_));
 sg13g2_nor2_1 _24619_ (.A(_09343_),
    .B(net5217),
    .Y(_07146_));
 sg13g2_o21ai_1 _24620_ (.B1(net6574),
    .Y(_07147_),
    .A1(net7546),
    .A2(net5212));
 sg13g2_a21oi_1 _24621_ (.A1(net5777),
    .A2(net5212),
    .Y(_01190_),
    .B1(_07147_));
 sg13g2_o21ai_1 _24622_ (.B1(net6575),
    .Y(_07148_),
    .A1(net7500),
    .A2(net5212));
 sg13g2_a21oi_1 _24623_ (.A1(net5798),
    .A2(_07145_),
    .Y(_01191_),
    .B1(_07148_));
 sg13g2_o21ai_1 _24624_ (.B1(net6574),
    .Y(_07149_),
    .A1(net7528),
    .A2(net5212));
 sg13g2_a21oi_1 _24625_ (.A1(net5728),
    .A2(net5212),
    .Y(_01192_),
    .B1(_07149_));
 sg13g2_o21ai_1 _24626_ (.B1(net6574),
    .Y(_07150_),
    .A1(net7543),
    .A2(net5212));
 sg13g2_a21oi_1 _24627_ (.A1(net5703),
    .A2(net5212),
    .Y(_01193_),
    .B1(_07150_));
 sg13g2_o21ai_1 _24628_ (.B1(net6567),
    .Y(_07151_),
    .A1(net6592),
    .A2(net5212));
 sg13g2_a21oi_1 _24629_ (.A1(net5684),
    .A2(_07146_),
    .Y(_01194_),
    .B1(_07151_));
 sg13g2_nand2_1 _24630_ (.Y(_07152_),
    .A(\atari2600.tia.audio_left_counter[1] ),
    .B(_05957_));
 sg13g2_nand4_1 _24631_ (.B(_05955_),
    .C(_05963_),
    .A(_00095_),
    .Y(_07153_),
    .D(_07152_));
 sg13g2_nor2_1 _24632_ (.A(_05956_),
    .B(_07153_),
    .Y(_07154_));
 sg13g2_and4_1 _24633_ (.A(_05951_),
    .B(_05953_),
    .C(_05968_),
    .D(_07154_),
    .X(_07155_));
 sg13g2_nand3_1 _24634_ (.B(_05974_),
    .C(_07155_),
    .A(_05949_),
    .Y(_07156_));
 sg13g2_or4_1 _24635_ (.A(_05971_),
    .B(_05975_),
    .C(_05977_),
    .D(_07156_),
    .X(_07157_));
 sg13g2_nor4_1 _24636_ (.A(_05943_),
    .B(_05947_),
    .C(_05981_),
    .D(_07157_),
    .Y(_07158_));
 sg13g2_xnor2_1 _24637_ (.Y(_07159_),
    .A(_00111_),
    .B(_05932_));
 sg13g2_and4_2 _24638_ (.A(_05935_),
    .B(_05938_),
    .C(_07158_),
    .D(_07159_),
    .X(_07160_));
 sg13g2_nand2b_1 _24639_ (.Y(_07161_),
    .B(\atari2600.tia.p4_l ),
    .A_N(net4969));
 sg13g2_nand2_1 _24640_ (.Y(_07162_),
    .A(net7372),
    .B(net4969));
 sg13g2_nand3_1 _24641_ (.B(_07161_),
    .C(_07162_),
    .A(net6579),
    .Y(_01195_));
 sg13g2_a21oi_1 _24642_ (.A1(net6873),
    .A2(net4970),
    .Y(_07163_),
    .B1(net6539));
 sg13g2_o21ai_1 _24643_ (.B1(_07163_),
    .Y(_01196_),
    .A1(_08500_),
    .A2(net4969));
 sg13g2_nand2b_1 _24644_ (.Y(_07164_),
    .B(net6873),
    .A_N(net4970));
 sg13g2_nand2_1 _24645_ (.Y(_07165_),
    .A(net7136),
    .B(net4970));
 sg13g2_nand3_1 _24646_ (.B(_07164_),
    .C(_07165_),
    .A(net6579),
    .Y(_01197_));
 sg13g2_nand2b_1 _24647_ (.Y(_07166_),
    .B(net7136),
    .A_N(net4970));
 sg13g2_xor2_1 _24648_ (.B(\atari2600.tia.p4_l ),
    .A(\atari2600.tia.poly4_l.x[1] ),
    .X(_07167_));
 sg13g2_nand2_1 _24649_ (.Y(_07168_),
    .A(net4970),
    .B(_07167_));
 sg13g2_nand3_1 _24650_ (.B(_07166_),
    .C(_07168_),
    .A(net6579),
    .Y(_01198_));
 sg13g2_a21oi_1 _24651_ (.A1(net4456),
    .A2(net4969),
    .Y(_07169_),
    .B1(net6539));
 sg13g2_o21ai_1 _24652_ (.B1(_07169_),
    .Y(_01199_),
    .A1(_08499_),
    .A2(net4969));
 sg13g2_nand2b_1 _24653_ (.Y(_07170_),
    .B(net4456),
    .A_N(net4969));
 sg13g2_nand2_1 _24654_ (.Y(_07171_),
    .A(net6916),
    .B(net4969));
 sg13g2_nand3_1 _24655_ (.B(_07170_),
    .C(_07171_),
    .A(net6579),
    .Y(_01200_));
 sg13g2_a21oi_1 _24656_ (.A1(net7122),
    .A2(net4973),
    .Y(_07172_),
    .B1(net6539));
 sg13g2_o21ai_1 _24657_ (.B1(_07172_),
    .Y(_01201_),
    .A1(_08498_),
    .A2(net4973));
 sg13g2_nand2b_1 _24658_ (.Y(_07173_),
    .B(net7122),
    .A_N(net4973));
 sg13g2_nand2_1 _24659_ (.Y(_07174_),
    .A(net7141),
    .B(net4973));
 sg13g2_nand3_1 _24660_ (.B(_07173_),
    .C(_07174_),
    .A(net6579),
    .Y(_01202_));
 sg13g2_nand2b_1 _24661_ (.Y(_07175_),
    .B(net7141),
    .A_N(net4973));
 sg13g2_xor2_1 _24662_ (.B(\atari2600.tia.p5_l ),
    .A(net6916),
    .X(_07176_));
 sg13g2_nand2_1 _24663_ (.Y(_07177_),
    .A(net4973),
    .B(_07176_));
 sg13g2_nand3_1 _24664_ (.B(_07175_),
    .C(_07177_),
    .A(net6580),
    .Y(_01203_));
 sg13g2_a21oi_1 _24665_ (.A1(net7225),
    .A2(net4971),
    .Y(_07178_),
    .B1(net6539));
 sg13g2_o21ai_1 _24666_ (.B1(_07178_),
    .Y(_01204_),
    .A1(_08497_),
    .A2(net4969));
 sg13g2_nand2b_1 _24667_ (.Y(_07179_),
    .B(net7225),
    .A_N(net4974));
 sg13g2_nand2_1 _24668_ (.Y(_07180_),
    .A(net7272),
    .B(net4974));
 sg13g2_nand3_1 _24669_ (.B(_07179_),
    .C(_07180_),
    .A(net6580),
    .Y(_01205_));
 sg13g2_nand2b_1 _24670_ (.Y(_07181_),
    .B(\atari2600.tia.poly9_l.x[2] ),
    .A_N(net4974));
 sg13g2_nand2_1 _24671_ (.Y(_07182_),
    .A(net7153),
    .B(net4973));
 sg13g2_nand3_1 _24672_ (.B(_07181_),
    .C(_07182_),
    .A(net6580),
    .Y(_01206_));
 sg13g2_nand2b_1 _24673_ (.Y(_07183_),
    .B(net7153),
    .A_N(net4973));
 sg13g2_nand2_1 _24674_ (.Y(_07184_),
    .A(net7209),
    .B(net4971));
 sg13g2_nand3_1 _24675_ (.B(_07183_),
    .C(_07184_),
    .A(net6579),
    .Y(_01207_));
 sg13g2_a21oi_1 _24676_ (.A1(net7162),
    .A2(net4971),
    .Y(_07185_),
    .B1(net6539));
 sg13g2_o21ai_1 _24677_ (.B1(_07185_),
    .Y(_01208_),
    .A1(_08496_),
    .A2(net4971));
 sg13g2_nand2b_1 _24678_ (.Y(_07186_),
    .B(\atari2600.tia.poly9_l.x[5] ),
    .A_N(net4971));
 sg13g2_nand2_1 _24679_ (.Y(_07187_),
    .A(net6945),
    .B(net4972));
 sg13g2_nand3_1 _24680_ (.B(_07186_),
    .C(_07187_),
    .A(net6581),
    .Y(_01209_));
 sg13g2_nand2b_1 _24681_ (.Y(_07188_),
    .B(net6945),
    .A_N(net4972));
 sg13g2_nand2_1 _24682_ (.Y(_07189_),
    .A(net6979),
    .B(net4972));
 sg13g2_nand3_1 _24683_ (.B(_07188_),
    .C(_07189_),
    .A(net6581),
    .Y(_01210_));
 sg13g2_nand2b_1 _24684_ (.Y(_07190_),
    .B(\atari2600.tia.poly9_l.x[7] ),
    .A_N(net4971));
 sg13g2_nand2_1 _24685_ (.Y(_07191_),
    .A(net4511),
    .B(net4971));
 sg13g2_nand3_1 _24686_ (.B(_07190_),
    .C(_07191_),
    .A(net6580),
    .Y(_01211_));
 sg13g2_nand2b_1 _24687_ (.Y(_07192_),
    .B(net4511),
    .A_N(net4971));
 sg13g2_xor2_1 _24688_ (.B(net7252),
    .A(net7209),
    .X(_07193_));
 sg13g2_nand2_1 _24689_ (.Y(_07194_),
    .A(net4972),
    .B(_07193_));
 sg13g2_nand3_1 _24690_ (.B(_07192_),
    .C(_07194_),
    .A(net6580),
    .Y(_01212_));
 sg13g2_xnor2_1 _24691_ (.Y(_07195_),
    .A(_00126_),
    .B(_05932_));
 sg13g2_or2_1 _24692_ (.X(_07196_),
    .B(_05934_),
    .A(_08624_));
 sg13g2_nand2_1 _24693_ (.Y(_07197_),
    .A(_08624_),
    .B(_05934_));
 sg13g2_and2_1 _24694_ (.A(_00124_),
    .B(_05936_),
    .X(_07198_));
 sg13g2_nor2_1 _24695_ (.A(_00124_),
    .B(_05936_),
    .Y(_07199_));
 sg13g2_nor2_1 _24696_ (.A(_00123_),
    .B(_05939_),
    .Y(_07200_));
 sg13g2_nand2_1 _24697_ (.Y(_07201_),
    .A(_00123_),
    .B(_05939_));
 sg13g2_or2_1 _24698_ (.X(_07202_),
    .B(_05941_),
    .A(_00122_));
 sg13g2_nand2_1 _24699_ (.Y(_07203_),
    .A(_00121_),
    .B(_05945_));
 sg13g2_or2_1 _24700_ (.X(_07204_),
    .B(_05945_),
    .A(_00121_));
 sg13g2_nand2_1 _24701_ (.Y(_07205_),
    .A(_00120_),
    .B(_05944_));
 sg13g2_nor2_1 _24702_ (.A(_00120_),
    .B(_05944_),
    .Y(_07206_));
 sg13g2_nor2_1 _24703_ (.A(_00119_),
    .B(_05973_),
    .Y(_07207_));
 sg13g2_and2_1 _24704_ (.A(_00119_),
    .B(_05973_),
    .X(_07208_));
 sg13g2_xnor2_1 _24705_ (.Y(_07209_),
    .A(\atari2600.tia.audio_right_counter[1] ),
    .B(_05957_));
 sg13g2_xor2_1 _24706_ (.B(_05961_),
    .A(_00113_),
    .X(_07210_));
 sg13g2_xnor2_1 _24707_ (.Y(_07211_),
    .A(_00114_),
    .B(_05954_));
 sg13g2_nor4_1 _24708_ (.A(\atari2600.tia.audio_right_counter[0] ),
    .B(_07209_),
    .C(_07210_),
    .D(_07211_),
    .Y(_07212_));
 sg13g2_xnor2_1 _24709_ (.Y(_07213_),
    .A(_00115_),
    .B(_05952_));
 sg13g2_xnor2_1 _24710_ (.Y(_07214_),
    .A(_08621_),
    .B(_05950_));
 sg13g2_xnor2_1 _24711_ (.Y(_07215_),
    .A(_00117_),
    .B(_05948_));
 sg13g2_nand4_1 _24712_ (.B(_07213_),
    .C(_07214_),
    .A(_07212_),
    .Y(_07216_),
    .D(_07215_));
 sg13g2_a21oi_1 _24713_ (.A1(_00118_),
    .A2(_05970_),
    .Y(_07217_),
    .B1(_07216_));
 sg13g2_o21ai_1 _24714_ (.B1(_07217_),
    .Y(_07218_),
    .A1(_00118_),
    .A2(_05970_));
 sg13g2_nor4_1 _24715_ (.A(_07206_),
    .B(_07207_),
    .C(_07208_),
    .D(_07218_),
    .Y(_07219_));
 sg13g2_nand4_1 _24716_ (.B(_07204_),
    .C(_07205_),
    .A(_07203_),
    .Y(_07220_),
    .D(_07219_));
 sg13g2_a21oi_1 _24717_ (.A1(_00122_),
    .A2(_05941_),
    .Y(_07221_),
    .B1(_07220_));
 sg13g2_nand3_1 _24718_ (.B(_07202_),
    .C(_07221_),
    .A(_07201_),
    .Y(_07222_));
 sg13g2_nor4_1 _24719_ (.A(_07198_),
    .B(_07199_),
    .C(_07200_),
    .D(_07222_),
    .Y(_07223_));
 sg13g2_nand4_1 _24720_ (.B(_07196_),
    .C(_07197_),
    .A(_07195_),
    .Y(_07224_),
    .D(_07223_));
 sg13g2_inv_1 _24721_ (.Y(_07225_),
    .A(net4968));
 sg13g2_nand2_1 _24722_ (.Y(_07226_),
    .A(net7325),
    .B(net4968));
 sg13g2_nand2_1 _24723_ (.Y(_07227_),
    .A(\atari2600.tia.poly4_r.x[1] ),
    .B(net4962));
 sg13g2_nand3_1 _24724_ (.B(_07226_),
    .C(_07227_),
    .A(net6579),
    .Y(_01213_));
 sg13g2_a21oi_1 _24725_ (.A1(net7244),
    .A2(net4961),
    .Y(_07228_),
    .B1(net6539));
 sg13g2_o21ai_1 _24726_ (.B1(_07228_),
    .Y(_01214_),
    .A1(_08495_),
    .A2(net4962));
 sg13g2_mux2_1 _24727_ (.A0(net4435),
    .A1(net7244),
    .S(net4968),
    .X(_07229_));
 sg13g2_or2_1 _24728_ (.X(_01215_),
    .B(_07229_),
    .A(net6539));
 sg13g2_nand2_1 _24729_ (.Y(_07230_),
    .A(net4435),
    .B(net4968));
 sg13g2_xor2_1 _24730_ (.B(\atari2600.tia.p4_r ),
    .A(\atari2600.tia.poly4_r.x[1] ),
    .X(_07231_));
 sg13g2_nand2_1 _24731_ (.Y(_07232_),
    .A(net4962),
    .B(_07231_));
 sg13g2_nand3_1 _24732_ (.B(_07230_),
    .C(_07232_),
    .A(net6579),
    .Y(_01216_));
 sg13g2_a21oi_1 _24733_ (.A1(net6815),
    .A2(net4962),
    .Y(_07233_),
    .B1(net6537));
 sg13g2_o21ai_1 _24734_ (.B1(_07233_),
    .Y(_01217_),
    .A1(_08494_),
    .A2(net4962));
 sg13g2_a21oi_1 _24735_ (.A1(net6815),
    .A2(net4968),
    .Y(_07234_),
    .B1(net6537));
 sg13g2_o21ai_1 _24736_ (.B1(_07234_),
    .Y(_01218_),
    .A1(_08493_),
    .A2(_07224_));
 sg13g2_a21oi_1 _24737_ (.A1(net4866),
    .A2(net4961),
    .Y(_07235_),
    .B1(net6537));
 sg13g2_o21ai_1 _24738_ (.B1(_07235_),
    .Y(_01219_),
    .A1(_08493_),
    .A2(net4961));
 sg13g2_mux2_1 _24739_ (.A0(net6984),
    .A1(net4866),
    .S(net4967),
    .X(_07236_));
 sg13g2_or2_1 _24740_ (.X(_01220_),
    .B(_07236_),
    .A(net6536));
 sg13g2_nand2_1 _24741_ (.Y(_07237_),
    .A(net6984),
    .B(net4968));
 sg13g2_xor2_1 _24742_ (.B(\atari2600.tia.p5_r ),
    .A(\atari2600.tia.poly5_r.x[2] ),
    .X(_07238_));
 sg13g2_nand2_1 _24743_ (.Y(_07239_),
    .A(net4961),
    .B(_07238_));
 sg13g2_nand3_1 _24744_ (.B(_07237_),
    .C(_07239_),
    .A(net6576),
    .Y(_01221_));
 sg13g2_a21oi_1 _24745_ (.A1(net7257),
    .A2(net4961),
    .Y(_07240_),
    .B1(net6537));
 sg13g2_o21ai_1 _24746_ (.B1(_07240_),
    .Y(_01222_),
    .A1(_08492_),
    .A2(net4962));
 sg13g2_mux2_1 _24747_ (.A0(net7498),
    .A1(net7257),
    .S(net4968),
    .X(_07241_));
 sg13g2_or2_1 _24748_ (.X(_01223_),
    .B(_07241_),
    .A(net6536));
 sg13g2_mux2_1 _24749_ (.A0(net4441),
    .A1(net7498),
    .S(net4967),
    .X(_07242_));
 sg13g2_or2_1 _24750_ (.X(_01224_),
    .B(_07242_),
    .A(net6536));
 sg13g2_a21oi_1 _24751_ (.A1(net4441),
    .A2(net4967),
    .Y(_07243_),
    .B1(net6536));
 sg13g2_o21ai_1 _24752_ (.B1(_07243_),
    .Y(_01225_),
    .A1(_08491_),
    .A2(net4967));
 sg13g2_a21oi_1 _24753_ (.A1(net7205),
    .A2(net4961),
    .Y(_07244_),
    .B1(net6536));
 sg13g2_o21ai_1 _24754_ (.B1(_07244_),
    .Y(_01226_),
    .A1(_08491_),
    .A2(net4961));
 sg13g2_mux2_1 _24755_ (.A0(net7486),
    .A1(net7205),
    .S(net4967),
    .X(_07245_));
 sg13g2_or2_1 _24756_ (.X(_01227_),
    .B(_07245_),
    .A(net6536));
 sg13g2_mux2_1 _24757_ (.A0(net7496),
    .A1(net7486),
    .S(net4967),
    .X(_07246_));
 sg13g2_or2_1 _24758_ (.X(_01228_),
    .B(_07246_),
    .A(net6536));
 sg13g2_mux2_1 _24759_ (.A0(net4410),
    .A1(net7496),
    .S(net4967),
    .X(_07247_));
 sg13g2_or2_1 _24760_ (.X(_01229_),
    .B(_07247_),
    .A(net6536));
 sg13g2_xor2_1 _24761_ (.B(\atari2600.tia.p9_r ),
    .A(\atari2600.tia.poly9_r.x[4] ),
    .X(_07248_));
 sg13g2_nand2_1 _24762_ (.Y(_07249_),
    .A(net4410),
    .B(net4967));
 sg13g2_nand2_1 _24763_ (.Y(_07250_),
    .A(net4961),
    .B(_07248_));
 sg13g2_nand3_1 _24764_ (.B(_07249_),
    .C(_07250_),
    .A(net6576),
    .Y(_01230_));
 sg13g2_nor2_1 _24765_ (.A(_03091_),
    .B(net5248),
    .Y(_07251_));
 sg13g2_nor2_1 _24766_ (.A(net3306),
    .B(net5109),
    .Y(_07252_));
 sg13g2_a21oi_1 _24767_ (.A1(net5772),
    .A2(net5109),
    .Y(_01231_),
    .B1(_07252_));
 sg13g2_nor2_1 _24768_ (.A(net3528),
    .B(net5110),
    .Y(_07253_));
 sg13g2_a21oi_1 _24769_ (.A1(net5793),
    .A2(net5110),
    .Y(_01232_),
    .B1(_07253_));
 sg13g2_nor2_1 _24770_ (.A(net3152),
    .B(net5110),
    .Y(_07254_));
 sg13g2_a21oi_1 _24771_ (.A1(net5722),
    .A2(net5110),
    .Y(_01233_),
    .B1(_07254_));
 sg13g2_nor2_1 _24772_ (.A(net4014),
    .B(net5110),
    .Y(_07255_));
 sg13g2_a21oi_1 _24773_ (.A1(net5698),
    .A2(net5110),
    .Y(_01234_),
    .B1(_07255_));
 sg13g2_nor2_1 _24774_ (.A(net3146),
    .B(net5109),
    .Y(_07256_));
 sg13g2_a21oi_1 _24775_ (.A1(net5679),
    .A2(net5109),
    .Y(_01235_),
    .B1(_07256_));
 sg13g2_nor2_1 _24776_ (.A(net4135),
    .B(net5109),
    .Y(_07257_));
 sg13g2_a21oi_1 _24777_ (.A1(net5599),
    .A2(net5109),
    .Y(_01236_),
    .B1(_07257_));
 sg13g2_nor2_1 _24778_ (.A(net3278),
    .B(net5110),
    .Y(_07258_));
 sg13g2_a21oi_1 _24779_ (.A1(net5662),
    .A2(_07251_),
    .Y(_01237_),
    .B1(_07258_));
 sg13g2_nor2_1 _24780_ (.A(net4362),
    .B(net5109),
    .Y(_07259_));
 sg13g2_a21oi_1 _24781_ (.A1(net5633),
    .A2(net5109),
    .Y(_01238_),
    .B1(_07259_));
 sg13g2_o21ai_1 _24782_ (.B1(net6547),
    .Y(_07260_),
    .A1(_09303_),
    .A2(_03134_));
 sg13g2_nor3_1 _24783_ (.A(net5450),
    .B(net5132),
    .C(_07260_),
    .Y(_07261_));
 sg13g2_nand3_1 _24784_ (.B(net6547),
    .C(net5132),
    .A(net7028),
    .Y(_07262_));
 sg13g2_a21oi_1 _24785_ (.A1(\atari2600.input_switches[3] ),
    .A2(net6526),
    .Y(_07263_),
    .B1(_07261_));
 sg13g2_nand2_1 _24786_ (.Y(_01239_),
    .A(_07262_),
    .B(_07263_));
 sg13g2_nand2_1 _24787_ (.Y(_07264_),
    .A(_05368_),
    .B(_05402_));
 sg13g2_nand3_1 _24788_ (.B(net5809),
    .C(_07264_),
    .A(net3121),
    .Y(_07265_));
 sg13g2_o21ai_1 _24789_ (.B1(_07265_),
    .Y(_01240_),
    .A1(_05283_),
    .A2(_05363_));
 sg13g2_nor2_1 _24790_ (.A(net5263),
    .B(net5238),
    .Y(_07266_));
 sg13g2_nor2_1 _24791_ (.A(net3304),
    .B(net5107),
    .Y(_07267_));
 sg13g2_a21oi_1 _24792_ (.A1(net5764),
    .A2(net5107),
    .Y(_01241_),
    .B1(_07267_));
 sg13g2_nor2_1 _24793_ (.A(net3835),
    .B(net5107),
    .Y(_07268_));
 sg13g2_a21oi_1 _24794_ (.A1(net5784),
    .A2(net5107),
    .Y(_01242_),
    .B1(_07268_));
 sg13g2_nor2_1 _24795_ (.A(net3471),
    .B(net5107),
    .Y(_07269_));
 sg13g2_a21oi_1 _24796_ (.A1(net5714),
    .A2(net5107),
    .Y(_01243_),
    .B1(_07269_));
 sg13g2_nor2_1 _24797_ (.A(net3392),
    .B(net5107),
    .Y(_07270_));
 sg13g2_a21oi_1 _24798_ (.A1(net5687),
    .A2(net5108),
    .Y(_01244_),
    .B1(_07270_));
 sg13g2_nor2_1 _24799_ (.A(net3285),
    .B(net5108),
    .Y(_07271_));
 sg13g2_a21oi_1 _24800_ (.A1(net5671),
    .A2(net5108),
    .Y(_01245_),
    .B1(_07271_));
 sg13g2_nor2_1 _24801_ (.A(net3545),
    .B(net5108),
    .Y(_07272_));
 sg13g2_a21oi_1 _24802_ (.A1(net5586),
    .A2(net5108),
    .Y(_01246_),
    .B1(_07272_));
 sg13g2_nor2_1 _24803_ (.A(net4073),
    .B(_07266_),
    .Y(_07273_));
 sg13g2_a21oi_1 _24804_ (.A1(net5654),
    .A2(net5107),
    .Y(_01247_),
    .B1(_07273_));
 sg13g2_nor2_1 _24805_ (.A(net3452),
    .B(net5108),
    .Y(_07274_));
 sg13g2_a21oi_1 _24806_ (.A1(net5623),
    .A2(net5108),
    .Y(_01248_),
    .B1(_07274_));
 sg13g2_nand2b_1 _24807_ (.Y(_07275_),
    .B(net5250),
    .A_N(net5263));
 sg13g2_nand2_1 _24808_ (.Y(_07276_),
    .A(net2980),
    .B(net5211));
 sg13g2_o21ai_1 _24809_ (.B1(_07276_),
    .Y(_01249_),
    .A1(net5761),
    .A2(net5211));
 sg13g2_nand2_1 _24810_ (.Y(_07277_),
    .A(net2976),
    .B(net5211));
 sg13g2_o21ai_1 _24811_ (.B1(_07277_),
    .Y(_01250_),
    .A1(net5785),
    .A2(net5211));
 sg13g2_nand2_1 _24812_ (.Y(_07278_),
    .A(net2968),
    .B(net5211));
 sg13g2_o21ai_1 _24813_ (.B1(_07278_),
    .Y(_01251_),
    .A1(net5710),
    .A2(net5211));
 sg13g2_nand2_1 _24814_ (.Y(_07279_),
    .A(net3035),
    .B(net5210));
 sg13g2_o21ai_1 _24815_ (.B1(_07279_),
    .Y(_01252_),
    .A1(net5688),
    .A2(net5210));
 sg13g2_nand2_1 _24816_ (.Y(_07280_),
    .A(net2967),
    .B(net5211));
 sg13g2_o21ai_1 _24817_ (.B1(_07280_),
    .Y(_01253_),
    .A1(net5671),
    .A2(net5211));
 sg13g2_nand2_1 _24818_ (.Y(_07281_),
    .A(net2971),
    .B(net5210));
 sg13g2_o21ai_1 _24819_ (.B1(_07281_),
    .Y(_01254_),
    .A1(net5586),
    .A2(net5210));
 sg13g2_nand2_1 _24820_ (.Y(_07282_),
    .A(net3087),
    .B(net5210));
 sg13g2_o21ai_1 _24821_ (.B1(_07282_),
    .Y(_01255_),
    .A1(net5648),
    .A2(net5210));
 sg13g2_nand2_1 _24822_ (.Y(_07283_),
    .A(net2962),
    .B(net5210));
 sg13g2_o21ai_1 _24823_ (.B1(_07283_),
    .Y(_01256_),
    .A1(net5624),
    .A2(net5210));
 sg13g2_nor2_1 _24824_ (.A(net5263),
    .B(net5259),
    .Y(_07284_));
 sg13g2_nor2_1 _24825_ (.A(net3693),
    .B(net5209),
    .Y(_07285_));
 sg13g2_a21oi_1 _24826_ (.A1(net5761),
    .A2(net5209),
    .Y(_01257_),
    .B1(_07285_));
 sg13g2_nor2_1 _24827_ (.A(net3620),
    .B(net5209),
    .Y(_07286_));
 sg13g2_a21oi_1 _24828_ (.A1(net5784),
    .A2(net5209),
    .Y(_01258_),
    .B1(_07286_));
 sg13g2_nor2_1 _24829_ (.A(net3989),
    .B(net5209),
    .Y(_07287_));
 sg13g2_a21oi_1 _24830_ (.A1(net5714),
    .A2(net5209),
    .Y(_01259_),
    .B1(_07287_));
 sg13g2_nor2_1 _24831_ (.A(net4317),
    .B(net5208),
    .Y(_07288_));
 sg13g2_a21oi_1 _24832_ (.A1(net5687),
    .A2(net5208),
    .Y(_01260_),
    .B1(_07288_));
 sg13g2_nor2_1 _24833_ (.A(net3098),
    .B(net5209),
    .Y(_07289_));
 sg13g2_a21oi_1 _24834_ (.A1(net5671),
    .A2(net5209),
    .Y(_01261_),
    .B1(_07289_));
 sg13g2_nor2_1 _24835_ (.A(net3660),
    .B(net5208),
    .Y(_07290_));
 sg13g2_a21oi_1 _24836_ (.A1(net5586),
    .A2(net5208),
    .Y(_01262_),
    .B1(_07290_));
 sg13g2_nor2_1 _24837_ (.A(net3689),
    .B(net5208),
    .Y(_07291_));
 sg13g2_a21oi_1 _24838_ (.A1(net5647),
    .A2(net5208),
    .Y(_01263_),
    .B1(_07291_));
 sg13g2_nor2_1 _24839_ (.A(net3245),
    .B(net5208),
    .Y(_07292_));
 sg13g2_a21oi_1 _24840_ (.A1(net5624),
    .A2(net5208),
    .Y(_01264_),
    .B1(_07292_));
 sg13g2_and4_1 _24841_ (.A(net5562),
    .B(net5400),
    .C(_09413_),
    .D(_03026_),
    .X(_07293_));
 sg13g2_nor2_1 _24842_ (.A(net3191),
    .B(net5048),
    .Y(_07294_));
 sg13g2_a21oi_1 _24843_ (.A1(net5762),
    .A2(net5048),
    .Y(_01265_),
    .B1(_07294_));
 sg13g2_nor2_1 _24844_ (.A(net3239),
    .B(net5048),
    .Y(_07295_));
 sg13g2_a21oi_1 _24845_ (.A1(net5783),
    .A2(net5048),
    .Y(_01266_),
    .B1(_07295_));
 sg13g2_nor2_1 _24846_ (.A(net3030),
    .B(net5048),
    .Y(_07296_));
 sg13g2_a21oi_1 _24847_ (.A1(net5713),
    .A2(net5048),
    .Y(_01267_),
    .B1(_07296_));
 sg13g2_nor2_1 _24848_ (.A(net4041),
    .B(net5047),
    .Y(_07297_));
 sg13g2_a21oi_1 _24849_ (.A1(net5691),
    .A2(net5047),
    .Y(_01268_),
    .B1(_07297_));
 sg13g2_nor2_1 _24850_ (.A(net3451),
    .B(net5048),
    .Y(_07298_));
 sg13g2_a21oi_1 _24851_ (.A1(net5669),
    .A2(net5048),
    .Y(_01269_),
    .B1(_07298_));
 sg13g2_nor2_1 _24852_ (.A(net3676),
    .B(net5047),
    .Y(_07299_));
 sg13g2_a21oi_1 _24853_ (.A1(net5592),
    .A2(net5047),
    .Y(_01270_),
    .B1(_07299_));
 sg13g2_nor2_1 _24854_ (.A(net4300),
    .B(net5047),
    .Y(_07300_));
 sg13g2_a21oi_1 _24855_ (.A1(net5650),
    .A2(net5047),
    .Y(_01271_),
    .B1(_07300_));
 sg13g2_nor2_1 _24856_ (.A(net4392),
    .B(net5047),
    .Y(_07301_));
 sg13g2_a21oi_1 _24857_ (.A1(net5631),
    .A2(net5047),
    .Y(_01272_),
    .B1(_07301_));
 sg13g2_nor2_1 _24858_ (.A(net5263),
    .B(net5249),
    .Y(_07302_));
 sg13g2_nor2_1 _24859_ (.A(net4237),
    .B(net5207),
    .Y(_07303_));
 sg13g2_a21oi_1 _24860_ (.A1(net5761),
    .A2(net5207),
    .Y(_01273_),
    .B1(_07303_));
 sg13g2_nor2_1 _24861_ (.A(net4501),
    .B(net5207),
    .Y(_07304_));
 sg13g2_a21oi_1 _24862_ (.A1(net5785),
    .A2(net5207),
    .Y(_01274_),
    .B1(_07304_));
 sg13g2_nor2_1 _24863_ (.A(net4199),
    .B(net5207),
    .Y(_07305_));
 sg13g2_a21oi_1 _24864_ (.A1(net5710),
    .A2(net5207),
    .Y(_01275_),
    .B1(_07305_));
 sg13g2_nor2_1 _24865_ (.A(net4090),
    .B(net5206),
    .Y(_07306_));
 sg13g2_a21oi_1 _24866_ (.A1(net5687),
    .A2(net5206),
    .Y(_01276_),
    .B1(_07306_));
 sg13g2_nor2_1 _24867_ (.A(net4098),
    .B(net5207),
    .Y(_07307_));
 sg13g2_a21oi_1 _24868_ (.A1(net5671),
    .A2(net5207),
    .Y(_01277_),
    .B1(_07307_));
 sg13g2_nor2_1 _24869_ (.A(net3014),
    .B(net5206),
    .Y(_07308_));
 sg13g2_a21oi_1 _24870_ (.A1(net5586),
    .A2(net5206),
    .Y(_01278_),
    .B1(_07308_));
 sg13g2_nor2_1 _24871_ (.A(net4338),
    .B(net5206),
    .Y(_07309_));
 sg13g2_a21oi_1 _24872_ (.A1(net5647),
    .A2(net5206),
    .Y(_01279_),
    .B1(_07309_));
 sg13g2_nor2_1 _24873_ (.A(net3103),
    .B(net5206),
    .Y(_07310_));
 sg13g2_a21oi_1 _24874_ (.A1(net5624),
    .A2(net5206),
    .Y(_01280_),
    .B1(_07310_));
 sg13g2_nor2_2 _24875_ (.A(_09422_),
    .B(net5255),
    .Y(_07311_));
 sg13g2_nor2_1 _24876_ (.A(net3718),
    .B(net5045),
    .Y(_07312_));
 sg13g2_a21oi_1 _24877_ (.A1(net5759),
    .A2(net5045),
    .Y(_01281_),
    .B1(_07312_));
 sg13g2_nor2_1 _24878_ (.A(net3696),
    .B(net5045),
    .Y(_07313_));
 sg13g2_a21oi_1 _24879_ (.A1(net5780),
    .A2(net5045),
    .Y(_01282_),
    .B1(_07313_));
 sg13g2_nor2_1 _24880_ (.A(net3105),
    .B(net5046),
    .Y(_07314_));
 sg13g2_a21oi_1 _24881_ (.A1(net5709),
    .A2(net5046),
    .Y(_01283_),
    .B1(_07314_));
 sg13g2_nor2_1 _24882_ (.A(net4091),
    .B(net5046),
    .Y(_07315_));
 sg13g2_a21oi_1 _24883_ (.A1(net5686),
    .A2(net5046),
    .Y(_01284_),
    .B1(_07315_));
 sg13g2_nor2_1 _24884_ (.A(net3104),
    .B(net5045),
    .Y(_07316_));
 sg13g2_a21oi_1 _24885_ (.A1(net5666),
    .A2(net5045),
    .Y(_01285_),
    .B1(_07316_));
 sg13g2_nor2_1 _24886_ (.A(net3717),
    .B(net5046),
    .Y(_07317_));
 sg13g2_a21oi_1 _24887_ (.A1(net5585),
    .A2(net5046),
    .Y(_01286_),
    .B1(_07317_));
 sg13g2_nor2_1 _24888_ (.A(net3238),
    .B(net5045),
    .Y(_07318_));
 sg13g2_a21oi_1 _24889_ (.A1(net5649),
    .A2(net5045),
    .Y(_01287_),
    .B1(_07318_));
 sg13g2_nor2_1 _24890_ (.A(net3869),
    .B(net5046),
    .Y(_07319_));
 sg13g2_a21oi_1 _24891_ (.A1(net5622),
    .A2(net5046),
    .Y(_01288_),
    .B1(_07319_));
 sg13g2_nor2_2 _24892_ (.A(net5548),
    .B(_09420_),
    .Y(_07320_));
 sg13g2_nand2_2 _24893_ (.Y(_07321_),
    .A(net5556),
    .B(_09421_));
 sg13g2_nand2_2 _24894_ (.Y(_07322_),
    .A(net5252),
    .B(_07320_));
 sg13g2_mux2_1 _24895_ (.A0(net5740),
    .A1(net6686),
    .S(_07322_),
    .X(_01289_));
 sg13g2_mux2_1 _24896_ (.A0(net5745),
    .A1(net6804),
    .S(_07322_),
    .X(_01290_));
 sg13g2_mux2_1 _24897_ (.A0(net5616),
    .A1(net4680),
    .S(_07322_),
    .X(_01291_));
 sg13g2_mux2_1 _24898_ (.A0(net5611),
    .A1(net6812),
    .S(_07322_),
    .X(_01292_));
 sg13g2_mux2_1 _24899_ (.A0(net5607),
    .A1(net4916),
    .S(_07322_),
    .X(_01293_));
 sg13g2_mux2_1 _24900_ (.A0(net5580),
    .A1(net4832),
    .S(_07322_),
    .X(_01294_));
 sg13g2_mux2_1 _24901_ (.A0(net5575),
    .A1(net6796),
    .S(_07322_),
    .X(_01295_));
 sg13g2_mux2_1 _24902_ (.A0(net5641),
    .A1(net6708),
    .S(_07322_),
    .X(_01296_));
 sg13g2_nor2_1 _24903_ (.A(_09422_),
    .B(net5249),
    .Y(_07323_));
 sg13g2_nor2_1 _24904_ (.A(net4295),
    .B(net5043),
    .Y(_07324_));
 sg13g2_a21oi_1 _24905_ (.A1(net5759),
    .A2(net5043),
    .Y(_01297_),
    .B1(_07324_));
 sg13g2_nor2_1 _24906_ (.A(net3526),
    .B(net5043),
    .Y(_07325_));
 sg13g2_a21oi_1 _24907_ (.A1(net5780),
    .A2(net5043),
    .Y(_01298_),
    .B1(_07325_));
 sg13g2_nor2_1 _24908_ (.A(net3386),
    .B(net5044),
    .Y(_07326_));
 sg13g2_a21oi_1 _24909_ (.A1(net5709),
    .A2(net5044),
    .Y(_01299_),
    .B1(_07326_));
 sg13g2_nor2_1 _24910_ (.A(net3071),
    .B(net5044),
    .Y(_07327_));
 sg13g2_a21oi_1 _24911_ (.A1(net5688),
    .A2(net5044),
    .Y(_01300_),
    .B1(_07327_));
 sg13g2_nor2_1 _24912_ (.A(net3033),
    .B(net5043),
    .Y(_07328_));
 sg13g2_a21oi_1 _24913_ (.A1(net5667),
    .A2(net5043),
    .Y(_01301_),
    .B1(_07328_));
 sg13g2_nor2_1 _24914_ (.A(net3395),
    .B(net5044),
    .Y(_07329_));
 sg13g2_a21oi_1 _24915_ (.A1(net5585),
    .A2(_07323_),
    .Y(_01302_),
    .B1(_07329_));
 sg13g2_nor2_1 _24916_ (.A(net4305),
    .B(net5044),
    .Y(_07330_));
 sg13g2_a21oi_1 _24917_ (.A1(net5647),
    .A2(net5044),
    .Y(_01303_),
    .B1(_07330_));
 sg13g2_nor2_1 _24918_ (.A(net3896),
    .B(net5043),
    .Y(_07331_));
 sg13g2_a21oi_1 _24919_ (.A1(net5622),
    .A2(net5043),
    .Y(_01304_),
    .B1(_07331_));
 sg13g2_nand2_2 _24920_ (.Y(_07332_),
    .A(_09061_),
    .B(_05129_));
 sg13g2_mux2_1 _24921_ (.A0(_05132_),
    .A1(net6671),
    .S(_07332_),
    .X(_01305_));
 sg13g2_mux2_1 _24922_ (.A0(_05139_),
    .A1(net7123),
    .S(_07332_),
    .X(_01306_));
 sg13g2_mux2_1 _24923_ (.A0(_05146_),
    .A1(net4639),
    .S(_07332_),
    .X(_01307_));
 sg13g2_mux2_1 _24924_ (.A0(_05151_),
    .A1(net6631),
    .S(_07332_),
    .X(_01308_));
 sg13g2_mux2_1 _24925_ (.A0(_05153_),
    .A1(net4498),
    .S(_07332_),
    .X(_01309_));
 sg13g2_mux2_1 _24926_ (.A0(_05159_),
    .A1(net4732),
    .S(_07332_),
    .X(_01310_));
 sg13g2_mux2_1 _24927_ (.A0(_05166_),
    .A1(net4811),
    .S(_07332_),
    .X(_01311_));
 sg13g2_mux2_1 _24928_ (.A0(_05171_),
    .A1(net7039),
    .S(_07332_),
    .X(_01312_));
 sg13g2_nor3_2 _24929_ (.A(_09128_),
    .B(net5432),
    .C(net5497),
    .Y(_07333_));
 sg13g2_o21ai_1 _24930_ (.B1(net6551),
    .Y(_07334_),
    .A1(net7213),
    .A2(_07333_));
 sg13g2_a21oi_1 _24931_ (.A1(net5683),
    .A2(_07333_),
    .Y(_01313_),
    .B1(_07334_));
 sg13g2_o21ai_1 _24932_ (.B1(net6551),
    .Y(_07335_),
    .A1(net7282),
    .A2(_07333_));
 sg13g2_a21oi_1 _24933_ (.A1(net5598),
    .A2(_07333_),
    .Y(_01314_),
    .B1(_07335_));
 sg13g2_nand2_1 _24934_ (.Y(_07336_),
    .A(net5662),
    .B(_07333_));
 sg13g2_o21ai_1 _24935_ (.B1(_07336_),
    .Y(_07337_),
    .A1(net7221),
    .A2(_07333_));
 sg13g2_nor2_1 _24936_ (.A(net6528),
    .B(_07337_),
    .Y(_01315_));
 sg13g2_nand2_1 _24937_ (.Y(_07338_),
    .A(net5632),
    .B(_07333_));
 sg13g2_o21ai_1 _24938_ (.B1(_07338_),
    .Y(_07339_),
    .A1(net7235),
    .A2(_07333_));
 sg13g2_nor2_1 _24939_ (.A(net6528),
    .B(_07339_),
    .Y(_01316_));
 sg13g2_and2_2 _24940_ (.A(_09127_),
    .B(_09398_),
    .X(_07340_));
 sg13g2_o21ai_1 _24941_ (.B1(net6551),
    .Y(_07341_),
    .A1(net6980),
    .A2(net5105));
 sg13g2_a21oi_1 _24942_ (.A1(net5632),
    .A2(net5105),
    .Y(_01317_),
    .B1(_07341_));
 sg13g2_o21ai_1 _24943_ (.B1(net6551),
    .Y(_07342_),
    .A1(net7211),
    .A2(net5105));
 sg13g2_a21oi_1 _24944_ (.A1(net5661),
    .A2(net5105),
    .Y(_01318_),
    .B1(_07342_));
 sg13g2_o21ai_1 _24945_ (.B1(net6551),
    .Y(_07343_),
    .A1(net7256),
    .A2(net5106));
 sg13g2_a21oi_1 _24946_ (.A1(net5598),
    .A2(net5106),
    .Y(_01319_),
    .B1(_07343_));
 sg13g2_o21ai_1 _24947_ (.B1(net6552),
    .Y(_07344_),
    .A1(net7091),
    .A2(net5106));
 sg13g2_a21oi_1 _24948_ (.A1(net5683),
    .A2(net5106),
    .Y(_01320_),
    .B1(_07344_));
 sg13g2_nand2_1 _24949_ (.Y(_07345_),
    .A(net5703),
    .B(net5105));
 sg13g2_o21ai_1 _24950_ (.B1(_07345_),
    .Y(_07346_),
    .A1(net7198),
    .A2(net5105));
 sg13g2_nor2_1 _24951_ (.A(net6528),
    .B(_07346_),
    .Y(_01321_));
 sg13g2_nand2_1 _24952_ (.Y(_07347_),
    .A(net5726),
    .B(net5106));
 sg13g2_o21ai_1 _24953_ (.B1(_07347_),
    .Y(_07348_),
    .A1(net7317),
    .A2(net5106));
 sg13g2_nor2_1 _24954_ (.A(net6528),
    .B(_07348_),
    .Y(_01322_));
 sg13g2_nand2_1 _24955_ (.Y(_07349_),
    .A(net5796),
    .B(net5105));
 sg13g2_o21ai_1 _24956_ (.B1(_07349_),
    .Y(_07350_),
    .A1(net7130),
    .A2(net5105));
 sg13g2_nor2_1 _24957_ (.A(net6528),
    .B(_07350_),
    .Y(_01323_));
 sg13g2_nand2_1 _24958_ (.Y(_07351_),
    .A(net5776),
    .B(net5106));
 sg13g2_o21ai_1 _24959_ (.B1(_07351_),
    .Y(_07352_),
    .A1(net7291),
    .A2(net5106));
 sg13g2_nor2_1 _24960_ (.A(net6528),
    .B(_07352_),
    .Y(_01324_));
 sg13g2_nor2_1 _24961_ (.A(net5257),
    .B(_07321_),
    .Y(_07353_));
 sg13g2_nor2_1 _24962_ (.A(net4474),
    .B(net5041),
    .Y(_07354_));
 sg13g2_a21oi_1 _24963_ (.A1(net5759),
    .A2(net5041),
    .Y(_01325_),
    .B1(_07354_));
 sg13g2_nor2_1 _24964_ (.A(net4081),
    .B(net5041),
    .Y(_07355_));
 sg13g2_a21oi_1 _24965_ (.A1(net5781),
    .A2(net5041),
    .Y(_01326_),
    .B1(_07355_));
 sg13g2_nor2_1 _24966_ (.A(net3307),
    .B(net5042),
    .Y(_07356_));
 sg13g2_a21oi_1 _24967_ (.A1(net5710),
    .A2(net5042),
    .Y(_01327_),
    .B1(_07356_));
 sg13g2_nor2_1 _24968_ (.A(net3826),
    .B(_07353_),
    .Y(_07357_));
 sg13g2_a21oi_1 _24969_ (.A1(net5687),
    .A2(net5042),
    .Y(_01328_),
    .B1(_07357_));
 sg13g2_nor2_1 _24970_ (.A(net3400),
    .B(net5042),
    .Y(_07358_));
 sg13g2_a21oi_1 _24971_ (.A1(net5670),
    .A2(net5042),
    .Y(_01329_),
    .B1(_07358_));
 sg13g2_nor2_1 _24972_ (.A(net3878),
    .B(net5041),
    .Y(_07359_));
 sg13g2_a21oi_1 _24973_ (.A1(net5585),
    .A2(net5041),
    .Y(_01330_),
    .B1(_07359_));
 sg13g2_nor2_1 _24974_ (.A(net3109),
    .B(net5042),
    .Y(_07360_));
 sg13g2_a21oi_1 _24975_ (.A1(net5647),
    .A2(net5042),
    .Y(_01331_),
    .B1(_07360_));
 sg13g2_nor2_1 _24976_ (.A(net3415),
    .B(net5041),
    .Y(_07361_));
 sg13g2_a21oi_1 _24977_ (.A1(net5622),
    .A2(net5041),
    .Y(_01332_),
    .B1(_07361_));
 sg13g2_nor2_1 _24978_ (.A(_09441_),
    .B(_04767_),
    .Y(_07362_));
 sg13g2_nor2_1 _24979_ (.A(net3204),
    .B(net5039),
    .Y(_07363_));
 sg13g2_a21oi_1 _24980_ (.A1(net5768),
    .A2(net5039),
    .Y(_01333_),
    .B1(_07363_));
 sg13g2_nor2_1 _24981_ (.A(net3929),
    .B(net5040),
    .Y(_07364_));
 sg13g2_a21oi_1 _24982_ (.A1(net5788),
    .A2(net5040),
    .Y(_01334_),
    .B1(_07364_));
 sg13g2_nor2_1 _24983_ (.A(net3753),
    .B(net5040),
    .Y(_07365_));
 sg13g2_a21oi_1 _24984_ (.A1(net5718),
    .A2(_07362_),
    .Y(_01335_),
    .B1(_07365_));
 sg13g2_nor2_1 _24985_ (.A(net4339),
    .B(net5039),
    .Y(_07366_));
 sg13g2_a21oi_1 _24986_ (.A1(net5695),
    .A2(net5039),
    .Y(_01336_),
    .B1(_07366_));
 sg13g2_nor2_1 _24987_ (.A(net3341),
    .B(net5040),
    .Y(_07367_));
 sg13g2_a21oi_1 _24988_ (.A1(net5674),
    .A2(net5040),
    .Y(_01337_),
    .B1(_07367_));
 sg13g2_nor2_1 _24989_ (.A(net3669),
    .B(net5040),
    .Y(_07368_));
 sg13g2_a21oi_1 _24990_ (.A1(net5593),
    .A2(net5040),
    .Y(_01338_),
    .B1(_07368_));
 sg13g2_nor2_1 _24991_ (.A(net3270),
    .B(net5039),
    .Y(_07369_));
 sg13g2_a21oi_1 _24992_ (.A1(net5657),
    .A2(net5039),
    .Y(_01339_),
    .B1(_07369_));
 sg13g2_nor2_1 _24993_ (.A(net3538),
    .B(net5039),
    .Y(_07370_));
 sg13g2_a21oi_1 _24994_ (.A1(net5635),
    .A2(net5039),
    .Y(_01340_),
    .B1(_07370_));
 sg13g2_nor2_2 _24995_ (.A(net5514),
    .B(_03023_),
    .Y(_07371_));
 sg13g2_nor2_2 _24996_ (.A(net5273),
    .B(_07371_),
    .Y(_07372_));
 sg13g2_nand2_1 _24997_ (.Y(_07373_),
    .A(\atari2600.ram_data[0] ),
    .B(net5534));
 sg13g2_nand4_1 _24998_ (.B(\flash_rom.addr_in[17] ),
    .C(\flash_rom.addr_in[18] ),
    .A(\flash_rom.addr_in[16] ),
    .Y(_07374_),
    .D(\flash_rom.addr_in[19] ));
 sg13g2_nand2b_1 _24999_ (.Y(_07375_),
    .B(net6040),
    .A_N(\external_rom_data[0] ));
 sg13g2_o21ai_1 _25000_ (.B1(_07375_),
    .Y(_07376_),
    .A1(\internal_rom_data[0] ),
    .A2(net6040));
 sg13g2_o21ai_1 _25001_ (.B1(_07373_),
    .Y(_07377_),
    .A1(net5534),
    .A2(_07376_));
 sg13g2_a22oi_1 _25002_ (.Y(_07378_),
    .B1(_07372_),
    .B2(_07377_),
    .A2(net5273),
    .A1(net7327));
 sg13g2_inv_1 _25003_ (.Y(_01341_),
    .A(net7328));
 sg13g2_nand2_1 _25004_ (.Y(_07379_),
    .A(net7366),
    .B(net5535));
 sg13g2_nand2b_1 _25005_ (.Y(_07380_),
    .B(net6040),
    .A_N(\external_rom_data[1] ));
 sg13g2_o21ai_1 _25006_ (.B1(_07380_),
    .Y(_07381_),
    .A1(\internal_rom_data[1] ),
    .A2(net6041));
 sg13g2_o21ai_1 _25007_ (.B1(_07379_),
    .Y(_07382_),
    .A1(net5534),
    .A2(_07381_));
 sg13g2_a22oi_1 _25008_ (.Y(_07383_),
    .B1(_07372_),
    .B2(net7367),
    .A2(net5273),
    .A1(net4492));
 sg13g2_inv_1 _25009_ (.Y(_01342_),
    .A(_07383_));
 sg13g2_nand2_1 _25010_ (.Y(_07384_),
    .A(net7346),
    .B(net5535));
 sg13g2_nand2b_1 _25011_ (.Y(_07385_),
    .B(net6041),
    .A_N(\external_rom_data[2] ));
 sg13g2_o21ai_1 _25012_ (.B1(_07385_),
    .Y(_07386_),
    .A1(\internal_rom_data[2] ),
    .A2(net6041));
 sg13g2_o21ai_1 _25013_ (.B1(_07384_),
    .Y(_07387_),
    .A1(net5535),
    .A2(_07386_));
 sg13g2_a22oi_1 _25014_ (.Y(_07388_),
    .B1(_07372_),
    .B2(net7347),
    .A2(net5273),
    .A1(net4643));
 sg13g2_inv_2 _25015_ (.Y(_01343_),
    .A(_07388_));
 sg13g2_nand2_1 _25016_ (.Y(_07389_),
    .A(net7340),
    .B(net5534));
 sg13g2_nand2b_1 _25017_ (.Y(_07390_),
    .B(net6041),
    .A_N(\external_rom_data[3] ));
 sg13g2_o21ai_1 _25018_ (.B1(_07390_),
    .Y(_07391_),
    .A1(\internal_rom_data[3] ),
    .A2(net6040));
 sg13g2_o21ai_1 _25019_ (.B1(_07389_),
    .Y(_07392_),
    .A1(net5535),
    .A2(_07391_));
 sg13g2_a22oi_1 _25020_ (.Y(_07393_),
    .B1(_07372_),
    .B2(_07392_),
    .A2(net5273),
    .A1(net7128));
 sg13g2_inv_1 _25021_ (.Y(_01344_),
    .A(_07393_));
 sg13g2_nand2_1 _25022_ (.Y(_07394_),
    .A(net7269),
    .B(net5534));
 sg13g2_nand2b_1 _25023_ (.Y(_07395_),
    .B(net6040),
    .A_N(\external_rom_data[4] ));
 sg13g2_o21ai_1 _25024_ (.B1(_07395_),
    .Y(_07396_),
    .A1(\internal_rom_data[4] ),
    .A2(net6040));
 sg13g2_o21ai_1 _25025_ (.B1(_07394_),
    .Y(_07397_),
    .A1(net5534),
    .A2(_07396_));
 sg13g2_a22oi_1 _25026_ (.Y(_07398_),
    .B1(_07372_),
    .B2(_07397_),
    .A2(net5273),
    .A1(net7167));
 sg13g2_inv_1 _25027_ (.Y(_01345_),
    .A(_07398_));
 sg13g2_nand2_1 _25028_ (.Y(_07399_),
    .A(net7259),
    .B(net5534));
 sg13g2_nand2b_1 _25029_ (.Y(_07400_),
    .B(net6040),
    .A_N(\external_rom_data[5] ));
 sg13g2_o21ai_1 _25030_ (.B1(_07400_),
    .Y(_07401_),
    .A1(\internal_rom_data[5] ),
    .A2(net6040));
 sg13g2_o21ai_1 _25031_ (.B1(_07399_),
    .Y(_07402_),
    .A1(net5534),
    .A2(_07401_));
 sg13g2_a22oi_1 _25032_ (.Y(_07403_),
    .B1(_07372_),
    .B2(net7260),
    .A2(net5273),
    .A1(net7157));
 sg13g2_inv_1 _25033_ (.Y(_01346_),
    .A(_07403_));
 sg13g2_mux2_1 _25034_ (.A0(\internal_rom_data[6] ),
    .A1(\external_rom_data[6] ),
    .S(net6041),
    .X(_07404_));
 sg13g2_a22oi_1 _25035_ (.Y(_07405_),
    .B1(_07371_),
    .B2(net4423),
    .A2(_03025_),
    .A1(\atari2600.ram_data[6] ));
 sg13g2_a22oi_1 _25036_ (.Y(_07406_),
    .B1(_07404_),
    .B2(_03023_),
    .A2(net5274),
    .A1(net4459));
 sg13g2_o21ai_1 _25037_ (.B1(_07406_),
    .Y(_01347_),
    .A1(net5274),
    .A2(_07405_));
 sg13g2_mux2_1 _25038_ (.A0(\internal_rom_data[7] ),
    .A1(net4380),
    .S(net6041),
    .X(_07407_));
 sg13g2_a22oi_1 _25039_ (.Y(_07408_),
    .B1(_07371_),
    .B2(net4341),
    .A2(_03025_),
    .A1(net7473));
 sg13g2_a22oi_1 _25040_ (.Y(_07409_),
    .B1(_07407_),
    .B2(_03023_),
    .A2(net5274),
    .A1(net4779));
 sg13g2_o21ai_1 _25041_ (.B1(_07409_),
    .Y(_01348_),
    .A1(net5274),
    .A2(_07408_));
 sg13g2_nor2_1 _25042_ (.A(net7065),
    .B(net5833),
    .Y(_07410_));
 sg13g2_a21oi_1 _25043_ (.A1(net5833),
    .A2(_08762_),
    .Y(_01349_),
    .B1(_07410_));
 sg13g2_nor2_1 _25044_ (.A(net7395),
    .B(net5833),
    .Y(_07411_));
 sg13g2_a21oi_1 _25045_ (.A1(net5833),
    .A2(_08757_),
    .Y(_01350_),
    .B1(_07411_));
 sg13g2_nor2_1 _25046_ (.A(net7292),
    .B(net5833),
    .Y(_07412_));
 sg13g2_a21oi_1 _25047_ (.A1(net5833),
    .A2(net5736),
    .Y(_01351_),
    .B1(_07412_));
 sg13g2_a22oi_1 _25048_ (.Y(_07413_),
    .B1(_08888_),
    .B2(_08896_),
    .A2(net5817),
    .A1(net6257));
 sg13g2_inv_1 _25049_ (.Y(_01352_),
    .A(_07413_));
 sg13g2_nand2_1 _25050_ (.Y(_07414_),
    .A(net7454),
    .B(net5817));
 sg13g2_o21ai_1 _25051_ (.B1(_07414_),
    .Y(_01353_),
    .A1(_08756_),
    .A2(_08954_));
 sg13g2_nor3_1 _25052_ (.A(_08746_),
    .B(_08756_),
    .C(net5818),
    .Y(_07415_));
 sg13g2_nand4_1 _25053_ (.B(net5732),
    .C(_08886_),
    .A(net5735),
    .Y(_07416_),
    .D(_07415_));
 sg13g2_o21ai_1 _25054_ (.B1(_07416_),
    .Y(_01354_),
    .A1(_08635_),
    .A2(net5824));
 sg13g2_nor2_1 _25055_ (.A(net5733),
    .B(net5732),
    .Y(_07417_));
 sg13g2_nand3_1 _25056_ (.B(_07415_),
    .C(_07417_),
    .A(_08886_),
    .Y(_07418_));
 sg13g2_o21ai_1 _25057_ (.B1(_07418_),
    .Y(_01355_),
    .A1(_08636_),
    .A2(net5822));
 sg13g2_nand2_1 _25058_ (.Y(_07419_),
    .A(net5732),
    .B(_08935_));
 sg13g2_nor2_2 _25059_ (.A(_08747_),
    .B(_08757_),
    .Y(_07420_));
 sg13g2_nand2_1 _25060_ (.Y(_07421_),
    .A(_08886_),
    .B(_07420_));
 sg13g2_nand2_1 _25061_ (.Y(_07422_),
    .A(net3246),
    .B(net5817));
 sg13g2_o21ai_1 _25062_ (.B1(_07422_),
    .Y(_01356_),
    .A1(_07419_),
    .A2(_07421_));
 sg13g2_nand2_1 _25063_ (.Y(_07423_),
    .A(net3208),
    .B(net5817));
 sg13g2_nand2_1 _25064_ (.Y(_07424_),
    .A(net5822),
    .B(_07417_));
 sg13g2_o21ai_1 _25065_ (.B1(_07423_),
    .Y(_01357_),
    .A1(_07421_),
    .A2(_07424_));
 sg13g2_nand3_1 _25066_ (.B(_08756_),
    .C(_08886_),
    .A(_08747_),
    .Y(_07425_));
 sg13g2_nand2_1 _25067_ (.Y(_07426_),
    .A(net3007),
    .B(net5817));
 sg13g2_o21ai_1 _25068_ (.B1(_07426_),
    .Y(_01358_),
    .A1(_07419_),
    .A2(_07425_));
 sg13g2_nand2_1 _25069_ (.Y(_07427_),
    .A(net3546),
    .B(net5817));
 sg13g2_o21ai_1 _25070_ (.B1(_07427_),
    .Y(_01359_),
    .A1(_07424_),
    .A2(_07425_));
 sg13g2_nor2_2 _25071_ (.A(net5736),
    .B(_08756_),
    .Y(_07428_));
 sg13g2_nor3_2 _25072_ (.A(net5736),
    .B(_08756_),
    .C(net5731),
    .Y(_07429_));
 sg13g2_nand3_1 _25073_ (.B(_08888_),
    .C(_07429_),
    .A(net5735),
    .Y(_07430_));
 sg13g2_o21ai_1 _25074_ (.B1(_07430_),
    .Y(_01360_),
    .A1(_08638_),
    .A2(net5824));
 sg13g2_nor2_1 _25075_ (.A(net7164),
    .B(net5824),
    .Y(_07431_));
 sg13g2_a21oi_1 _25076_ (.A1(net5824),
    .A2(_09004_),
    .Y(_01361_),
    .B1(_07431_));
 sg13g2_nand2_1 _25077_ (.Y(_07432_),
    .A(net7296),
    .B(net5818));
 sg13g2_nand4_1 _25078_ (.B(net5822),
    .C(_08836_),
    .A(net5736),
    .Y(_07433_),
    .D(_08989_));
 sg13g2_o21ai_1 _25079_ (.B1(_07432_),
    .Y(_01362_),
    .A1(net5732),
    .A2(_07433_));
 sg13g2_a21oi_2 _25080_ (.B1(net5820),
    .Y(_07434_),
    .A2(_08989_),
    .A1(net5736));
 sg13g2_o21ai_1 _25081_ (.B1(net5822),
    .Y(_07435_),
    .A1(_08746_),
    .A2(_08990_));
 sg13g2_o21ai_1 _25082_ (.B1(_07435_),
    .Y(_07436_),
    .A1(_08756_),
    .A2(net5819));
 sg13g2_a21oi_1 _25083_ (.A1(_08587_),
    .A2(net5819),
    .Y(_01363_),
    .B1(_07436_));
 sg13g2_nand2_1 _25084_ (.Y(_07437_),
    .A(net5734),
    .B(_07420_));
 sg13g2_inv_1 _25085_ (.Y(_07438_),
    .A(_07437_));
 sg13g2_nand3_1 _25086_ (.B(net5730),
    .C(_07438_),
    .A(_08739_),
    .Y(_07439_));
 sg13g2_nand2_1 _25087_ (.Y(_07440_),
    .A(_08830_),
    .B(_07420_));
 sg13g2_nand3_1 _25088_ (.B(_08830_),
    .C(_07420_),
    .A(net5731),
    .Y(_07441_));
 sg13g2_nand3_1 _25089_ (.B(_07439_),
    .C(_07441_),
    .A(net5823),
    .Y(_07442_));
 sg13g2_o21ai_1 _25090_ (.B1(_07442_),
    .Y(_07443_),
    .A1(net7446),
    .A2(net5824));
 sg13g2_inv_1 _25091_ (.Y(_01364_),
    .A(_07443_));
 sg13g2_o21ai_1 _25092_ (.B1(net5856),
    .Y(_07444_),
    .A1(net6034),
    .A2(_08872_));
 sg13g2_nand2_1 _25093_ (.Y(_07445_),
    .A(net7161),
    .B(_07444_));
 sg13g2_nand2_1 _25094_ (.Y(_07446_),
    .A(net4937),
    .B(net5736));
 sg13g2_nand3b_1 _25095_ (.B(_08830_),
    .C(_08763_),
    .Y(_07447_),
    .A_N(_07444_));
 sg13g2_o21ai_1 _25096_ (.B1(_07445_),
    .Y(_01365_),
    .A1(_07446_),
    .A2(_07447_));
 sg13g2_o21ai_1 _25097_ (.B1(_07433_),
    .Y(_01366_),
    .A1(_08590_),
    .A2(net5822));
 sg13g2_nand2_1 _25098_ (.Y(_07448_),
    .A(net7170),
    .B(_07444_));
 sg13g2_nand2_1 _25099_ (.Y(_01367_),
    .A(_07447_),
    .B(_07448_));
 sg13g2_a22oi_1 _25100_ (.Y(_07449_),
    .B1(_08888_),
    .B2(_07438_),
    .A2(net5818),
    .A1(net7280));
 sg13g2_nand3_1 _25101_ (.B(net5822),
    .C(_08989_),
    .A(net5755),
    .Y(_07450_));
 sg13g2_nand2_1 _25102_ (.Y(_07451_),
    .A(_08761_),
    .B(_07420_));
 sg13g2_o21ai_1 _25103_ (.B1(_07449_),
    .Y(_01368_),
    .A1(_07450_),
    .A2(_07451_));
 sg13g2_mux2_1 _25104_ (.A0(net7290),
    .A1(_07429_),
    .S(net5824),
    .X(_01369_));
 sg13g2_nand2_1 _25105_ (.Y(_07452_),
    .A(net3316),
    .B(net5817));
 sg13g2_o21ai_1 _25106_ (.B1(_07452_),
    .Y(_01370_),
    .A1(_07428_),
    .A2(_07450_));
 sg13g2_nand2_1 _25107_ (.Y(_07453_),
    .A(_08746_),
    .B(_08762_));
 sg13g2_nand2_2 _25108_ (.Y(_07454_),
    .A(net5731),
    .B(_07428_));
 sg13g2_a21oi_1 _25109_ (.A1(_08726_),
    .A2(_08733_),
    .Y(_07455_),
    .B1(_08830_));
 sg13g2_nor3_1 _25110_ (.A(net5820),
    .B(_07454_),
    .C(_07455_),
    .Y(_07456_));
 sg13g2_a21o_1 _25111_ (.A2(net5819),
    .A1(net7464),
    .B1(_07456_),
    .X(_01371_));
 sg13g2_and4_1 _25112_ (.A(net5755),
    .B(_08751_),
    .C(_08989_),
    .D(_07428_),
    .X(_07457_));
 sg13g2_nand2_1 _25113_ (.Y(_07458_),
    .A(net7102),
    .B(net5821));
 sg13g2_o21ai_1 _25114_ (.B1(net5823),
    .Y(_07459_),
    .A1(_08833_),
    .A2(_07457_));
 sg13g2_nand3_1 _25115_ (.B(_07458_),
    .C(_07459_),
    .A(_08936_),
    .Y(_01372_));
 sg13g2_o21ai_1 _25116_ (.B1(net6546),
    .Y(_01373_),
    .A1(_08490_),
    .A2(net5824));
 sg13g2_nand2_1 _25117_ (.Y(_07460_),
    .A(net5755),
    .B(_07428_));
 sg13g2_nand3_1 _25118_ (.B(net5735),
    .C(_07429_),
    .A(net5755),
    .Y(_07461_));
 sg13g2_o21ai_1 _25119_ (.B1(_07461_),
    .Y(_07462_),
    .A1(net5730),
    .A2(_07454_));
 sg13g2_nand2_1 _25120_ (.Y(_07463_),
    .A(net5754),
    .B(_07462_));
 sg13g2_nor3_1 _25121_ (.A(_08761_),
    .B(_08991_),
    .C(_07437_),
    .Y(_07464_));
 sg13g2_nand2b_1 _25122_ (.Y(_07465_),
    .B(net5822),
    .A_N(_07464_));
 sg13g2_nand2_1 _25123_ (.Y(_07466_),
    .A(_08989_),
    .B(_07429_));
 sg13g2_nor3_1 _25124_ (.A(net5734),
    .B(_08832_),
    .C(_07466_),
    .Y(_07467_));
 sg13g2_nand3_1 _25125_ (.B(net5734),
    .C(_07429_),
    .A(net5754),
    .Y(_07468_));
 sg13g2_a22oi_1 _25126_ (.Y(_07469_),
    .B1(_07453_),
    .B2(_08830_),
    .A2(_08992_),
    .A1(_08753_));
 sg13g2_nand3_1 _25127_ (.B(_07468_),
    .C(_07469_),
    .A(_09018_),
    .Y(_07470_));
 sg13g2_nor3_1 _25128_ (.A(_07465_),
    .B(_07467_),
    .C(_07470_),
    .Y(_07471_));
 sg13g2_nor2_1 _25129_ (.A(net5819),
    .B(_07467_),
    .Y(_07472_));
 sg13g2_a22oi_1 _25130_ (.Y(_01374_),
    .B1(_07463_),
    .B2(_07471_),
    .A2(net5820),
    .A1(_08639_));
 sg13g2_and2_1 _25131_ (.A(net6256),
    .B(net6544),
    .X(_07473_));
 sg13g2_nor3_1 _25132_ (.A(net6522),
    .B(net5862),
    .C(_04868_),
    .Y(_07474_));
 sg13g2_a21o_1 _25133_ (.A2(_07473_),
    .A1(net5821),
    .B1(net5801),
    .X(_01375_));
 sg13g2_nor2_1 _25134_ (.A(net4640),
    .B(net5802),
    .Y(_07475_));
 sg13g2_a21oi_1 _25135_ (.A1(_08731_),
    .A2(net5802),
    .Y(_01376_),
    .B1(_07475_));
 sg13g2_mux2_1 _25136_ (.A0(net7266),
    .A1(\atari2600.cpu.DIMUX[1] ),
    .S(net5801),
    .X(_01377_));
 sg13g2_mux2_1 _25137_ (.A0(net7181),
    .A1(\atari2600.cpu.DIMUX[2] ),
    .S(net5802),
    .X(_01378_));
 sg13g2_mux2_1 _25138_ (.A0(net7187),
    .A1(\atari2600.cpu.DIMUX[3] ),
    .S(net5801),
    .X(_01379_));
 sg13g2_nor2_1 _25139_ (.A(net4471),
    .B(net5801),
    .Y(_07476_));
 sg13g2_a21oi_1 _25140_ (.A1(_08749_),
    .A2(net5801),
    .Y(_01380_),
    .B1(_07476_));
 sg13g2_nor2_1 _25141_ (.A(net7036),
    .B(net5801),
    .Y(_07477_));
 sg13g2_a21oi_1 _25142_ (.A1(_08759_),
    .A2(net5801),
    .Y(_01381_),
    .B1(_07477_));
 sg13g2_mux2_1 _25143_ (.A0(net7250),
    .A1(\atari2600.cpu.DIMUX[6] ),
    .S(net5801),
    .X(_01382_));
 sg13g2_nor2_1 _25144_ (.A(net7217),
    .B(net5802),
    .Y(_07478_));
 sg13g2_a21oi_1 _25145_ (.A1(_08744_),
    .A2(net5802),
    .Y(_01383_),
    .B1(_07478_));
 sg13g2_nor2_1 _25146_ (.A(net6034),
    .B(net5998),
    .Y(_07479_));
 sg13g2_inv_1 _25147_ (.Y(_07480_),
    .A(_07479_));
 sg13g2_nor2_1 _25148_ (.A(\atari2600.cpu.cld ),
    .B(\atari2600.cpu.sed ),
    .Y(_07481_));
 sg13g2_a21oi_1 _25149_ (.A1(_05126_),
    .A2(_07481_),
    .Y(_07482_),
    .B1(_07479_));
 sg13g2_nor2b_1 _25150_ (.A(net6257),
    .B_N(_00164_),
    .Y(_07483_));
 sg13g2_a21oi_1 _25151_ (.A1(\atari2600.cpu.ADD[3] ),
    .A2(net6257),
    .Y(_07484_),
    .B1(_07483_));
 sg13g2_o21ai_1 _25152_ (.B1(_07482_),
    .Y(_07485_),
    .A1(net5998),
    .A2(_07484_));
 sg13g2_a21oi_1 _25153_ (.A1(net5826),
    .A2(net5998),
    .Y(_07486_),
    .B1(_07485_));
 sg13g2_nor2_1 _25154_ (.A(\atari2600.cpu.D ),
    .B(_07482_),
    .Y(_07487_));
 sg13g2_nor4_1 _25155_ (.A(net2946),
    .B(net6524),
    .C(_07486_),
    .D(_07487_),
    .Y(_01384_));
 sg13g2_nor2b_1 _25156_ (.A(net5827),
    .B_N(net5999),
    .Y(_07488_));
 sg13g2_nor3_1 _25157_ (.A(\atari2600.cpu.sei ),
    .B(\atari2600.cpu.cli ),
    .C(_08804_),
    .Y(_07489_));
 sg13g2_a221oi_1 _25158_ (.B2(_07479_),
    .C1(_07489_),
    .B1(_08995_),
    .A1(net6518),
    .Y(_07490_),
    .A2(_00134_));
 sg13g2_nand2_1 _25159_ (.Y(_07491_),
    .A(_00165_),
    .B(_08994_));
 sg13g2_a21oi_1 _25160_ (.A1(\atari2600.cpu.ADD[2] ),
    .A2(_08995_),
    .Y(_07492_),
    .B1(net5998));
 sg13g2_a21oi_1 _25161_ (.A1(_07491_),
    .A2(_07492_),
    .Y(_07493_),
    .B1(_07488_));
 sg13g2_nand2_1 _25162_ (.Y(_07494_),
    .A(_07490_),
    .B(_07493_));
 sg13g2_nand2b_1 _25163_ (.Y(_07495_),
    .B(net7191),
    .A_N(_07490_));
 sg13g2_nand3_1 _25164_ (.B(_07494_),
    .C(_07495_),
    .A(_08847_),
    .Y(_01385_));
 sg13g2_a21oi_1 _25165_ (.A1(\atari2600.cpu.bit_ins ),
    .A2(_08795_),
    .Y(_07496_),
    .B1(_07480_));
 sg13g2_nor3_1 _25166_ (.A(net6257),
    .B(\atari2600.cpu.clv ),
    .C(_08771_),
    .Y(_07497_));
 sg13g2_a21oi_1 _25167_ (.A1(_08637_),
    .A2(_07497_),
    .Y(_07498_),
    .B1(_07496_));
 sg13g2_nand3_1 _25168_ (.B(net6257),
    .C(net6034),
    .A(\atari2600.cpu.ADD[6] ),
    .Y(_07499_));
 sg13g2_xor2_1 _25169_ (.B(\atari2600.cpu.ALU.AI7 ),
    .A(\atari2600.cpu.ALU.BI7 ),
    .X(_07500_));
 sg13g2_xor2_1 _25170_ (.B(_00091_),
    .A(net6247),
    .X(_07501_));
 sg13g2_xnor2_1 _25171_ (.Y(_07502_),
    .A(_07500_),
    .B(_07501_));
 sg13g2_a22oi_1 _25172_ (.Y(_07503_),
    .B1(_07497_),
    .B2(_07502_),
    .A2(_08771_),
    .A1(net5825));
 sg13g2_nand2_1 _25173_ (.Y(_07504_),
    .A(_07499_),
    .B(_07503_));
 sg13g2_mux2_1 _25174_ (.A0(net7218),
    .A1(_07504_),
    .S(_07498_),
    .X(_01386_));
 sg13g2_o21ai_1 _25175_ (.B1(_05126_),
    .Y(_07505_),
    .A1(_08639_),
    .A2(_09062_));
 sg13g2_nor2_1 _25176_ (.A(\atari2600.cpu.compare ),
    .B(_07505_),
    .Y(_07506_));
 sg13g2_a21oi_1 _25177_ (.A1(_08815_),
    .A2(_07496_),
    .Y(_07507_),
    .B1(_07506_));
 sg13g2_nor2_1 _25178_ (.A(net6034),
    .B(_08814_),
    .Y(_07508_));
 sg13g2_mux2_1 _25179_ (.A0(\atari2600.cpu.ADD[7] ),
    .A1(\atari2600.cpu.DIMUX[7] ),
    .S(_07508_),
    .X(_07509_));
 sg13g2_mux2_1 _25180_ (.A0(net4176),
    .A1(_07509_),
    .S(_07507_),
    .X(_01387_));
 sg13g2_nor4_1 _25181_ (.A(net6248),
    .B(\atari2600.cpu.ADD[7] ),
    .C(\atari2600.cpu.ADD[5] ),
    .D(net6250),
    .Y(_07510_));
 sg13g2_nor4_1 _25182_ (.A(\atari2600.cpu.ADD[1] ),
    .B(net6251),
    .C(net6253),
    .D(\atari2600.cpu.ADD[3] ),
    .Y(_07511_));
 sg13g2_nand2_1 _25183_ (.Y(_07512_),
    .A(_07510_),
    .B(_07511_));
 sg13g2_or2_1 _25184_ (.X(_07513_),
    .B(_07512_),
    .A(net6257));
 sg13g2_a21oi_1 _25185_ (.A1(net6252),
    .A2(net6257),
    .Y(_07514_),
    .B1(net5998));
 sg13g2_a221oi_1 _25186_ (.B2(_07514_),
    .C1(_08814_),
    .B1(_07513_),
    .A1(_08735_),
    .Y(_07515_),
    .A2(net5998));
 sg13g2_nor2_1 _25187_ (.A(_08815_),
    .B(_07512_),
    .Y(_07516_));
 sg13g2_nand2b_1 _25188_ (.Y(_07517_),
    .B(_07506_),
    .A_N(\atari2600.cpu.bit_ins ));
 sg13g2_o21ai_1 _25189_ (.B1(_07517_),
    .Y(_07518_),
    .A1(_08814_),
    .A2(_07480_));
 sg13g2_nor3_1 _25190_ (.A(_07515_),
    .B(_07516_),
    .C(_07518_),
    .Y(_07519_));
 sg13g2_a21oi_1 _25191_ (.A1(_08578_),
    .A2(_07518_),
    .Y(_01388_),
    .B1(_07519_));
 sg13g2_a22oi_1 _25192_ (.Y(_07520_),
    .B1(_08814_),
    .B2(\atari2600.cpu.shift ),
    .A2(net6034),
    .A1(_00133_));
 sg13g2_nor3_1 _25193_ (.A(\atari2600.cpu.shift ),
    .B(\atari2600.cpu.compare ),
    .C(\atari2600.cpu.adc_sbc ),
    .Y(_07521_));
 sg13g2_nor3_1 _25194_ (.A(\atari2600.cpu.clc ),
    .B(\atari2600.cpu.plp ),
    .C(\atari2600.cpu.sec ),
    .Y(_07522_));
 sg13g2_a21oi_1 _25195_ (.A1(_07521_),
    .A2(_07522_),
    .Y(_07523_),
    .B1(_07520_));
 sg13g2_nor2b_1 _25196_ (.A(\atari2600.cpu.plp ),
    .B_N(_00166_),
    .Y(_07524_));
 sg13g2_a21oi_1 _25197_ (.A1(net6253),
    .A2(\atari2600.cpu.plp ),
    .Y(_07525_),
    .B1(_07524_));
 sg13g2_nor2_1 _25198_ (.A(net6247),
    .B(_07521_),
    .Y(_07526_));
 sg13g2_a21oi_1 _25199_ (.A1(_07521_),
    .A2(_07525_),
    .Y(_07527_),
    .B1(_07526_));
 sg13g2_nand2_1 _25200_ (.Y(_07528_),
    .A(_07523_),
    .B(_07527_));
 sg13g2_o21ai_1 _25201_ (.B1(_07528_),
    .Y(_07529_),
    .A1(_08582_),
    .A2(_07523_));
 sg13g2_nor2_1 _25202_ (.A(net5998),
    .B(_07529_),
    .Y(_07530_));
 sg13g2_a21oi_1 _25203_ (.A1(net7517),
    .A2(net5998),
    .Y(_01389_),
    .B1(_07530_));
 sg13g2_mux2_1 _25204_ (.A0(net7143),
    .A1(\atari2600.cpu.backwards ),
    .S(net5866),
    .X(_01390_));
 sg13g2_mux2_1 _25205_ (.A0(_09152_),
    .A1(net7096),
    .S(net5815),
    .X(_01391_));
 sg13g2_mux2_1 _25206_ (.A0(_09134_),
    .A1(net7248),
    .S(net5815),
    .X(_01392_));
 sg13g2_mux2_1 _25207_ (.A0(_09144_),
    .A1(net7003),
    .S(net5813),
    .X(_01393_));
 sg13g2_mux2_1 _25208_ (.A0(_09164_),
    .A1(net7059),
    .S(net5813),
    .X(_01394_));
 sg13g2_mux2_1 _25209_ (.A0(_09091_),
    .A1(net7150),
    .S(net5813),
    .X(_01395_));
 sg13g2_mux2_1 _25210_ (.A0(_09103_),
    .A1(net7115),
    .S(net5813),
    .X(_01396_));
 sg13g2_mux2_1 _25211_ (.A0(_09258_),
    .A1(net7183),
    .S(net5814),
    .X(_01397_));
 sg13g2_nand2_1 _25212_ (.Y(_07531_),
    .A(net3521),
    .B(net5813));
 sg13g2_o21ai_1 _25213_ (.B1(_07531_),
    .Y(_01398_),
    .A1(_09121_),
    .A2(net5813));
 sg13g2_mux2_1 _25214_ (.A0(net4482),
    .A1(_05271_),
    .S(net5828),
    .X(_01399_));
 sg13g2_nor2_1 _25215_ (.A(net6253),
    .B(net5855),
    .Y(_07532_));
 sg13g2_nor2_1 _25216_ (.A(_05236_),
    .B(net5916),
    .Y(_07533_));
 sg13g2_nor3_1 _25217_ (.A(net5934),
    .B(_05259_),
    .C(_07533_),
    .Y(_07534_));
 sg13g2_nand2_1 _25218_ (.Y(_07535_),
    .A(\atari2600.cpu.PC[0] ),
    .B(net5991));
 sg13g2_o21ai_1 _25219_ (.B1(_07535_),
    .Y(_07536_),
    .A1(_08731_),
    .A2(_05244_));
 sg13g2_xnor2_1 _25220_ (.Y(_07537_),
    .A(net5916),
    .B(_07536_));
 sg13g2_nand2_1 _25221_ (.Y(_07538_),
    .A(net5917),
    .B(_07537_));
 sg13g2_a22oi_1 _25222_ (.Y(_07539_),
    .B1(net5928),
    .B2(net6252),
    .A2(net5995),
    .A1(\atari2600.cpu.ABH[1] ));
 sg13g2_a22oi_1 _25223_ (.Y(_07540_),
    .B1(_05268_),
    .B2(_09129_),
    .A2(_05237_),
    .A1(\atari2600.cpu.DIMUX[1] ));
 sg13g2_nand2_2 _25224_ (.Y(_07541_),
    .A(_07539_),
    .B(_07540_));
 sg13g2_a22oi_1 _25225_ (.Y(_07542_),
    .B1(_09072_),
    .B2(net6253),
    .A2(net5995),
    .A1(\atari2600.cpu.ABH[0] ));
 sg13g2_o21ai_1 _25226_ (.B1(_07542_),
    .Y(_07543_),
    .A1(_08731_),
    .A2(_05238_));
 sg13g2_a21o_1 _25227_ (.A2(_05268_),
    .A1(_09148_),
    .B1(_07543_),
    .X(_07544_));
 sg13g2_nand3_1 _25228_ (.B(_07536_),
    .C(_07544_),
    .A(_05265_),
    .Y(_07545_));
 sg13g2_and2_1 _25229_ (.A(_05263_),
    .B(_07536_),
    .X(_07546_));
 sg13g2_a21o_1 _25230_ (.A2(_07545_),
    .A1(_05266_),
    .B1(_07546_),
    .X(_07547_));
 sg13g2_a21oi_1 _25231_ (.A1(_05265_),
    .A2(_07536_),
    .Y(_07548_),
    .B1(_07544_));
 sg13g2_nor2_1 _25232_ (.A(_05250_),
    .B(_07548_),
    .Y(_07549_));
 sg13g2_a22oi_1 _25233_ (.Y(_07550_),
    .B1(_07547_),
    .B2(_07549_),
    .A2(_07541_),
    .A1(_05250_));
 sg13g2_a21oi_1 _25234_ (.A1(_05278_),
    .A2(_07538_),
    .Y(_07551_),
    .B1(_07550_));
 sg13g2_nand2_1 _25235_ (.Y(_07552_),
    .A(_07538_),
    .B(_07550_));
 sg13g2_nand2b_1 _25236_ (.Y(_07553_),
    .B(_07552_),
    .A_N(_07551_));
 sg13g2_xor2_1 _25237_ (.B(_07553_),
    .A(_07534_),
    .X(_07554_));
 sg13g2_a21oi_1 _25238_ (.A1(net5829),
    .A2(_07554_),
    .Y(_01400_),
    .B1(_07532_));
 sg13g2_nor2_1 _25239_ (.A(net6252),
    .B(net5854),
    .Y(_07555_));
 sg13g2_a21oi_1 _25240_ (.A1(_07534_),
    .A2(_07552_),
    .Y(_07556_),
    .B1(_07551_));
 sg13g2_nand2_1 _25241_ (.Y(_07557_),
    .A(\atari2600.cpu.PC[1] ),
    .B(net5991));
 sg13g2_o21ai_1 _25242_ (.B1(_07557_),
    .Y(_07558_),
    .A1(_08735_),
    .A2(_05244_));
 sg13g2_xnor2_1 _25243_ (.Y(_07559_),
    .A(net5916),
    .B(_07558_));
 sg13g2_and2_1 _25244_ (.A(net5917),
    .B(_07559_),
    .X(_07560_));
 sg13g2_a22oi_1 _25245_ (.Y(_07561_),
    .B1(net5928),
    .B2(net6251),
    .A2(net5994),
    .A1(\atari2600.cpu.ABH[2] ));
 sg13g2_a22oi_1 _25246_ (.Y(_07562_),
    .B1(_05268_),
    .B2(_09139_),
    .A2(_05237_),
    .A1(net5827));
 sg13g2_and2_1 _25247_ (.A(_07561_),
    .B(_07562_),
    .X(_07563_));
 sg13g2_inv_1 _25248_ (.Y(_07564_),
    .A(_07563_));
 sg13g2_a21oi_1 _25249_ (.A1(_05266_),
    .A2(_07541_),
    .Y(_07565_),
    .B1(_07558_));
 sg13g2_nor2_1 _25250_ (.A(_05265_),
    .B(_07541_),
    .Y(_07566_));
 sg13g2_and4_1 _25251_ (.A(_05262_),
    .B(net5875),
    .C(_07541_),
    .D(_07558_),
    .X(_07567_));
 sg13g2_nor4_1 _25252_ (.A(net5934),
    .B(_07565_),
    .C(_07566_),
    .D(_07567_),
    .Y(_07568_));
 sg13g2_a21oi_2 _25253_ (.B1(_07568_),
    .Y(_07569_),
    .A2(_07564_),
    .A1(net5934));
 sg13g2_nor2b_1 _25254_ (.A(_07560_),
    .B_N(_07569_),
    .Y(_07570_));
 sg13g2_nor2_1 _25255_ (.A(_05277_),
    .B(_07560_),
    .Y(_07571_));
 sg13g2_or2_1 _25256_ (.X(_07572_),
    .B(_07571_),
    .A(_07569_));
 sg13g2_mux2_1 _25257_ (.A0(_07571_),
    .A1(_07560_),
    .S(_07569_),
    .X(_07573_));
 sg13g2_xnor2_1 _25258_ (.Y(_07574_),
    .A(_07556_),
    .B(_07573_));
 sg13g2_inv_1 _25259_ (.Y(_07575_),
    .A(_07574_));
 sg13g2_a21oi_1 _25260_ (.A1(net5828),
    .A2(_07575_),
    .Y(_01401_),
    .B1(_07555_));
 sg13g2_nor2_1 _25261_ (.A(net6251),
    .B(net5854),
    .Y(_07576_));
 sg13g2_o21ai_1 _25262_ (.B1(_07572_),
    .Y(_07577_),
    .A1(_07556_),
    .A2(_07570_));
 sg13g2_a22oi_1 _25263_ (.Y(_07578_),
    .B1(net5928),
    .B2(\atari2600.cpu.ADD[3] ),
    .A2(net5996),
    .A1(\atari2600.cpu.ABH[3] ));
 sg13g2_a22oi_1 _25264_ (.Y(_07579_),
    .B1(_05268_),
    .B2(_09159_),
    .A2(_05237_),
    .A1(net5826));
 sg13g2_nand2_1 _25265_ (.Y(_07580_),
    .A(_07578_),
    .B(_07579_));
 sg13g2_a22oi_1 _25266_ (.Y(_07581_),
    .B1(_05243_),
    .B2(net5827),
    .A2(net5991),
    .A1(_08585_));
 sg13g2_nand2b_1 _25267_ (.Y(_07582_),
    .B(net5875),
    .A_N(_07581_));
 sg13g2_o21ai_1 _25268_ (.B1(_05266_),
    .Y(_07583_),
    .A1(_07563_),
    .A2(_07582_));
 sg13g2_o21ai_1 _25269_ (.B1(_07583_),
    .Y(_07584_),
    .A1(_05264_),
    .A2(_07581_));
 sg13g2_a21oi_1 _25270_ (.A1(_07563_),
    .A2(_07582_),
    .Y(_07585_),
    .B1(_05250_));
 sg13g2_a22oi_1 _25271_ (.Y(_07586_),
    .B1(_07584_),
    .B2(_07585_),
    .A2(_07580_),
    .A1(net5934));
 sg13g2_o21ai_1 _25272_ (.B1(_05236_),
    .Y(_07587_),
    .A1(net5916),
    .A2(_07581_));
 sg13g2_a21o_1 _25273_ (.A2(_07581_),
    .A1(net5916),
    .B1(_07587_),
    .X(_07588_));
 sg13g2_nand2_1 _25274_ (.Y(_07589_),
    .A(_05278_),
    .B(_07588_));
 sg13g2_nor2b_1 _25275_ (.A(_07586_),
    .B_N(_07589_),
    .Y(_07590_));
 sg13g2_nand2_1 _25276_ (.Y(_07591_),
    .A(_07586_),
    .B(_07588_));
 sg13g2_mux2_1 _25277_ (.A0(_07589_),
    .A1(_07588_),
    .S(_07586_),
    .X(_07592_));
 sg13g2_xor2_1 _25278_ (.B(_07592_),
    .A(_07577_),
    .X(_07593_));
 sg13g2_a21oi_1 _25279_ (.A1(net5828),
    .A2(_07593_),
    .Y(_01402_),
    .B1(_07576_));
 sg13g2_nor2_1 _25280_ (.A(net7480),
    .B(net5854),
    .Y(_07594_));
 sg13g2_a22oi_1 _25281_ (.Y(_07595_),
    .B1(net5928),
    .B2(net6250),
    .A2(net5993),
    .A1(\atari2600.cpu.ABH[4] ));
 sg13g2_a22oi_1 _25282_ (.Y(_07596_),
    .B1(_05268_),
    .B2(_09064_),
    .A2(_05237_),
    .A1(\atari2600.cpu.DIMUX[4] ));
 sg13g2_nand2_1 _25283_ (.Y(_07597_),
    .A(_07595_),
    .B(_07596_));
 sg13g2_inv_1 _25284_ (.Y(_07598_),
    .A(_07597_));
 sg13g2_a22oi_1 _25285_ (.Y(_07599_),
    .B1(_05243_),
    .B2(net5826),
    .A2(net5991),
    .A1(\atari2600.cpu.PC[3] ));
 sg13g2_inv_1 _25286_ (.Y(_07600_),
    .A(_07599_));
 sg13g2_nor2b_1 _25287_ (.A(_07599_),
    .B_N(net5875),
    .Y(_07601_));
 sg13g2_nand2_1 _25288_ (.Y(_07602_),
    .A(_07580_),
    .B(_07601_));
 sg13g2_a22oi_1 _25289_ (.Y(_07603_),
    .B1(_07602_),
    .B2(_05266_),
    .A2(_07600_),
    .A1(_05263_));
 sg13g2_nor2_1 _25290_ (.A(_07580_),
    .B(_07601_),
    .Y(_07604_));
 sg13g2_nor3_1 _25291_ (.A(net5933),
    .B(_07603_),
    .C(_07604_),
    .Y(_07605_));
 sg13g2_a21oi_1 _25292_ (.A1(net5933),
    .A2(_07597_),
    .Y(_07606_),
    .B1(_07605_));
 sg13g2_inv_1 _25293_ (.Y(_07607_),
    .A(_07606_));
 sg13g2_o21ai_1 _25294_ (.B1(net5917),
    .Y(_07608_),
    .A1(net5915),
    .A2(_07599_));
 sg13g2_a21o_1 _25295_ (.A2(_07599_),
    .A1(net5915),
    .B1(_07608_),
    .X(_07609_));
 sg13g2_nand2_1 _25296_ (.Y(_07610_),
    .A(_05278_),
    .B(_07609_));
 sg13g2_mux2_1 _25297_ (.A0(_07610_),
    .A1(_07609_),
    .S(_07606_),
    .X(_07611_));
 sg13g2_a21oi_1 _25298_ (.A1(_07577_),
    .A2(_07591_),
    .Y(_07612_),
    .B1(_07590_));
 sg13g2_nor2_1 _25299_ (.A(_07611_),
    .B(_07612_),
    .Y(_07613_));
 sg13g2_nand2_1 _25300_ (.Y(_07614_),
    .A(_07611_),
    .B(_07612_));
 sg13g2_nand2b_1 _25301_ (.Y(_07615_),
    .B(_07614_),
    .A_N(_07613_));
 sg13g2_a21oi_1 _25302_ (.A1(net5828),
    .A2(_07615_),
    .Y(_01403_),
    .B1(_07594_));
 sg13g2_nand2_1 _25303_ (.Y(_07616_),
    .A(net6250),
    .B(net5858));
 sg13g2_a22oi_1 _25304_ (.Y(_07617_),
    .B1(net5928),
    .B2(net6249),
    .A2(net5993),
    .A1(\atari2600.cpu.ABH[5] ));
 sg13g2_a22oi_1 _25305_ (.Y(_07618_),
    .B1(_05268_),
    .B2(_09098_),
    .A2(_05237_),
    .A1(\atari2600.cpu.DIMUX[5] ));
 sg13g2_and2_1 _25306_ (.A(_07617_),
    .B(_07618_),
    .X(_07619_));
 sg13g2_inv_1 _25307_ (.Y(_07620_),
    .A(_07619_));
 sg13g2_a22oi_1 _25308_ (.Y(_07621_),
    .B1(_05243_),
    .B2(\atari2600.cpu.DIMUX[4] ),
    .A2(net5991),
    .A1(\atari2600.cpu.PC[4] ));
 sg13g2_nand2b_1 _25309_ (.Y(_07622_),
    .B(net5875),
    .A_N(_07621_));
 sg13g2_o21ai_1 _25310_ (.B1(_05266_),
    .Y(_07623_),
    .A1(_07598_),
    .A2(_07622_));
 sg13g2_o21ai_1 _25311_ (.B1(_07623_),
    .Y(_07624_),
    .A1(_05264_),
    .A2(_07621_));
 sg13g2_a21oi_1 _25312_ (.A1(_07598_),
    .A2(_07622_),
    .Y(_07625_),
    .B1(net5933));
 sg13g2_a22oi_1 _25313_ (.Y(_07626_),
    .B1(_07624_),
    .B2(_07625_),
    .A2(_07620_),
    .A1(net5933));
 sg13g2_xor2_1 _25314_ (.B(_07621_),
    .A(net5915),
    .X(_07627_));
 sg13g2_nand2_1 _25315_ (.Y(_07628_),
    .A(net5917),
    .B(_07627_));
 sg13g2_and2_1 _25316_ (.A(_07626_),
    .B(_07628_),
    .X(_07629_));
 sg13g2_a21o_1 _25317_ (.A2(_07628_),
    .A1(_05278_),
    .B1(_07626_),
    .X(_07630_));
 sg13g2_nand2b_1 _25318_ (.Y(_07631_),
    .B(_07630_),
    .A_N(_07629_));
 sg13g2_nand2_1 _25319_ (.Y(_07632_),
    .A(\atari2600.cpu.adc_bcd ),
    .B(_08795_));
 sg13g2_a21oi_1 _25320_ (.A1(_07575_),
    .A2(_07593_),
    .Y(_07633_),
    .B1(_07632_));
 sg13g2_a221oi_1 _25321_ (.B2(_07633_),
    .C1(_07613_),
    .B1(_07614_),
    .A1(_07607_),
    .Y(_07634_),
    .A2(_07610_));
 sg13g2_xnor2_1 _25322_ (.Y(_07635_),
    .A(_07631_),
    .B(_07634_));
 sg13g2_o21ai_1 _25323_ (.B1(_07616_),
    .Y(_01404_),
    .A1(net5853),
    .A2(_07635_));
 sg13g2_nor2_1 _25324_ (.A(net6249),
    .B(net5854),
    .Y(_07636_));
 sg13g2_o21ai_1 _25325_ (.B1(_07630_),
    .Y(_07637_),
    .A1(_07629_),
    .A2(_07634_));
 sg13g2_a22oi_1 _25326_ (.Y(_07638_),
    .B1(_05237_),
    .B2(net5825),
    .A2(net5993),
    .A1(\atari2600.cpu.ABH[6] ));
 sg13g2_a22oi_1 _25327_ (.Y(_07639_),
    .B1(_09253_),
    .B2(_05268_),
    .A2(net5928),
    .A1(net6248));
 sg13g2_and2_1 _25328_ (.A(_07638_),
    .B(_07639_),
    .X(_07640_));
 sg13g2_nor2b_1 _25329_ (.A(_07640_),
    .B_N(net5933),
    .Y(_07641_));
 sg13g2_nand2_1 _25330_ (.Y(_07642_),
    .A(\atari2600.cpu.DIMUX[5] ),
    .B(_05243_));
 sg13g2_o21ai_1 _25331_ (.B1(_07642_),
    .Y(_07643_),
    .A1(_08595_),
    .A2(_08920_));
 sg13g2_nand2_1 _25332_ (.Y(_07644_),
    .A(net5875),
    .B(_07643_));
 sg13g2_o21ai_1 _25333_ (.B1(_05266_),
    .Y(_07645_),
    .A1(_07619_),
    .A2(_07644_));
 sg13g2_nand2_1 _25334_ (.Y(_07646_),
    .A(_05263_),
    .B(_07643_));
 sg13g2_a221oi_1 _25335_ (.B2(_07646_),
    .C1(net5933),
    .B1(_07645_),
    .A1(_07619_),
    .Y(_07647_),
    .A2(_07644_));
 sg13g2_or2_1 _25336_ (.X(_07648_),
    .B(_07647_),
    .A(_07641_));
 sg13g2_xnor2_1 _25337_ (.Y(_07649_),
    .A(net5915),
    .B(_07643_));
 sg13g2_nand2_1 _25338_ (.Y(_07650_),
    .A(net5917),
    .B(_07649_));
 sg13g2_nand2_1 _25339_ (.Y(_07651_),
    .A(_05278_),
    .B(_07650_));
 sg13g2_mux2_1 _25340_ (.A0(_07650_),
    .A1(_07651_),
    .S(_07648_),
    .X(_07652_));
 sg13g2_nor2b_1 _25341_ (.A(_07652_),
    .B_N(_07637_),
    .Y(_07653_));
 sg13g2_xor2_1 _25342_ (.B(_07652_),
    .A(_07637_),
    .X(_07654_));
 sg13g2_a21oi_1 _25343_ (.A1(net5829),
    .A2(_07654_),
    .Y(_01405_),
    .B1(_07636_));
 sg13g2_nor2_1 _25344_ (.A(net6248),
    .B(net5854),
    .Y(_07655_));
 sg13g2_a22oi_1 _25345_ (.Y(_07656_),
    .B1(_05243_),
    .B2(net5825),
    .A2(net5991),
    .A1(\atari2600.cpu.PC[6] ));
 sg13g2_nand2b_1 _25346_ (.Y(_07657_),
    .B(net5875),
    .A_N(_07656_));
 sg13g2_o21ai_1 _25347_ (.B1(_05266_),
    .Y(_07658_),
    .A1(_07640_),
    .A2(_07657_));
 sg13g2_o21ai_1 _25348_ (.B1(_07658_),
    .Y(_07659_),
    .A1(_05264_),
    .A2(_07656_));
 sg13g2_a21oi_1 _25349_ (.A1(_07640_),
    .A2(_07657_),
    .Y(_07660_),
    .B1(net5933));
 sg13g2_a22oi_1 _25350_ (.Y(_07661_),
    .B1(_07659_),
    .B2(_07660_),
    .A2(_05271_),
    .A1(net5933));
 sg13g2_o21ai_1 _25351_ (.B1(net5917),
    .Y(_07662_),
    .A1(net5915),
    .A2(_07656_));
 sg13g2_a21o_1 _25352_ (.A2(_07656_),
    .A1(net5915),
    .B1(_07662_),
    .X(_07663_));
 sg13g2_a21oi_1 _25353_ (.A1(_05278_),
    .A2(_07663_),
    .Y(_07664_),
    .B1(_07661_));
 sg13g2_a21o_1 _25354_ (.A2(_07663_),
    .A1(_07661_),
    .B1(_07664_),
    .X(_07665_));
 sg13g2_a21oi_1 _25355_ (.A1(_07648_),
    .A2(_07651_),
    .Y(_07666_),
    .B1(_07653_));
 sg13g2_nor2_1 _25356_ (.A(_07665_),
    .B(_07666_),
    .Y(_07667_));
 sg13g2_xnor2_1 _25357_ (.Y(_07668_),
    .A(_07665_),
    .B(_07666_));
 sg13g2_a21oi_1 _25358_ (.A1(net5829),
    .A2(_07668_),
    .Y(_01406_),
    .B1(_07655_));
 sg13g2_o21ai_1 _25359_ (.B1(_05279_),
    .Y(_07669_),
    .A1(_05260_),
    .A2(_05275_));
 sg13g2_nor2b_1 _25360_ (.A(_05276_),
    .B_N(_07669_),
    .Y(_07670_));
 sg13g2_nor2_1 _25361_ (.A(_07664_),
    .B(_07667_),
    .Y(_07671_));
 sg13g2_xnor2_1 _25362_ (.Y(_07672_),
    .A(_07670_),
    .B(_07671_));
 sg13g2_mux2_1 _25363_ (.A0(net7501),
    .A1(_07672_),
    .S(net5828),
    .X(_01407_));
 sg13g2_nor2_1 _25364_ (.A(net7155),
    .B(net5854),
    .Y(_07673_));
 sg13g2_a21oi_1 _25365_ (.A1(net5828),
    .A2(_07634_),
    .Y(_01408_),
    .B1(_07673_));
 sg13g2_nand2_1 _25366_ (.Y(_07674_),
    .A(net5934),
    .B(_07544_));
 sg13g2_o21ai_1 _25367_ (.B1(_07669_),
    .Y(_07675_),
    .A1(_05276_),
    .A2(_07671_));
 sg13g2_xor2_1 _25368_ (.B(_07675_),
    .A(_07674_),
    .X(_07676_));
 sg13g2_a21oi_1 _25369_ (.A1(_07654_),
    .A2(_07668_),
    .Y(_07677_),
    .B1(_07632_));
 sg13g2_a21oi_1 _25370_ (.A1(_07672_),
    .A2(_07677_),
    .Y(_07678_),
    .B1(net5858));
 sg13g2_a22oi_1 _25371_ (.Y(_01409_),
    .B1(_07676_),
    .B2(_07678_),
    .A2(net5858),
    .A1(_08592_));
 sg13g2_nand2_1 _25372_ (.Y(_07679_),
    .A(net7068),
    .B(net5858));
 sg13g2_o21ai_1 _25373_ (.B1(_08943_),
    .Y(_07680_),
    .A1(net6106),
    .A2(_08957_));
 sg13g2_nand2_1 _25374_ (.Y(_07681_),
    .A(_08771_),
    .B(_08920_));
 sg13g2_nor4_1 _25375_ (.A(_08788_),
    .B(_09033_),
    .C(_07680_),
    .D(_07681_),
    .Y(_07682_));
 sg13g2_nand4_1 _25376_ (.B(net5990),
    .C(_09074_),
    .A(_08847_),
    .Y(_07683_),
    .D(_07682_));
 sg13g2_nand2_1 _25377_ (.Y(_07684_),
    .A(_08810_),
    .B(_09074_));
 sg13g2_nor2_1 _25378_ (.A(net5994),
    .B(_07684_),
    .Y(_07685_));
 sg13g2_nand2_1 _25379_ (.Y(_07686_),
    .A(_08850_),
    .B(_07685_));
 sg13g2_nor2_2 _25380_ (.A(_08974_),
    .B(_07686_),
    .Y(_07687_));
 sg13g2_nand3_1 _25381_ (.B(net5990),
    .C(_07685_),
    .A(_08850_),
    .Y(_07688_));
 sg13g2_o21ai_1 _25382_ (.B1(net6253),
    .Y(_07689_),
    .A1(net5996),
    .A2(net5932));
 sg13g2_and2_1 _25383_ (.A(\atari2600.cpu.PC[0] ),
    .B(_08974_),
    .X(_07690_));
 sg13g2_o21ai_1 _25384_ (.B1(_07689_),
    .Y(_07691_),
    .A1(_00087_),
    .A2(_07688_));
 sg13g2_nor2_1 _25385_ (.A(_07690_),
    .B(_07691_),
    .Y(_07692_));
 sg13g2_o21ai_1 _25386_ (.B1(_07683_),
    .Y(_07693_),
    .A1(_07690_),
    .A2(_07691_));
 sg13g2_xor2_1 _25387_ (.B(_07692_),
    .A(_07683_),
    .X(_07694_));
 sg13g2_o21ai_1 _25388_ (.B1(_07679_),
    .Y(_01410_),
    .A1(net5858),
    .A2(_07694_));
 sg13g2_a221oi_1 _25389_ (.B2(net6252),
    .C1(_09130_),
    .B1(net5932),
    .A1(_08490_),
    .Y(_07695_),
    .A2(_08849_));
 sg13g2_o21ai_1 _25390_ (.B1(_07695_),
    .Y(_07696_),
    .A1(_00088_),
    .A2(net5870));
 sg13g2_nand2b_1 _25391_ (.Y(_07697_),
    .B(_07696_),
    .A_N(_07693_));
 sg13g2_nor2_1 _25392_ (.A(net4443),
    .B(net5854),
    .Y(_07698_));
 sg13g2_xor2_1 _25393_ (.B(_07696_),
    .A(_07693_),
    .X(_07699_));
 sg13g2_a21oi_1 _25394_ (.A1(net5854),
    .A2(_07699_),
    .Y(_01411_),
    .B1(_07698_));
 sg13g2_o21ai_1 _25395_ (.B1(_08850_),
    .Y(_07700_),
    .A1(_00076_),
    .A2(net5992));
 sg13g2_a21oi_1 _25396_ (.A1(net6251),
    .A2(net5932),
    .Y(_07701_),
    .B1(_07700_));
 sg13g2_o21ai_1 _25397_ (.B1(_07701_),
    .Y(_07702_),
    .A1(_00078_),
    .A2(net5870));
 sg13g2_nand2b_1 _25398_ (.Y(_07703_),
    .B(_07702_),
    .A_N(_07697_));
 sg13g2_nor2_1 _25399_ (.A(net3642),
    .B(net5855),
    .Y(_07704_));
 sg13g2_xor2_1 _25400_ (.B(_07702_),
    .A(_07697_),
    .X(_07705_));
 sg13g2_a21oi_1 _25401_ (.A1(net5855),
    .A2(_07705_),
    .Y(_01412_),
    .B1(_07704_));
 sg13g2_a21oi_1 _25402_ (.A1(\atari2600.cpu.ADD[3] ),
    .A2(net5931),
    .Y(_07706_),
    .B1(_08849_));
 sg13g2_o21ai_1 _25403_ (.B1(_07706_),
    .Y(_07707_),
    .A1(_00089_),
    .A2(net5870));
 sg13g2_nor2_1 _25404_ (.A(_09160_),
    .B(_07707_),
    .Y(_07708_));
 sg13g2_or2_1 _25405_ (.X(_07709_),
    .B(_07708_),
    .A(_07703_));
 sg13g2_nand2_1 _25406_ (.Y(_07710_),
    .A(net5830),
    .B(_07709_));
 sg13g2_a21oi_1 _25407_ (.A1(_07703_),
    .A2(_07708_),
    .Y(_07711_),
    .B1(_07710_));
 sg13g2_a21o_1 _25408_ (.A2(net5859),
    .A1(net7253),
    .B1(_07711_),
    .X(_01413_));
 sg13g2_nor2_1 _25409_ (.A(net7008),
    .B(net5830),
    .Y(_07712_));
 sg13g2_o21ai_1 _25410_ (.B1(net5870),
    .Y(_07713_),
    .A1(net6250),
    .A2(_08849_));
 sg13g2_o21ai_1 _25411_ (.B1(_07713_),
    .Y(_07714_),
    .A1(_00085_),
    .A2(net5870));
 sg13g2_nor2b_1 _25412_ (.A(_07709_),
    .B_N(_07714_),
    .Y(_07715_));
 sg13g2_xor2_1 _25413_ (.B(_07714_),
    .A(_07709_),
    .X(_07716_));
 sg13g2_a21oi_1 _25414_ (.A1(net5831),
    .A2(_07716_),
    .Y(_01414_),
    .B1(_07712_));
 sg13g2_a221oi_1 _25415_ (.B2(net6249),
    .C1(_08849_),
    .B1(net5932),
    .A1(_08596_),
    .Y(_07717_),
    .A2(net5994));
 sg13g2_o21ai_1 _25416_ (.B1(_07717_),
    .Y(_07718_),
    .A1(_00060_),
    .A2(net5870));
 sg13g2_nand2_1 _25417_ (.Y(_07719_),
    .A(_07715_),
    .B(_07718_));
 sg13g2_o21ai_1 _25418_ (.B1(net5831),
    .Y(_07720_),
    .A1(_07715_),
    .A2(_07718_));
 sg13g2_nand2b_1 _25419_ (.Y(_07721_),
    .B(_07719_),
    .A_N(_07720_));
 sg13g2_o21ai_1 _25420_ (.B1(_07721_),
    .Y(_01415_),
    .A1(_08595_),
    .A2(net5831));
 sg13g2_nor2_1 _25421_ (.A(net7145),
    .B(net5829),
    .Y(_07722_));
 sg13g2_o21ai_1 _25422_ (.B1(_08850_),
    .Y(_07723_),
    .A1(_00092_),
    .A2(net5992));
 sg13g2_a21oi_1 _25423_ (.A1(net6248),
    .A2(net5931),
    .Y(_07724_),
    .B1(_07723_));
 sg13g2_o21ai_1 _25424_ (.B1(_07724_),
    .Y(_07725_),
    .A1(_00061_),
    .A2(net5870));
 sg13g2_nor2b_1 _25425_ (.A(_07719_),
    .B_N(_07725_),
    .Y(_07726_));
 sg13g2_xor2_1 _25426_ (.B(_07725_),
    .A(_07719_),
    .X(_07727_));
 sg13g2_a21oi_1 _25427_ (.A1(net5828),
    .A2(_07727_),
    .Y(_01416_),
    .B1(_07722_));
 sg13g2_nor2_1 _25428_ (.A(net7196),
    .B(net5829),
    .Y(_07728_));
 sg13g2_a21oi_1 _25429_ (.A1(\atari2600.cpu.ADD[7] ),
    .A2(net5931),
    .Y(_07729_),
    .B1(_08849_));
 sg13g2_o21ai_1 _25430_ (.B1(_07729_),
    .Y(_07730_),
    .A1(_00062_),
    .A2(net5870));
 sg13g2_a21oi_1 _25431_ (.A1(_08599_),
    .A2(net5996),
    .Y(_07731_),
    .B1(_07730_));
 sg13g2_nor2b_2 _25432_ (.A(_07731_),
    .B_N(_07726_),
    .Y(_07732_));
 sg13g2_xor2_1 _25433_ (.B(_07731_),
    .A(_07726_),
    .X(_07733_));
 sg13g2_a21oi_1 _25434_ (.A1(net5829),
    .A2(_07733_),
    .Y(_01417_),
    .B1(_07728_));
 sg13g2_nand2_1 _25435_ (.Y(_07734_),
    .A(\atari2600.cpu.DIMUX[0] ),
    .B(net5932));
 sg13g2_nand2_2 _25436_ (.Y(_07735_),
    .A(_08850_),
    .B(_07688_));
 sg13g2_a221oi_1 _25437_ (.B2(net6253),
    .C1(_07735_),
    .B1(_08974_),
    .A1(\atari2600.cpu.ABH[0] ),
    .Y(_07736_),
    .A2(net5995));
 sg13g2_a22oi_1 _25438_ (.Y(_07737_),
    .B1(_07734_),
    .B2(_07736_),
    .A2(_07687_),
    .A1(_00063_));
 sg13g2_nand2_2 _25439_ (.Y(_07738_),
    .A(_07732_),
    .B(_07737_));
 sg13g2_o21ai_1 _25440_ (.B1(net5832),
    .Y(_07739_),
    .A1(_07732_),
    .A2(_07737_));
 sg13g2_nand2b_1 _25441_ (.Y(_07740_),
    .B(_07738_),
    .A_N(_07739_));
 sg13g2_o21ai_1 _25442_ (.B1(_07740_),
    .Y(_01418_),
    .A1(_08584_),
    .A2(net5832));
 sg13g2_a21oi_1 _25443_ (.A1(\atari2600.cpu.ABH[1] ),
    .A2(net5996),
    .Y(_07741_),
    .B1(_07735_));
 sg13g2_o21ai_1 _25444_ (.B1(_07741_),
    .Y(_07742_),
    .A1(_00074_),
    .A2(_08975_));
 sg13g2_a21oi_1 _25445_ (.A1(\atari2600.cpu.DIMUX[1] ),
    .A2(net5932),
    .Y(_07743_),
    .B1(_07742_));
 sg13g2_a21o_1 _25446_ (.A2(_07687_),
    .A1(_00064_),
    .B1(_07743_),
    .X(_07744_));
 sg13g2_a21oi_1 _25447_ (.A1(_07738_),
    .A2(_07744_),
    .Y(_07745_),
    .B1(net5859));
 sg13g2_o21ai_1 _25448_ (.B1(_07745_),
    .Y(_07746_),
    .A1(_07738_),
    .A2(_07744_));
 sg13g2_o21ai_1 _25449_ (.B1(_07746_),
    .Y(_01419_),
    .A1(_08579_),
    .A2(net5855));
 sg13g2_a221oi_1 _25450_ (.B2(net5827),
    .C1(_07735_),
    .B1(net5932),
    .A1(\atari2600.cpu.ABH[2] ),
    .Y(_07747_),
    .A2(net5994));
 sg13g2_o21ai_1 _25451_ (.B1(_07747_),
    .Y(_07748_),
    .A1(_00076_),
    .A2(net5990));
 sg13g2_o21ai_1 _25452_ (.B1(_07748_),
    .Y(_07749_),
    .A1(_08672_),
    .A2(_07688_));
 sg13g2_or3_1 _25453_ (.A(_07738_),
    .B(_07744_),
    .C(_07749_),
    .X(_07750_));
 sg13g2_o21ai_1 _25454_ (.B1(_07749_),
    .Y(_07751_),
    .A1(_07738_),
    .A2(_07744_));
 sg13g2_a21oi_1 _25455_ (.A1(_07750_),
    .A2(_07751_),
    .Y(_07752_),
    .B1(net5859));
 sg13g2_a21oi_1 _25456_ (.A1(_08581_),
    .A2(net5853),
    .Y(_01420_),
    .B1(_07752_));
 sg13g2_a221oi_1 _25457_ (.B2(net5826),
    .C1(_07735_),
    .B1(net5931),
    .A1(\atari2600.cpu.ABH[3] ),
    .Y(_07753_),
    .A2(net5994));
 sg13g2_o21ai_1 _25458_ (.B1(_07753_),
    .Y(_07754_),
    .A1(_00090_),
    .A2(net5990));
 sg13g2_o21ai_1 _25459_ (.B1(_07754_),
    .Y(_07755_),
    .A1(_08673_),
    .A2(_07688_));
 sg13g2_nor2_1 _25460_ (.A(_07750_),
    .B(_07755_),
    .Y(_07756_));
 sg13g2_a21oi_1 _25461_ (.A1(_07750_),
    .A2(_07755_),
    .Y(_07757_),
    .B1(net5859));
 sg13g2_nand2b_1 _25462_ (.Y(_07758_),
    .B(_07757_),
    .A_N(_07756_));
 sg13g2_o21ai_1 _25463_ (.B1(_07758_),
    .Y(_01421_),
    .A1(_08605_),
    .A2(net5830));
 sg13g2_nand2_1 _25464_ (.Y(_07759_),
    .A(\atari2600.cpu.DIMUX[4] ),
    .B(net5931));
 sg13g2_a221oi_1 _25465_ (.B2(net6250),
    .C1(_07735_),
    .B1(_08974_),
    .A1(\atari2600.cpu.ABH[4] ),
    .Y(_07760_),
    .A2(net5993));
 sg13g2_a22oi_1 _25466_ (.Y(_07761_),
    .B1(_07759_),
    .B2(_07760_),
    .A2(_07687_),
    .A1(_00067_));
 sg13g2_or2_1 _25467_ (.X(_07762_),
    .B(_07761_),
    .A(_07756_));
 sg13g2_nand2_1 _25468_ (.Y(_07763_),
    .A(_07756_),
    .B(_07761_));
 sg13g2_nand3_1 _25469_ (.B(_07762_),
    .C(_07763_),
    .A(net5830),
    .Y(_07764_));
 sg13g2_o21ai_1 _25470_ (.B1(_07764_),
    .Y(_01422_),
    .A1(_08598_),
    .A2(net5830));
 sg13g2_nor2_1 _25471_ (.A(net7214),
    .B(net5855),
    .Y(_07765_));
 sg13g2_nand2_1 _25472_ (.Y(_07766_),
    .A(\atari2600.cpu.DIMUX[5] ),
    .B(net5931));
 sg13g2_a221oi_1 _25473_ (.B2(_08596_),
    .C1(_07735_),
    .B1(_08974_),
    .A1(\atari2600.cpu.ABH[5] ),
    .Y(_07767_),
    .A2(net5993));
 sg13g2_a22oi_1 _25474_ (.Y(_07768_),
    .B1(_07766_),
    .B2(_07767_),
    .A2(_07687_),
    .A1(_00068_));
 sg13g2_nor2b_1 _25475_ (.A(_07763_),
    .B_N(_07768_),
    .Y(_07769_));
 sg13g2_xor2_1 _25476_ (.B(_07768_),
    .A(_07763_),
    .X(_07770_));
 sg13g2_a21oi_1 _25477_ (.A1(net5830),
    .A2(_07770_),
    .Y(_01423_),
    .B1(_07765_));
 sg13g2_nand2b_1 _25478_ (.Y(_07771_),
    .B(_08974_),
    .A_N(_00092_));
 sg13g2_a221oi_1 _25479_ (.B2(net5825),
    .C1(_07735_),
    .B1(net5931),
    .A1(\atari2600.cpu.ABH[6] ),
    .Y(_07772_),
    .A2(net5993));
 sg13g2_a22oi_1 _25480_ (.Y(_07773_),
    .B1(_07771_),
    .B2(_07772_),
    .A2(_07687_),
    .A1(_08659_));
 sg13g2_nand2_1 _25481_ (.Y(_07774_),
    .A(_07769_),
    .B(_07773_));
 sg13g2_o21ai_1 _25482_ (.B1(net5830),
    .Y(_07775_),
    .A1(_07769_),
    .A2(_07773_));
 sg13g2_nand2b_1 _25483_ (.Y(_07776_),
    .B(_07774_),
    .A_N(_07775_));
 sg13g2_o21ai_1 _25484_ (.B1(_07776_),
    .Y(_01424_),
    .A1(_08659_),
    .A2(net5830));
 sg13g2_nor2_1 _25485_ (.A(net7381),
    .B(net5855),
    .Y(_07777_));
 sg13g2_a221oi_1 _25486_ (.B2(\atari2600.cpu.DIMUX[7] ),
    .C1(_07735_),
    .B1(net5931),
    .A1(\atari2600.cpu.ABH[7] ),
    .Y(_07778_),
    .A2(net5993));
 sg13g2_o21ai_1 _25487_ (.B1(_07778_),
    .Y(_07779_),
    .A1(_00091_),
    .A2(net5990));
 sg13g2_o21ai_1 _25488_ (.B1(_07779_),
    .Y(_07780_),
    .A1(\atari2600.cpu.PC[15] ),
    .A2(_07688_));
 sg13g2_xnor2_1 _25489_ (.Y(_07781_),
    .A(_07774_),
    .B(_07780_));
 sg13g2_a21oi_1 _25490_ (.A1(net5831),
    .A2(_07781_),
    .Y(_01425_),
    .B1(_07777_));
 sg13g2_nor2_1 _25491_ (.A(net5255),
    .B(_07321_),
    .Y(_07782_));
 sg13g2_nor2_1 _25492_ (.A(net4841),
    .B(net5037),
    .Y(_07783_));
 sg13g2_a21oi_1 _25493_ (.A1(net5759),
    .A2(net5037),
    .Y(_01426_),
    .B1(_07783_));
 sg13g2_nor2_1 _25494_ (.A(net3720),
    .B(net5037),
    .Y(_07784_));
 sg13g2_a21oi_1 _25495_ (.A1(net5780),
    .A2(net5037),
    .Y(_01427_),
    .B1(_07784_));
 sg13g2_nor2_1 _25496_ (.A(net4250),
    .B(net5038),
    .Y(_07785_));
 sg13g2_a21oi_1 _25497_ (.A1(net5710),
    .A2(net5038),
    .Y(_01428_),
    .B1(_07785_));
 sg13g2_nor2_1 _25498_ (.A(net3296),
    .B(_07782_),
    .Y(_07786_));
 sg13g2_a21oi_1 _25499_ (.A1(net5687),
    .A2(net5038),
    .Y(_01429_),
    .B1(_07786_));
 sg13g2_nor2_1 _25500_ (.A(net3060),
    .B(net5038),
    .Y(_07787_));
 sg13g2_a21oi_1 _25501_ (.A1(net5670),
    .A2(net5038),
    .Y(_01430_),
    .B1(_07787_));
 sg13g2_nor2_1 _25502_ (.A(net3662),
    .B(net5037),
    .Y(_07788_));
 sg13g2_a21oi_1 _25503_ (.A1(net5585),
    .A2(net5037),
    .Y(_01431_),
    .B1(_07788_));
 sg13g2_nor2_1 _25504_ (.A(net3292),
    .B(net5038),
    .Y(_07789_));
 sg13g2_a21oi_1 _25505_ (.A1(net5647),
    .A2(net5038),
    .Y(_01432_),
    .B1(_07789_));
 sg13g2_nor2_1 _25506_ (.A(net3814),
    .B(net5037),
    .Y(_07790_));
 sg13g2_a21oi_1 _25507_ (.A1(net5622),
    .A2(net5037),
    .Y(_01433_),
    .B1(_07790_));
 sg13g2_nor2_1 _25508_ (.A(net5238),
    .B(_07321_),
    .Y(_07791_));
 sg13g2_nor2_1 _25509_ (.A(net3561),
    .B(net5035),
    .Y(_07792_));
 sg13g2_a21oi_1 _25510_ (.A1(net5759),
    .A2(net5035),
    .Y(_01434_),
    .B1(_07792_));
 sg13g2_nor2_1 _25511_ (.A(net7088),
    .B(net5035),
    .Y(_07793_));
 sg13g2_a21oi_1 _25512_ (.A1(net5780),
    .A2(net5035),
    .Y(_01435_),
    .B1(_07793_));
 sg13g2_nor2_1 _25513_ (.A(net3394),
    .B(net5036),
    .Y(_07794_));
 sg13g2_a21oi_1 _25514_ (.A1(net5710),
    .A2(net5036),
    .Y(_01436_),
    .B1(_07794_));
 sg13g2_nor2_1 _25515_ (.A(net3463),
    .B(net5036),
    .Y(_07795_));
 sg13g2_a21oi_1 _25516_ (.A1(net5687),
    .A2(net5036),
    .Y(_01437_),
    .B1(_07795_));
 sg13g2_nor2_1 _25517_ (.A(net3408),
    .B(net5036),
    .Y(_07796_));
 sg13g2_a21oi_1 _25518_ (.A1(net5667),
    .A2(net5036),
    .Y(_01438_),
    .B1(_07796_));
 sg13g2_nor2_1 _25519_ (.A(net3728),
    .B(net5035),
    .Y(_07797_));
 sg13g2_a21oi_1 _25520_ (.A1(net5585),
    .A2(net5035),
    .Y(_01439_),
    .B1(_07797_));
 sg13g2_nor2_1 _25521_ (.A(net3427),
    .B(net5036),
    .Y(_07798_));
 sg13g2_a21oi_1 _25522_ (.A1(net5647),
    .A2(net5036),
    .Y(_01440_),
    .B1(_07798_));
 sg13g2_nor2_1 _25523_ (.A(net3197),
    .B(net5035),
    .Y(_07799_));
 sg13g2_a21oi_1 _25524_ (.A1(net5622),
    .A2(net5035),
    .Y(_01441_),
    .B1(_07799_));
 sg13g2_a21oi_1 _25525_ (.A1(net7447),
    .A2(net5929),
    .Y(_07800_),
    .B1(_05281_));
 sg13g2_nor2_1 _25526_ (.A(net6530),
    .B(_07800_),
    .Y(_01442_));
 sg13g2_a21oi_1 _25527_ (.A1(net6246),
    .A2(net7447),
    .Y(_07801_),
    .B1(_08679_));
 sg13g2_o21ai_1 _25528_ (.B1(_07801_),
    .Y(_07802_),
    .A1(net6246),
    .A2(net7447));
 sg13g2_o21ai_1 _25529_ (.B1(net6571),
    .Y(_07803_),
    .A1(net6246),
    .A2(_08710_));
 sg13g2_a21oi_1 _25530_ (.A1(_08710_),
    .A2(_07802_),
    .Y(_01443_),
    .B1(_07803_));
 sg13g2_and3_1 _25531_ (.X(_01444_),
    .A(net2941),
    .B(net6570),
    .C(net5930));
 sg13g2_and3_1 _25532_ (.X(_01445_),
    .A(net2942),
    .B(net6570),
    .C(net5930));
 sg13g2_and3_1 _25533_ (.X(_01446_),
    .A(net2951),
    .B(net6570),
    .C(net5930));
 sg13g2_and3_1 _25534_ (.X(_01447_),
    .A(net2954),
    .B(net6570),
    .C(net5930));
 sg13g2_and3_1 _25535_ (.X(_01448_),
    .A(net2945),
    .B(net6570),
    .C(net5929));
 sg13g2_and3_1 _25536_ (.X(_01449_),
    .A(net2948),
    .B(net6571),
    .C(net5929));
 sg13g2_nand3_1 _25537_ (.B(net6571),
    .C(net5929),
    .A(\atari2600.clk_counter[8] ),
    .Y(_07804_));
 sg13g2_nand2_1 _25538_ (.Y(_07805_),
    .A(_08634_),
    .B(_07801_));
 sg13g2_o21ai_1 _25539_ (.B1(_07804_),
    .Y(_01450_),
    .A1(_09471_),
    .A2(net3066));
 sg13g2_nand3_1 _25540_ (.B(_09345_),
    .C(net5251),
    .A(_09262_),
    .Y(_07806_));
 sg13g2_mux2_1 _25541_ (.A0(net5742),
    .A1(net4699),
    .S(_07806_),
    .X(_01451_));
 sg13g2_mux2_1 _25542_ (.A0(net5747),
    .A1(net4587),
    .S(_07806_),
    .X(_01452_));
 sg13g2_mux2_1 _25543_ (.A0(net5619),
    .A1(net4907),
    .S(_07806_),
    .X(_01453_));
 sg13g2_mux2_1 _25544_ (.A0(net5612),
    .A1(net6638),
    .S(_07806_),
    .X(_01454_));
 sg13g2_mux2_1 _25545_ (.A0(net5609),
    .A1(net4857),
    .S(_07806_),
    .X(_01455_));
 sg13g2_mux2_1 _25546_ (.A0(net5583),
    .A1(net7093),
    .S(_07806_),
    .X(_01456_));
 sg13g2_mux2_1 _25547_ (.A0(net5579),
    .A1(net6630),
    .S(_07806_),
    .X(_01457_));
 sg13g2_mux2_1 _25548_ (.A0(net5645),
    .A1(net4630),
    .S(_07806_),
    .X(_01458_));
 sg13g2_nor2_1 _25549_ (.A(net5255),
    .B(_03134_),
    .Y(_07807_));
 sg13g2_nor2_1 _25550_ (.A(net4382),
    .B(net5034),
    .Y(_07808_));
 sg13g2_a21oi_1 _25551_ (.A1(net5769),
    .A2(net5034),
    .Y(_01459_),
    .B1(_07808_));
 sg13g2_nor2_1 _25552_ (.A(net3819),
    .B(net5032),
    .Y(_07809_));
 sg13g2_a21oi_1 _25553_ (.A1(net5789),
    .A2(net5032),
    .Y(_01460_),
    .B1(_07809_));
 sg13g2_nor2_1 _25554_ (.A(net3228),
    .B(net5034),
    .Y(_07810_));
 sg13g2_a21oi_1 _25555_ (.A1(net5719),
    .A2(net5034),
    .Y(_01461_),
    .B1(_07810_));
 sg13g2_nor2_1 _25556_ (.A(net3922),
    .B(net5033),
    .Y(_07811_));
 sg13g2_a21oi_1 _25557_ (.A1(net5695),
    .A2(net5033),
    .Y(_01462_),
    .B1(_07811_));
 sg13g2_nor2_1 _25558_ (.A(net3251),
    .B(net5032),
    .Y(_07812_));
 sg13g2_a21oi_1 _25559_ (.A1(net5672),
    .A2(net5032),
    .Y(_01463_),
    .B1(_07812_));
 sg13g2_nor2_1 _25560_ (.A(net3076),
    .B(net5033),
    .Y(_07813_));
 sg13g2_a21oi_1 _25561_ (.A1(net5593),
    .A2(net5033),
    .Y(_01464_),
    .B1(_07813_));
 sg13g2_nor2_1 _25562_ (.A(net4437),
    .B(net5032),
    .Y(_07814_));
 sg13g2_a21oi_1 _25563_ (.A1(net5656),
    .A2(net5032),
    .Y(_01465_),
    .B1(_07814_));
 sg13g2_nor2_1 _25564_ (.A(net3650),
    .B(net5032),
    .Y(_07815_));
 sg13g2_a21oi_1 _25565_ (.A1(net5630),
    .A2(net5032),
    .Y(_01466_),
    .B1(_07815_));
 sg13g2_nor2_1 _25566_ (.A(_09441_),
    .B(_04792_),
    .Y(_07816_));
 sg13g2_nor2_1 _25567_ (.A(net3532),
    .B(net5030),
    .Y(_07817_));
 sg13g2_a21oi_1 _25568_ (.A1(net5768),
    .A2(net5030),
    .Y(_01467_),
    .B1(_07817_));
 sg13g2_nor2_1 _25569_ (.A(net4414),
    .B(net5031),
    .Y(_07818_));
 sg13g2_a21oi_1 _25570_ (.A1(net5788),
    .A2(net5031),
    .Y(_01468_),
    .B1(_07818_));
 sg13g2_nor2_1 _25571_ (.A(net3120),
    .B(_07816_),
    .Y(_07819_));
 sg13g2_a21oi_1 _25572_ (.A1(net5718),
    .A2(net5031),
    .Y(_01469_),
    .B1(_07819_));
 sg13g2_nor2_1 _25573_ (.A(net3402),
    .B(net5030),
    .Y(_07820_));
 sg13g2_a21oi_1 _25574_ (.A1(net5695),
    .A2(net5030),
    .Y(_01470_),
    .B1(_07820_));
 sg13g2_nor2_1 _25575_ (.A(net3196),
    .B(net5031),
    .Y(_07821_));
 sg13g2_a21oi_1 _25576_ (.A1(net5674),
    .A2(net5031),
    .Y(_01471_),
    .B1(_07821_));
 sg13g2_nor2_1 _25577_ (.A(net3059),
    .B(net5031),
    .Y(_07822_));
 sg13g2_a21oi_1 _25578_ (.A1(net5593),
    .A2(net5031),
    .Y(_01472_),
    .B1(_07822_));
 sg13g2_nor2_1 _25579_ (.A(net3302),
    .B(net5030),
    .Y(_07823_));
 sg13g2_a21oi_1 _25580_ (.A1(net5657),
    .A2(net5030),
    .Y(_01473_),
    .B1(_07823_));
 sg13g2_nor2_1 _25581_ (.A(net3330),
    .B(net5030),
    .Y(_07824_));
 sg13g2_a21oi_1 _25582_ (.A1(net5635),
    .A2(net5030),
    .Y(_01474_),
    .B1(_07824_));
 sg13g2_o21ai_1 _25583_ (.B1(net6544),
    .Y(_07825_),
    .A1(\flash_rom.spi_select ),
    .A2(_03188_));
 sg13g2_inv_2 _25584_ (.Y(_07826_),
    .A(_07825_));
 sg13g2_nor2_2 _25585_ (.A(net7303),
    .B(_11054_),
    .Y(_07827_));
 sg13g2_nand2_2 _25586_ (.Y(_07828_),
    .A(net6245),
    .B(_11056_));
 sg13g2_nor3_2 _25587_ (.A(\flash_rom.nibbles_remaining[2] ),
    .B(\flash_rom.nibbles_remaining[1] ),
    .C(\flash_rom.nibbles_remaining[0] ),
    .Y(_07829_));
 sg13g2_nand2_1 _25588_ (.Y(_07830_),
    .A(net7495),
    .B(_07829_));
 sg13g2_nor2_1 _25589_ (.A(_07828_),
    .B(_07830_),
    .Y(_07831_));
 sg13g2_nor2_1 _25590_ (.A(_07827_),
    .B(_07831_),
    .Y(_07832_));
 sg13g2_nor2_1 _25591_ (.A(_07825_),
    .B(_07832_),
    .Y(_01475_));
 sg13g2_nor2b_1 _25592_ (.A(\gamepad_pmod.driver.pmod_clk_prev ),
    .B_N(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .Y(_07833_));
 sg13g2_nor2_1 _25593_ (.A(net6523),
    .B(net6038),
    .Y(_07834_));
 sg13g2_a22oi_1 _25594_ (.Y(_01476_),
    .B1(net6004),
    .B2(_08486_),
    .A2(net6038),
    .A1(_08488_));
 sg13g2_a22oi_1 _25595_ (.Y(_01477_),
    .B1(net6004),
    .B2(_08485_),
    .A2(net6038),
    .A1(_08486_));
 sg13g2_a22oi_1 _25596_ (.Y(_01478_),
    .B1(net6004),
    .B2(_08484_),
    .A2(net6038),
    .A1(_08485_));
 sg13g2_a22oi_1 _25597_ (.Y(_01479_),
    .B1(net6004),
    .B2(_08483_),
    .A2(net6038),
    .A1(_08484_));
 sg13g2_a22oi_1 _25598_ (.Y(_01480_),
    .B1(net6004),
    .B2(_08482_),
    .A2(net6038),
    .A1(_08483_));
 sg13g2_a22oi_1 _25599_ (.Y(_01481_),
    .B1(net6004),
    .B2(_08481_),
    .A2(net6038),
    .A1(_08482_));
 sg13g2_a22oi_1 _25600_ (.Y(_01482_),
    .B1(net6004),
    .B2(_08480_),
    .A2(net6038),
    .A1(_08481_));
 sg13g2_a22oi_1 _25601_ (.Y(_01483_),
    .B1(net6005),
    .B2(_08479_),
    .A2(net6039),
    .A1(_08480_));
 sg13g2_a22oi_1 _25602_ (.Y(_01484_),
    .B1(net6004),
    .B2(_08478_),
    .A2(net6039),
    .A1(_08479_));
 sg13g2_a22oi_1 _25603_ (.Y(_01485_),
    .B1(net6005),
    .B2(_08477_),
    .A2(net6039),
    .A1(_08478_));
 sg13g2_a22oi_1 _25604_ (.Y(_01486_),
    .B1(net6005),
    .B2(_08476_),
    .A2(net6039),
    .A1(_08477_));
 sg13g2_a22oi_1 _25605_ (.Y(_01487_),
    .B1(net6005),
    .B2(_08475_),
    .A2(net6039),
    .A1(_08476_));
 sg13g2_nor2_1 _25606_ (.A(net6523),
    .B(_08657_),
    .Y(_01488_));
 sg13g2_and2_1 _25607_ (.A(net6544),
    .B(net2940),
    .X(_01489_));
 sg13g2_and2_1 _25608_ (.A(net6544),
    .B(net6),
    .X(_01490_));
 sg13g2_and2_1 _25609_ (.A(net6544),
    .B(net2938),
    .X(_01491_));
 sg13g2_nor2_1 _25610_ (.A(_03021_),
    .B(net5248),
    .Y(_07835_));
 sg13g2_nor2_1 _25611_ (.A(net3042),
    .B(net5103),
    .Y(_07836_));
 sg13g2_a21oi_1 _25612_ (.A1(net5774),
    .A2(net5103),
    .Y(_01492_),
    .B1(_07836_));
 sg13g2_nor2_1 _25613_ (.A(net3572),
    .B(net5103),
    .Y(_07837_));
 sg13g2_a21oi_1 _25614_ (.A1(net5794),
    .A2(net5103),
    .Y(_01493_),
    .B1(_07837_));
 sg13g2_nor2_1 _25615_ (.A(net3610),
    .B(net5104),
    .Y(_07838_));
 sg13g2_a21oi_1 _25616_ (.A1(net5724),
    .A2(net5104),
    .Y(_01494_),
    .B1(_07838_));
 sg13g2_nor2_1 _25617_ (.A(net3070),
    .B(net5103),
    .Y(_07839_));
 sg13g2_a21oi_1 _25618_ (.A1(net5700),
    .A2(net5103),
    .Y(_01495_),
    .B1(_07839_));
 sg13g2_nor2_1 _25619_ (.A(net3943),
    .B(net5103),
    .Y(_07840_));
 sg13g2_a21oi_1 _25620_ (.A1(net5680),
    .A2(net5103),
    .Y(_01496_),
    .B1(_07840_));
 sg13g2_nor2_1 _25621_ (.A(net3588),
    .B(_07835_),
    .Y(_07841_));
 sg13g2_a21oi_1 _25622_ (.A1(net5601),
    .A2(net5104),
    .Y(_01497_),
    .B1(_07841_));
 sg13g2_nor2_1 _25623_ (.A(net3851),
    .B(net5104),
    .Y(_07842_));
 sg13g2_a21oi_1 _25624_ (.A1(net5658),
    .A2(net5104),
    .Y(_01498_),
    .B1(_07842_));
 sg13g2_nor2_1 _25625_ (.A(net3385),
    .B(net5104),
    .Y(_07843_));
 sg13g2_a21oi_1 _25626_ (.A1(net5636),
    .A2(net5104),
    .Y(_01499_),
    .B1(_07843_));
 sg13g2_nor2_1 _25627_ (.A(_09331_),
    .B(net5249),
    .Y(_07844_));
 sg13g2_nor2_1 _25628_ (.A(net3222),
    .B(net5029),
    .Y(_07845_));
 sg13g2_a21oi_1 _25629_ (.A1(net5761),
    .A2(net5029),
    .Y(_01500_),
    .B1(_07845_));
 sg13g2_nor2_1 _25630_ (.A(net3085),
    .B(net5028),
    .Y(_07846_));
 sg13g2_a21oi_1 _25631_ (.A1(net5781),
    .A2(net5028),
    .Y(_01501_),
    .B1(_07846_));
 sg13g2_nor2_1 _25632_ (.A(net4078),
    .B(net5029),
    .Y(_07847_));
 sg13g2_a21oi_1 _25633_ (.A1(net5710),
    .A2(net5029),
    .Y(_01502_),
    .B1(_07847_));
 sg13g2_nor2_1 _25634_ (.A(net3737),
    .B(net5028),
    .Y(_07848_));
 sg13g2_a21oi_1 _25635_ (.A1(net5686),
    .A2(net5028),
    .Y(_01503_),
    .B1(_07848_));
 sg13g2_nor2_1 _25636_ (.A(net3151),
    .B(net5029),
    .Y(_07849_));
 sg13g2_a21oi_1 _25637_ (.A1(net5667),
    .A2(_07844_),
    .Y(_01504_),
    .B1(_07849_));
 sg13g2_nor2_1 _25638_ (.A(net3032),
    .B(net5028),
    .Y(_07850_));
 sg13g2_a21oi_1 _25639_ (.A1(net5587),
    .A2(net5028),
    .Y(_01505_),
    .B1(_07850_));
 sg13g2_nor2_1 _25640_ (.A(net3279),
    .B(net5028),
    .Y(_07851_));
 sg13g2_a21oi_1 _25641_ (.A1(net5649),
    .A2(net5028),
    .Y(_01506_),
    .B1(_07851_));
 sg13g2_nor2_1 _25642_ (.A(net3090),
    .B(net5029),
    .Y(_07852_));
 sg13g2_a21oi_1 _25643_ (.A1(net5625),
    .A2(net5029),
    .Y(_01507_),
    .B1(_07852_));
 sg13g2_nand2_1 _25644_ (.Y(_07853_),
    .A(\hvsync_gen.vga.vpos[0] ),
    .B(_03198_));
 sg13g2_nand2_1 _25645_ (.Y(_07854_),
    .A(\hvsync_gen.vga.vpos[3] ),
    .B(\hvsync_gen.vga.vpos[2] ));
 sg13g2_nor4_1 _25646_ (.A(_08572_),
    .B(\hvsync_gen.vga.vpos[8] ),
    .C(\hvsync_gen.vga.vpos[0] ),
    .D(_07854_),
    .Y(_07855_));
 sg13g2_a21oi_1 _25647_ (.A1(_09040_),
    .A2(_07855_),
    .Y(_07856_),
    .B1(net6541));
 sg13g2_nand2_1 _25648_ (.Y(_07857_),
    .A(_03197_),
    .B(_07856_));
 sg13g2_o21ai_1 _25649_ (.B1(_07853_),
    .Y(_01508_),
    .A1(_08487_),
    .A2(_07857_));
 sg13g2_nand2_1 _25650_ (.Y(_07858_),
    .A(net7321),
    .B(_03198_));
 sg13g2_nand2_1 _25651_ (.Y(_07859_),
    .A(net7321),
    .B(\hvsync_gen.vga.vpos[0] ));
 sg13g2_xnor2_1 _25652_ (.Y(_07860_),
    .A(net7321),
    .B(\hvsync_gen.vga.vpos[0] ));
 sg13g2_o21ai_1 _25653_ (.B1(_07858_),
    .Y(_01509_),
    .A1(_07857_),
    .A2(_07860_));
 sg13g2_nor2_1 _25654_ (.A(_03198_),
    .B(_07859_),
    .Y(_07861_));
 sg13g2_and2_1 _25655_ (.A(net7412),
    .B(_07861_),
    .X(_07862_));
 sg13g2_nor2_2 _25656_ (.A(_03198_),
    .B(_07856_),
    .Y(_07863_));
 sg13g2_nor2_1 _25657_ (.A(net7412),
    .B(_07861_),
    .Y(_07864_));
 sg13g2_nor3_1 _25658_ (.A(_07862_),
    .B(_07863_),
    .C(_07864_),
    .Y(_01510_));
 sg13g2_nor2_1 _25659_ (.A(net7456),
    .B(_07862_),
    .Y(_07865_));
 sg13g2_and2_1 _25660_ (.A(net7456),
    .B(_07862_),
    .X(_07866_));
 sg13g2_nor3_1 _25661_ (.A(_07863_),
    .B(_07865_),
    .C(_07866_),
    .Y(_01511_));
 sg13g2_nand3_1 _25662_ (.B(\hvsync_gen.vga.vpos[3] ),
    .C(\hvsync_gen.vga.vpos[2] ),
    .A(\hvsync_gen.vga.vpos[4] ),
    .Y(_07867_));
 sg13g2_xnor2_1 _25663_ (.Y(_07868_),
    .A(net7442),
    .B(_07866_));
 sg13g2_nor2_1 _25664_ (.A(_07863_),
    .B(_07868_),
    .Y(_01512_));
 sg13g2_a21oi_1 _25665_ (.A1(\hvsync_gen.vga.vpos[4] ),
    .A2(_07866_),
    .Y(_07869_),
    .B1(net7178));
 sg13g2_and3_1 _25666_ (.X(_07870_),
    .A(net7178),
    .B(\hvsync_gen.vga.vpos[4] ),
    .C(_07866_));
 sg13g2_nor3_1 _25667_ (.A(_07863_),
    .B(net7179),
    .C(_07870_),
    .Y(_01513_));
 sg13g2_nor2_1 _25668_ (.A(net7433),
    .B(_07870_),
    .Y(_07871_));
 sg13g2_and2_1 _25669_ (.A(net7433),
    .B(_07870_),
    .X(_07872_));
 sg13g2_nor3_1 _25670_ (.A(_07863_),
    .B(net7434),
    .C(_07872_),
    .Y(_01514_));
 sg13g2_xnor2_1 _25671_ (.Y(_07873_),
    .A(net7437),
    .B(_07872_));
 sg13g2_nor2_1 _25672_ (.A(_07863_),
    .B(_07873_),
    .Y(_01515_));
 sg13g2_a21oi_1 _25673_ (.A1(\hvsync_gen.vga.vpos[7] ),
    .A2(_07872_),
    .Y(_07874_),
    .B1(net7239));
 sg13g2_nor3_1 _25674_ (.A(_09233_),
    .B(_07859_),
    .C(_07867_),
    .Y(_07875_));
 sg13g2_a21oi_1 _25675_ (.A1(_03199_),
    .A2(_07875_),
    .Y(_07876_),
    .B1(_07863_));
 sg13g2_nor2b_1 _25676_ (.A(net7240),
    .B_N(_07876_),
    .Y(_01516_));
 sg13g2_nand2_1 _25677_ (.Y(_07877_),
    .A(net7131),
    .B(_07876_));
 sg13g2_nand2_1 _25678_ (.Y(_07878_),
    .A(_08572_),
    .B(_07875_));
 sg13g2_o21ai_1 _25679_ (.B1(_07877_),
    .Y(_01517_),
    .A1(_07857_),
    .A2(_07878_));
 sg13g2_and2_1 _25680_ (.A(net6546),
    .B(net5),
    .X(_01518_));
 sg13g2_and2_1 _25681_ (.A(net6546),
    .B(net2937),
    .X(_01519_));
 sg13g2_nand3_1 _25682_ (.B(_09321_),
    .C(net5253),
    .A(net5551),
    .Y(_07879_));
 sg13g2_mux2_1 _25683_ (.A0(net5739),
    .A1(net4715),
    .S(_07879_),
    .X(_01520_));
 sg13g2_mux2_1 _25684_ (.A0(net5749),
    .A1(net6607),
    .S(_07879_),
    .X(_01521_));
 sg13g2_mux2_1 _25685_ (.A0(net5618),
    .A1(net4678),
    .S(_07879_),
    .X(_01522_));
 sg13g2_mux2_1 _25686_ (.A0(net5612),
    .A1(net4743),
    .S(_07879_),
    .X(_01523_));
 sg13g2_mux2_1 _25687_ (.A0(net5606),
    .A1(net4702),
    .S(_07879_),
    .X(_01524_));
 sg13g2_mux2_1 _25688_ (.A0(net5581),
    .A1(net4763),
    .S(_07879_),
    .X(_01525_));
 sg13g2_mux2_1 _25689_ (.A0(net5576),
    .A1(net6735),
    .S(_07879_),
    .X(_01526_));
 sg13g2_mux2_1 _25690_ (.A0(net5644),
    .A1(net7034),
    .S(_07879_),
    .X(_01527_));
 sg13g2_nor2_1 _25691_ (.A(_09422_),
    .B(net5237),
    .Y(_07880_));
 sg13g2_nor2_1 _25692_ (.A(net3269),
    .B(net5027),
    .Y(_07881_));
 sg13g2_a21oi_1 _25693_ (.A1(net5760),
    .A2(net5027),
    .Y(_01528_),
    .B1(_07881_));
 sg13g2_nor2_1 _25694_ (.A(net3543),
    .B(net5026),
    .Y(_07882_));
 sg13g2_a21oi_1 _25695_ (.A1(net5780),
    .A2(net5026),
    .Y(_01529_),
    .B1(_07882_));
 sg13g2_nor2_1 _25696_ (.A(net3236),
    .B(net5026),
    .Y(_07883_));
 sg13g2_a21oi_1 _25697_ (.A1(net5709),
    .A2(net5026),
    .Y(_01530_),
    .B1(_07883_));
 sg13g2_nor2_1 _25698_ (.A(net4490),
    .B(net5027),
    .Y(_07884_));
 sg13g2_a21oi_1 _25699_ (.A1(net5686),
    .A2(net5027),
    .Y(_01531_),
    .B1(_07884_));
 sg13g2_nor2_1 _25700_ (.A(net3149),
    .B(net5026),
    .Y(_07885_));
 sg13g2_a21oi_1 _25701_ (.A1(net5666),
    .A2(net5026),
    .Y(_01532_),
    .B1(_07885_));
 sg13g2_nor2_1 _25702_ (.A(net3600),
    .B(net5027),
    .Y(_07886_));
 sg13g2_a21oi_1 _25703_ (.A1(net5586),
    .A2(_07880_),
    .Y(_01533_),
    .B1(_07886_));
 sg13g2_nor2_1 _25704_ (.A(net4304),
    .B(net5027),
    .Y(_07887_));
 sg13g2_a21oi_1 _25705_ (.A1(net5647),
    .A2(net5027),
    .Y(_01534_),
    .B1(_07887_));
 sg13g2_nor2_1 _25706_ (.A(net4030),
    .B(net5026),
    .Y(_07888_));
 sg13g2_a21oi_1 _25707_ (.A1(net5623),
    .A2(net5026),
    .Y(_01535_),
    .B1(_07888_));
 sg13g2_nor2_1 _25708_ (.A(_09441_),
    .B(net5238),
    .Y(_07889_));
 sg13g2_nor2_1 _25709_ (.A(net3216),
    .B(net5025),
    .Y(_07890_));
 sg13g2_a21oi_1 _25710_ (.A1(net5768),
    .A2(net5025),
    .Y(_01536_),
    .B1(_07890_));
 sg13g2_nor2_1 _25711_ (.A(net3368),
    .B(net5024),
    .Y(_07891_));
 sg13g2_a21oi_1 _25712_ (.A1(net5788),
    .A2(net5024),
    .Y(_01537_),
    .B1(_07891_));
 sg13g2_nor2_1 _25713_ (.A(net3607),
    .B(net5025),
    .Y(_07892_));
 sg13g2_a21oi_1 _25714_ (.A1(net5718),
    .A2(net5025),
    .Y(_01538_),
    .B1(_07892_));
 sg13g2_nor2_1 _25715_ (.A(net3459),
    .B(net5025),
    .Y(_07893_));
 sg13g2_a21oi_1 _25716_ (.A1(net5695),
    .A2(net5025),
    .Y(_01539_),
    .B1(_07893_));
 sg13g2_nor2_1 _25717_ (.A(net3845),
    .B(net5024),
    .Y(_07894_));
 sg13g2_a21oi_1 _25718_ (.A1(net5674),
    .A2(net5024),
    .Y(_01540_),
    .B1(_07894_));
 sg13g2_nor2_1 _25719_ (.A(net4522),
    .B(net5024),
    .Y(_07895_));
 sg13g2_a21oi_1 _25720_ (.A1(net5593),
    .A2(net5024),
    .Y(_01541_),
    .B1(_07895_));
 sg13g2_nor2_1 _25721_ (.A(net3298),
    .B(net5024),
    .Y(_07896_));
 sg13g2_a21oi_1 _25722_ (.A1(net5655),
    .A2(net5024),
    .Y(_01542_),
    .B1(_07896_));
 sg13g2_nor2_1 _25723_ (.A(net3328),
    .B(net5025),
    .Y(_07897_));
 sg13g2_a21oi_1 _25724_ (.A1(net5630),
    .A2(net5025),
    .Y(_01543_),
    .B1(_07897_));
 sg13g2_nor2_1 _25725_ (.A(_09422_),
    .B(net5259),
    .Y(_07898_));
 sg13g2_nor2_1 _25726_ (.A(net4259),
    .B(net5023),
    .Y(_07899_));
 sg13g2_a21oi_1 _25727_ (.A1(net5759),
    .A2(net5023),
    .Y(_01544_),
    .B1(_07899_));
 sg13g2_nor2_1 _25728_ (.A(net4141),
    .B(net5022),
    .Y(_07900_));
 sg13g2_a21oi_1 _25729_ (.A1(net5780),
    .A2(net5022),
    .Y(_01545_),
    .B1(_07900_));
 sg13g2_nor2_1 _25730_ (.A(net3361),
    .B(net5022),
    .Y(_07901_));
 sg13g2_a21oi_1 _25731_ (.A1(net5709),
    .A2(net5022),
    .Y(_01546_),
    .B1(_07901_));
 sg13g2_nor2_1 _25732_ (.A(net3351),
    .B(_07898_),
    .Y(_07902_));
 sg13g2_a21oi_1 _25733_ (.A1(net5686),
    .A2(net5023),
    .Y(_01547_),
    .B1(_07902_));
 sg13g2_nor2_1 _25734_ (.A(net3242),
    .B(net5022),
    .Y(_07903_));
 sg13g2_a21oi_1 _25735_ (.A1(net5666),
    .A2(net5022),
    .Y(_01548_),
    .B1(_07903_));
 sg13g2_nor2_1 _25736_ (.A(net4439),
    .B(net5023),
    .Y(_07904_));
 sg13g2_a21oi_1 _25737_ (.A1(net5585),
    .A2(net5023),
    .Y(_01549_),
    .B1(_07904_));
 sg13g2_nor2_1 _25738_ (.A(net3125),
    .B(net5023),
    .Y(_07905_));
 sg13g2_a21oi_1 _25739_ (.A1(net5647),
    .A2(net5023),
    .Y(_01550_),
    .B1(_07905_));
 sg13g2_nor2_1 _25740_ (.A(net3202),
    .B(net5022),
    .Y(_07906_));
 sg13g2_a21oi_1 _25741_ (.A1(net5622),
    .A2(net5022),
    .Y(_01551_),
    .B1(_07906_));
 sg13g2_nor2b_1 _25742_ (.A(\gamepad_pmod.driver.pmod_latch_prev ),
    .B_N(net2928),
    .Y(_07907_));
 sg13g2_nor2_1 _25743_ (.A(net6523),
    .B(net6037),
    .Y(_07908_));
 sg13g2_a22oi_1 _25744_ (.Y(_01552_),
    .B1(net6002),
    .B2(_08640_),
    .A2(net6036),
    .A1(_08486_));
 sg13g2_a22oi_1 _25745_ (.Y(_01553_),
    .B1(net6002),
    .B2(_08641_),
    .A2(net6036),
    .A1(_08485_));
 sg13g2_a22oi_1 _25746_ (.Y(_01554_),
    .B1(net6002),
    .B2(_08643_),
    .A2(net6036),
    .A1(_08484_));
 sg13g2_a22oi_1 _25747_ (.Y(_01555_),
    .B1(net6002),
    .B2(_08642_),
    .A2(net6036),
    .A1(_08483_));
 sg13g2_a22oi_1 _25748_ (.Y(_01556_),
    .B1(net6002),
    .B2(_08644_),
    .A2(net6036),
    .A1(_08482_));
 sg13g2_a22oi_1 _25749_ (.Y(_01557_),
    .B1(net6002),
    .B2(_08645_),
    .A2(net6036),
    .A1(_08481_));
 sg13g2_a22oi_1 _25750_ (.Y(_01558_),
    .B1(net6002),
    .B2(_08646_),
    .A2(net6036),
    .A1(_08480_));
 sg13g2_a22oi_1 _25751_ (.Y(_01559_),
    .B1(net6003),
    .B2(_08647_),
    .A2(net6037),
    .A1(_08479_));
 sg13g2_a22oi_1 _25752_ (.Y(_01560_),
    .B1(net6003),
    .B2(_08648_),
    .A2(net6037),
    .A1(_08478_));
 sg13g2_a22oi_1 _25753_ (.Y(_01561_),
    .B1(net6003),
    .B2(_08649_),
    .A2(net6037),
    .A1(_08477_));
 sg13g2_a22oi_1 _25754_ (.Y(_01562_),
    .B1(net6003),
    .B2(_08650_),
    .A2(net6037),
    .A1(_08476_));
 sg13g2_a22oi_1 _25755_ (.Y(_01563_),
    .B1(net6002),
    .B2(_08651_),
    .A2(net6036),
    .A1(_08475_));
 sg13g2_nand3_1 _25756_ (.B(_09321_),
    .C(net5251),
    .A(net5555),
    .Y(_07909_));
 sg13g2_mux2_1 _25757_ (.A0(net5742),
    .A1(net4655),
    .S(_07909_),
    .X(_01564_));
 sg13g2_mux2_1 _25758_ (.A0(net5744),
    .A1(net4831),
    .S(_07909_),
    .X(_01565_));
 sg13g2_mux2_1 _25759_ (.A0(net5618),
    .A1(net7023),
    .S(_07909_),
    .X(_01566_));
 sg13g2_mux2_1 _25760_ (.A0(net5612),
    .A1(net4784),
    .S(_07909_),
    .X(_01567_));
 sg13g2_mux2_1 _25761_ (.A0(net5606),
    .A1(net6962),
    .S(_07909_),
    .X(_01568_));
 sg13g2_mux2_1 _25762_ (.A0(net5581),
    .A1(net6596),
    .S(_07909_),
    .X(_01569_));
 sg13g2_mux2_1 _25763_ (.A0(net5578),
    .A1(net6585),
    .S(_07909_),
    .X(_01570_));
 sg13g2_mux2_1 _25764_ (.A0(net5644),
    .A1(net4647),
    .S(_07909_),
    .X(_01571_));
 sg13g2_nand3_1 _25765_ (.B(_09321_),
    .C(net5252),
    .A(net5555),
    .Y(_07910_));
 sg13g2_mux2_1 _25766_ (.A0(net5739),
    .A1(net6642),
    .S(_07910_),
    .X(_01572_));
 sg13g2_mux2_1 _25767_ (.A0(net5744),
    .A1(net6930),
    .S(_07910_),
    .X(_01573_));
 sg13g2_mux2_1 _25768_ (.A0(net5618),
    .A1(net4662),
    .S(_07910_),
    .X(_01574_));
 sg13g2_mux2_1 _25769_ (.A0(net5612),
    .A1(net4847),
    .S(_07910_),
    .X(_01575_));
 sg13g2_mux2_1 _25770_ (.A0(net5606),
    .A1(net6743),
    .S(_07910_),
    .X(_01576_));
 sg13g2_mux2_1 _25771_ (.A0(net5581),
    .A1(net4940),
    .S(_07910_),
    .X(_01577_));
 sg13g2_mux2_1 _25772_ (.A0(net5578),
    .A1(net4906),
    .S(_07910_),
    .X(_01578_));
 sg13g2_mux2_1 _25773_ (.A0(net5644),
    .A1(net6601),
    .S(_07910_),
    .X(_01579_));
 sg13g2_nor2_1 _25774_ (.A(_09422_),
    .B(net5238),
    .Y(_07911_));
 sg13g2_nor2_1 _25775_ (.A(net3604),
    .B(net5020),
    .Y(_07912_));
 sg13g2_a21oi_1 _25776_ (.A1(net5759),
    .A2(net5020),
    .Y(_01580_),
    .B1(_07912_));
 sg13g2_nor2_1 _25777_ (.A(net3178),
    .B(net5021),
    .Y(_07913_));
 sg13g2_a21oi_1 _25778_ (.A1(net5780),
    .A2(net5021),
    .Y(_01581_),
    .B1(_07913_));
 sg13g2_nor2_1 _25779_ (.A(net3229),
    .B(net5020),
    .Y(_07914_));
 sg13g2_a21oi_1 _25780_ (.A1(net5709),
    .A2(net5020),
    .Y(_01582_),
    .B1(_07914_));
 sg13g2_nor2_1 _25781_ (.A(net3313),
    .B(_07911_),
    .Y(_07915_));
 sg13g2_a21oi_1 _25782_ (.A1(net5686),
    .A2(net5021),
    .Y(_01583_),
    .B1(_07915_));
 sg13g2_nor2_1 _25783_ (.A(net4556),
    .B(net5020),
    .Y(_07916_));
 sg13g2_a21oi_1 _25784_ (.A1(net5666),
    .A2(net5020),
    .Y(_01584_),
    .B1(_07916_));
 sg13g2_nor2_1 _25785_ (.A(net3347),
    .B(net5021),
    .Y(_07917_));
 sg13g2_a21oi_1 _25786_ (.A1(net5585),
    .A2(net5021),
    .Y(_01585_),
    .B1(_07917_));
 sg13g2_nor2_1 _25787_ (.A(net4400),
    .B(net5020),
    .Y(_07918_));
 sg13g2_a21oi_1 _25788_ (.A1(net5649),
    .A2(net5020),
    .Y(_01586_),
    .B1(_07918_));
 sg13g2_nor2_1 _25789_ (.A(net4292),
    .B(net5021),
    .Y(_07919_));
 sg13g2_a21oi_1 _25790_ (.A1(net5622),
    .A2(net5021),
    .Y(_01587_),
    .B1(_07919_));
 sg13g2_nor3_2 _25791_ (.A(_09053_),
    .B(_09057_),
    .C(_05128_),
    .Y(_07920_));
 sg13g2_mux2_1 _25792_ (.A0(net4419),
    .A1(_05132_),
    .S(_07920_),
    .X(_01588_));
 sg13g2_mux2_1 _25793_ (.A0(net3716),
    .A1(_05139_),
    .S(_07920_),
    .X(_01589_));
 sg13g2_mux2_1 _25794_ (.A0(net3243),
    .A1(_05146_),
    .S(_07920_),
    .X(_01590_));
 sg13g2_mux2_1 _25795_ (.A0(net3638),
    .A1(_05151_),
    .S(_07920_),
    .X(_01591_));
 sg13g2_mux2_1 _25796_ (.A0(net3894),
    .A1(_05153_),
    .S(_07920_),
    .X(_01592_));
 sg13g2_mux2_1 _25797_ (.A0(net3465),
    .A1(_05159_),
    .S(_07920_),
    .X(_01593_));
 sg13g2_mux2_1 _25798_ (.A0(net3652),
    .A1(_05166_),
    .S(_07920_),
    .X(_01594_));
 sg13g2_mux2_1 _25799_ (.A0(net3383),
    .A1(_05171_),
    .S(_07920_),
    .X(_01595_));
 sg13g2_and2_2 _25800_ (.A(_09062_),
    .B(_05129_),
    .X(_07921_));
 sg13g2_mux2_1 _25801_ (.A0(net3672),
    .A1(_05132_),
    .S(_07921_),
    .X(_01596_));
 sg13g2_mux2_1 _25802_ (.A0(net3827),
    .A1(_05139_),
    .S(_07921_),
    .X(_01597_));
 sg13g2_mux2_1 _25803_ (.A0(net4228),
    .A1(_05146_),
    .S(_07921_),
    .X(_01598_));
 sg13g2_mux2_1 _25804_ (.A0(net3337),
    .A1(_05151_),
    .S(_07921_),
    .X(_01599_));
 sg13g2_mux2_1 _25805_ (.A0(net3437),
    .A1(_05153_),
    .S(_07921_),
    .X(_01600_));
 sg13g2_mux2_1 _25806_ (.A0(net3629),
    .A1(_05159_),
    .S(_07921_),
    .X(_01601_));
 sg13g2_mux2_1 _25807_ (.A0(net4342),
    .A1(_05166_),
    .S(_07921_),
    .X(_01602_));
 sg13g2_mux2_1 _25808_ (.A0(net3964),
    .A1(_05171_),
    .S(_07921_),
    .X(_01603_));
 sg13g2_nor2_1 _25809_ (.A(net5263),
    .B(net5257),
    .Y(_07922_));
 sg13g2_nor2_1 _25810_ (.A(net3237),
    .B(net5204),
    .Y(_07923_));
 sg13g2_a21oi_1 _25811_ (.A1(net5764),
    .A2(net5204),
    .Y(_01604_),
    .B1(_07923_));
 sg13g2_nor2_1 _25812_ (.A(net4146),
    .B(net5205),
    .Y(_07924_));
 sg13g2_a21oi_1 _25813_ (.A1(net5786),
    .A2(net5205),
    .Y(_01605_),
    .B1(_07924_));
 sg13g2_nor2_1 _25814_ (.A(net4364),
    .B(net5205),
    .Y(_07925_));
 sg13g2_a21oi_1 _25815_ (.A1(net5714),
    .A2(net5205),
    .Y(_01606_),
    .B1(_07925_));
 sg13g2_nor2_1 _25816_ (.A(net3988),
    .B(net5205),
    .Y(_07926_));
 sg13g2_a21oi_1 _25817_ (.A1(net5687),
    .A2(net5205),
    .Y(_01607_),
    .B1(_07926_));
 sg13g2_nor2_1 _25818_ (.A(net4227),
    .B(net5204),
    .Y(_07927_));
 sg13g2_a21oi_1 _25819_ (.A1(net5671),
    .A2(net5204),
    .Y(_01608_),
    .B1(_07927_));
 sg13g2_nor2_1 _25820_ (.A(net4368),
    .B(net5204),
    .Y(_07928_));
 sg13g2_a21oi_1 _25821_ (.A1(net5586),
    .A2(net5204),
    .Y(_01609_),
    .B1(_07928_));
 sg13g2_nor2_1 _25822_ (.A(net4313),
    .B(_07922_),
    .Y(_07929_));
 sg13g2_a21oi_1 _25823_ (.A1(net5654),
    .A2(net5205),
    .Y(_01610_),
    .B1(_07929_));
 sg13g2_nor2_1 _25824_ (.A(net3404),
    .B(net5204),
    .Y(_07930_));
 sg13g2_a21oi_1 _25825_ (.A1(net5623),
    .A2(net5204),
    .Y(_01611_),
    .B1(_07930_));
 sg13g2_nand2b_2 _25826_ (.Y(_07931_),
    .B(net5252),
    .A_N(net5263));
 sg13g2_mux2_1 _25827_ (.A0(net5739),
    .A1(net4879),
    .S(_07931_),
    .X(_01612_));
 sg13g2_mux2_1 _25828_ (.A0(net5744),
    .A1(net4770),
    .S(_07931_),
    .X(_01613_));
 sg13g2_mux2_1 _25829_ (.A0(net5616),
    .A1(net6655),
    .S(_07931_),
    .X(_01614_));
 sg13g2_mux2_1 _25830_ (.A0(net5611),
    .A1(net7050),
    .S(_07931_),
    .X(_01615_));
 sg13g2_mux2_1 _25831_ (.A0(net5606),
    .A1(net4722),
    .S(_07931_),
    .X(_01616_));
 sg13g2_mux2_1 _25832_ (.A0(net5580),
    .A1(net4497),
    .S(_07931_),
    .X(_01617_));
 sg13g2_mux2_1 _25833_ (.A0(net5576),
    .A1(net7057),
    .S(_07931_),
    .X(_01618_));
 sg13g2_mux2_1 _25834_ (.A0(net5642),
    .A1(net6712),
    .S(_07931_),
    .X(_01619_));
 sg13g2_nor2_1 _25835_ (.A(_09432_),
    .B(net5249),
    .Y(_07932_));
 sg13g2_nor2_1 _25836_ (.A(net3514),
    .B(_07932_),
    .Y(_07933_));
 sg13g2_a21oi_1 _25837_ (.A1(net5764),
    .A2(net5101),
    .Y(_01620_),
    .B1(_07933_));
 sg13g2_nor2_1 _25838_ (.A(net3311),
    .B(net5101),
    .Y(_07934_));
 sg13g2_a21oi_1 _25839_ (.A1(net5785),
    .A2(net5101),
    .Y(_01621_),
    .B1(_07934_));
 sg13g2_nor2_1 _25840_ (.A(net3077),
    .B(net5101),
    .Y(_07935_));
 sg13g2_a21oi_1 _25841_ (.A1(net5717),
    .A2(net5102),
    .Y(_01622_),
    .B1(_07935_));
 sg13g2_nor2_1 _25842_ (.A(net3973),
    .B(net5101),
    .Y(_07936_));
 sg13g2_a21oi_1 _25843_ (.A1(net5688),
    .A2(net5101),
    .Y(_01623_),
    .B1(_07936_));
 sg13g2_nor2_1 _25844_ (.A(net3593),
    .B(net5102),
    .Y(_07937_));
 sg13g2_a21oi_1 _25845_ (.A1(net5667),
    .A2(net5102),
    .Y(_01624_),
    .B1(_07937_));
 sg13g2_nor2_1 _25846_ (.A(net3177),
    .B(net5102),
    .Y(_07938_));
 sg13g2_a21oi_1 _25847_ (.A1(net5587),
    .A2(net5102),
    .Y(_01625_),
    .B1(_07938_));
 sg13g2_nor2_1 _25848_ (.A(net3260),
    .B(net5101),
    .Y(_07939_));
 sg13g2_a21oi_1 _25849_ (.A1(net5654),
    .A2(net5101),
    .Y(_01626_),
    .B1(_07939_));
 sg13g2_nor2_1 _25850_ (.A(net3597),
    .B(net5102),
    .Y(_07940_));
 sg13g2_a21oi_1 _25851_ (.A1(net5624),
    .A2(net5102),
    .Y(_01627_),
    .B1(_07940_));
 sg13g2_nor2_1 _25852_ (.A(_09432_),
    .B(net5237),
    .Y(_07941_));
 sg13g2_nor2_1 _25853_ (.A(net4031),
    .B(_07941_),
    .Y(_07942_));
 sg13g2_a21oi_1 _25854_ (.A1(net5764),
    .A2(net5099),
    .Y(_01628_),
    .B1(_07942_));
 sg13g2_nor2_1 _25855_ (.A(net3247),
    .B(net5099),
    .Y(_07943_));
 sg13g2_a21oi_1 _25856_ (.A1(net5785),
    .A2(net5100),
    .Y(_01629_),
    .B1(_07943_));
 sg13g2_nor2_1 _25857_ (.A(net3164),
    .B(net5099),
    .Y(_07944_));
 sg13g2_a21oi_1 _25858_ (.A1(net5714),
    .A2(net5099),
    .Y(_01630_),
    .B1(_07944_));
 sg13g2_nor2_1 _25859_ (.A(net3163),
    .B(net5099),
    .Y(_07945_));
 sg13g2_a21oi_1 _25860_ (.A1(net5688),
    .A2(net5099),
    .Y(_01631_),
    .B1(_07945_));
 sg13g2_nor2_1 _25861_ (.A(net3297),
    .B(net5100),
    .Y(_07946_));
 sg13g2_a21oi_1 _25862_ (.A1(net5667),
    .A2(net5100),
    .Y(_01632_),
    .B1(_07946_));
 sg13g2_nor2_1 _25863_ (.A(net3080),
    .B(net5100),
    .Y(_07947_));
 sg13g2_a21oi_1 _25864_ (.A1(net5587),
    .A2(net5100),
    .Y(_01633_),
    .B1(_07947_));
 sg13g2_nor2_1 _25865_ (.A(net3068),
    .B(net5099),
    .Y(_07948_));
 sg13g2_a21oi_1 _25866_ (.A1(net5654),
    .A2(net5099),
    .Y(_01634_),
    .B1(_07948_));
 sg13g2_nor2_1 _25867_ (.A(net3362),
    .B(net5100),
    .Y(_07949_));
 sg13g2_a21oi_1 _25868_ (.A1(net5624),
    .A2(net5100),
    .Y(_01635_),
    .B1(_07949_));
 sg13g2_nor2_1 _25869_ (.A(_09432_),
    .B(net5259),
    .Y(_07950_));
 sg13g2_nor2_1 _25870_ (.A(net4397),
    .B(net5098),
    .Y(_07951_));
 sg13g2_a21oi_1 _25871_ (.A1(net5767),
    .A2(net5098),
    .Y(_01636_),
    .B1(_07951_));
 sg13g2_nor2_1 _25872_ (.A(net3963),
    .B(_07950_),
    .Y(_07952_));
 sg13g2_a21oi_1 _25873_ (.A1(net5785),
    .A2(net5098),
    .Y(_01637_),
    .B1(_07952_));
 sg13g2_nor2_1 _25874_ (.A(net3758),
    .B(net5098),
    .Y(_07953_));
 sg13g2_a21oi_1 _25875_ (.A1(net5714),
    .A2(net5098),
    .Y(_01638_),
    .B1(_07953_));
 sg13g2_nor2_1 _25876_ (.A(net4486),
    .B(net5097),
    .Y(_07954_));
 sg13g2_a21oi_1 _25877_ (.A1(net5688),
    .A2(net5097),
    .Y(_01639_),
    .B1(_07954_));
 sg13g2_nor2_1 _25878_ (.A(net3291),
    .B(net5097),
    .Y(_07955_));
 sg13g2_a21oi_1 _25879_ (.A1(net5672),
    .A2(net5097),
    .Y(_01640_),
    .B1(_07955_));
 sg13g2_nor2_1 _25880_ (.A(net4009),
    .B(net5097),
    .Y(_07956_));
 sg13g2_a21oi_1 _25881_ (.A1(net5587),
    .A2(net5097),
    .Y(_01641_),
    .B1(_07956_));
 sg13g2_nor2_1 _25882_ (.A(net3446),
    .B(net5098),
    .Y(_07957_));
 sg13g2_a21oi_1 _25883_ (.A1(net5654),
    .A2(net5098),
    .Y(_01642_),
    .B1(_07957_));
 sg13g2_nor2_1 _25884_ (.A(net3761),
    .B(net5097),
    .Y(_07958_));
 sg13g2_a21oi_1 _25885_ (.A1(net5627),
    .A2(net5097),
    .Y(_01643_),
    .B1(_07958_));
 sg13g2_nor2_1 _25886_ (.A(net5203),
    .B(net5255),
    .Y(_07959_));
 sg13g2_nor2_1 _25887_ (.A(net3982),
    .B(net5019),
    .Y(_07960_));
 sg13g2_a21oi_1 _25888_ (.A1(net5762),
    .A2(net5019),
    .Y(_01644_),
    .B1(_07960_));
 sg13g2_nor2_1 _25889_ (.A(net3026),
    .B(net5019),
    .Y(_07961_));
 sg13g2_a21oi_1 _25890_ (.A1(net5783),
    .A2(net5019),
    .Y(_01645_),
    .B1(_07961_));
 sg13g2_nor2_1 _25891_ (.A(net3775),
    .B(net5019),
    .Y(_07962_));
 sg13g2_a21oi_1 _25892_ (.A1(net5713),
    .A2(net5019),
    .Y(_01646_),
    .B1(_07962_));
 sg13g2_nor2_1 _25893_ (.A(net3671),
    .B(net5018),
    .Y(_07963_));
 sg13g2_a21oi_1 _25894_ (.A1(net5691),
    .A2(net5018),
    .Y(_01647_),
    .B1(_07963_));
 sg13g2_nor2_1 _25895_ (.A(net3025),
    .B(net5019),
    .Y(_07964_));
 sg13g2_a21oi_1 _25896_ (.A1(net5668),
    .A2(net5019),
    .Y(_01648_),
    .B1(_07964_));
 sg13g2_nor2_1 _25897_ (.A(net3706),
    .B(net5018),
    .Y(_07965_));
 sg13g2_a21oi_1 _25898_ (.A1(net5592),
    .A2(net5018),
    .Y(_01649_),
    .B1(_07965_));
 sg13g2_nor2_1 _25899_ (.A(net3798),
    .B(net5018),
    .Y(_07966_));
 sg13g2_a21oi_1 _25900_ (.A1(net5651),
    .A2(net5018),
    .Y(_01650_),
    .B1(_07966_));
 sg13g2_nor2_1 _25901_ (.A(net4340),
    .B(net5018),
    .Y(_07967_));
 sg13g2_a21oi_1 _25902_ (.A1(net5629),
    .A2(net5018),
    .Y(_01651_),
    .B1(_07967_));
 sg13g2_nor2_1 _25903_ (.A(_09432_),
    .B(net5238),
    .Y(_07968_));
 sg13g2_nor2_1 _25904_ (.A(net4299),
    .B(net5096),
    .Y(_07969_));
 sg13g2_a21oi_1 _25905_ (.A1(net5764),
    .A2(net5096),
    .Y(_01652_),
    .B1(_07969_));
 sg13g2_nor2_1 _25906_ (.A(net3029),
    .B(net5096),
    .Y(_07970_));
 sg13g2_a21oi_1 _25907_ (.A1(net5785),
    .A2(net5096),
    .Y(_01653_),
    .B1(_07970_));
 sg13g2_nor2_1 _25908_ (.A(net3887),
    .B(net5096),
    .Y(_07971_));
 sg13g2_a21oi_1 _25909_ (.A1(net5717),
    .A2(net5096),
    .Y(_01654_),
    .B1(_07971_));
 sg13g2_nor2_1 _25910_ (.A(net3253),
    .B(net5095),
    .Y(_07972_));
 sg13g2_a21oi_1 _25911_ (.A1(net5694),
    .A2(net5095),
    .Y(_01655_),
    .B1(_07972_));
 sg13g2_nor2_1 _25912_ (.A(net3487),
    .B(net5095),
    .Y(_07973_));
 sg13g2_a21oi_1 _25913_ (.A1(net5672),
    .A2(net5095),
    .Y(_01656_),
    .B1(_07973_));
 sg13g2_nor2_1 _25914_ (.A(net4161),
    .B(net5095),
    .Y(_07974_));
 sg13g2_a21oi_1 _25915_ (.A1(net5590),
    .A2(net5095),
    .Y(_01657_),
    .B1(_07974_));
 sg13g2_nor2_1 _25916_ (.A(net3885),
    .B(net5095),
    .Y(_07975_));
 sg13g2_a21oi_1 _25917_ (.A1(net5654),
    .A2(net5095),
    .Y(_01658_),
    .B1(_07975_));
 sg13g2_nor2_1 _25918_ (.A(net3367),
    .B(net5096),
    .Y(_07976_));
 sg13g2_a21oi_1 _25919_ (.A1(net5628),
    .A2(net5096),
    .Y(_01659_),
    .B1(_07976_));
 sg13g2_nor2_1 _25920_ (.A(_09432_),
    .B(net5255),
    .Y(_07977_));
 sg13g2_nor2_1 _25921_ (.A(net4116),
    .B(net5094),
    .Y(_07978_));
 sg13g2_a21oi_1 _25922_ (.A1(net5764),
    .A2(_07977_),
    .Y(_01660_),
    .B1(_07978_));
 sg13g2_nor2_1 _25923_ (.A(net3327),
    .B(net5093),
    .Y(_07979_));
 sg13g2_a21oi_1 _25924_ (.A1(net5784),
    .A2(net5093),
    .Y(_01661_),
    .B1(_07979_));
 sg13g2_nor2_1 _25925_ (.A(net4109),
    .B(net5093),
    .Y(_07980_));
 sg13g2_a21oi_1 _25926_ (.A1(net5714),
    .A2(net5093),
    .Y(_01662_),
    .B1(_07980_));
 sg13g2_nor2_1 _25927_ (.A(net3036),
    .B(net5094),
    .Y(_07981_));
 sg13g2_a21oi_1 _25928_ (.A1(net5694),
    .A2(net5094),
    .Y(_01663_),
    .B1(_07981_));
 sg13g2_nor2_1 _25929_ (.A(net3381),
    .B(net5093),
    .Y(_07982_));
 sg13g2_a21oi_1 _25930_ (.A1(net5671),
    .A2(net5093),
    .Y(_01664_),
    .B1(_07982_));
 sg13g2_nor2_1 _25931_ (.A(net3782),
    .B(net5094),
    .Y(_07983_));
 sg13g2_a21oi_1 _25932_ (.A1(net5590),
    .A2(net5094),
    .Y(_01665_),
    .B1(_07983_));
 sg13g2_nor2_1 _25933_ (.A(net3722),
    .B(net5093),
    .Y(_07984_));
 sg13g2_a21oi_1 _25934_ (.A1(net5652),
    .A2(net5093),
    .Y(_01666_),
    .B1(_07984_));
 sg13g2_nor2_1 _25935_ (.A(net3244),
    .B(net5094),
    .Y(_07985_));
 sg13g2_a21oi_1 _25936_ (.A1(net5626),
    .A2(net5094),
    .Y(_01667_),
    .B1(_07985_));
 sg13g2_nor2_1 _25937_ (.A(_09432_),
    .B(net5257),
    .Y(_07986_));
 sg13g2_nor2_1 _25938_ (.A(net3315),
    .B(net5092),
    .Y(_07987_));
 sg13g2_a21oi_1 _25939_ (.A1(net5764),
    .A2(net5092),
    .Y(_01668_),
    .B1(_07987_));
 sg13g2_nor2_1 _25940_ (.A(net3180),
    .B(net5092),
    .Y(_07988_));
 sg13g2_a21oi_1 _25941_ (.A1(net5784),
    .A2(net5092),
    .Y(_01669_),
    .B1(_07988_));
 sg13g2_nor2_1 _25942_ (.A(net4065),
    .B(net5092),
    .Y(_07989_));
 sg13g2_a21oi_1 _25943_ (.A1(net5714),
    .A2(net5092),
    .Y(_01670_),
    .B1(_07989_));
 sg13g2_nor2_1 _25944_ (.A(net4101),
    .B(net5091),
    .Y(_07990_));
 sg13g2_a21oi_1 _25945_ (.A1(net5694),
    .A2(net5091),
    .Y(_01671_),
    .B1(_07990_));
 sg13g2_nor2_1 _25946_ (.A(net3912),
    .B(net5091),
    .Y(_07991_));
 sg13g2_a21oi_1 _25947_ (.A1(net5673),
    .A2(net5091),
    .Y(_01672_),
    .B1(_07991_));
 sg13g2_nor2_1 _25948_ (.A(net3433),
    .B(net5091),
    .Y(_07992_));
 sg13g2_a21oi_1 _25949_ (.A1(net5590),
    .A2(net5091),
    .Y(_01673_),
    .B1(_07992_));
 sg13g2_nor2_1 _25950_ (.A(net3688),
    .B(net5092),
    .Y(_07993_));
 sg13g2_a21oi_1 _25951_ (.A1(net5652),
    .A2(net5092),
    .Y(_01674_),
    .B1(_07993_));
 sg13g2_nor2_1 _25952_ (.A(net3082),
    .B(net5091),
    .Y(_07994_));
 sg13g2_a21oi_1 _25953_ (.A1(net5626),
    .A2(net5091),
    .Y(_01675_),
    .B1(_07994_));
 sg13g2_nand3_1 _25954_ (.B(_09318_),
    .C(net5252),
    .A(_09262_),
    .Y(_07995_));
 sg13g2_mux2_1 _25955_ (.A0(net5739),
    .A1(net4833),
    .S(_07995_),
    .X(_01676_));
 sg13g2_mux2_1 _25956_ (.A0(net5744),
    .A1(net6894),
    .S(_07995_),
    .X(_01677_));
 sg13g2_mux2_1 _25957_ (.A0(net5616),
    .A1(net6589),
    .S(_07995_),
    .X(_01678_));
 sg13g2_mux2_1 _25958_ (.A0(net5611),
    .A1(net4952),
    .S(_07995_),
    .X(_01679_));
 sg13g2_mux2_1 _25959_ (.A0(net5606),
    .A1(net4718),
    .S(_07995_),
    .X(_01680_));
 sg13g2_mux2_1 _25960_ (.A0(net5581),
    .A1(net4898),
    .S(_07995_),
    .X(_01681_));
 sg13g2_mux2_1 _25961_ (.A0(net5576),
    .A1(net6694),
    .S(_07995_),
    .X(_01682_));
 sg13g2_mux2_1 _25962_ (.A0(net5642),
    .A1(net4649),
    .S(_07995_),
    .X(_01683_));
 sg13g2_nor2_1 _25963_ (.A(_03124_),
    .B(net5248),
    .Y(_07996_));
 sg13g2_nor2_1 _25964_ (.A(net3267),
    .B(net5089),
    .Y(_07997_));
 sg13g2_a21oi_1 _25965_ (.A1(net5775),
    .A2(net5089),
    .Y(_01684_),
    .B1(_07997_));
 sg13g2_nor2_1 _25966_ (.A(net3585),
    .B(net5090),
    .Y(_07998_));
 sg13g2_a21oi_1 _25967_ (.A1(net5792),
    .A2(net5090),
    .Y(_01685_),
    .B1(_07998_));
 sg13g2_nor2_1 _25968_ (.A(net4108),
    .B(net5090),
    .Y(_07999_));
 sg13g2_a21oi_1 _25969_ (.A1(net5722),
    .A2(net5090),
    .Y(_01686_),
    .B1(_07999_));
 sg13g2_nor2_1 _25970_ (.A(net3314),
    .B(net5090),
    .Y(_08000_));
 sg13g2_a21oi_1 _25971_ (.A1(net5701),
    .A2(net5090),
    .Y(_01687_),
    .B1(_08000_));
 sg13g2_nor2_1 _25972_ (.A(net3158),
    .B(net5089),
    .Y(_08001_));
 sg13g2_a21oi_1 _25973_ (.A1(net5680),
    .A2(net5089),
    .Y(_01688_),
    .B1(_08001_));
 sg13g2_nor2_1 _25974_ (.A(net4230),
    .B(net5089),
    .Y(_08002_));
 sg13g2_a21oi_1 _25975_ (.A1(net5602),
    .A2(net5089),
    .Y(_01689_),
    .B1(_08002_));
 sg13g2_nor2_1 _25976_ (.A(net3938),
    .B(net5090),
    .Y(_08003_));
 sg13g2_a21oi_1 _25977_ (.A1(net5661),
    .A2(_07996_),
    .Y(_01690_),
    .B1(_08003_));
 sg13g2_nor2_1 _25978_ (.A(net7058),
    .B(net5089),
    .Y(_08004_));
 sg13g2_a21oi_1 _25979_ (.A1(net5638),
    .A2(net5089),
    .Y(_01691_),
    .B1(_08004_));
 sg13g2_nor2_1 _25980_ (.A(_03124_),
    .B(net5236),
    .Y(_08005_));
 sg13g2_nor2_1 _25981_ (.A(net4038),
    .B(net5087),
    .Y(_08006_));
 sg13g2_a21oi_1 _25982_ (.A1(net5775),
    .A2(net5087),
    .Y(_01692_),
    .B1(_08006_));
 sg13g2_nor2_1 _25983_ (.A(net4168),
    .B(net5088),
    .Y(_08007_));
 sg13g2_a21oi_1 _25984_ (.A1(net5792),
    .A2(net5088),
    .Y(_01693_),
    .B1(_08007_));
 sg13g2_nor2_1 _25985_ (.A(net3309),
    .B(net5088),
    .Y(_08008_));
 sg13g2_a21oi_1 _25986_ (.A1(net5722),
    .A2(net5088),
    .Y(_01694_),
    .B1(_08008_));
 sg13g2_nor2_1 _25987_ (.A(net4029),
    .B(net5088),
    .Y(_08009_));
 sg13g2_a21oi_1 _25988_ (.A1(net5702),
    .A2(net5088),
    .Y(_01695_),
    .B1(_08009_));
 sg13g2_nor2_1 _25989_ (.A(net3608),
    .B(_08005_),
    .Y(_08010_));
 sg13g2_a21oi_1 _25990_ (.A1(net5680),
    .A2(net5088),
    .Y(_01696_),
    .B1(_08010_));
 sg13g2_nor2_1 _25991_ (.A(net3220),
    .B(net5087),
    .Y(_08011_));
 sg13g2_a21oi_1 _25992_ (.A1(net5602),
    .A2(net5087),
    .Y(_01697_),
    .B1(_08011_));
 sg13g2_nor2_1 _25993_ (.A(net3123),
    .B(net5087),
    .Y(_08012_));
 sg13g2_a21oi_1 _25994_ (.A1(net5662),
    .A2(net5087),
    .Y(_01698_),
    .B1(_08012_));
 sg13g2_nor2_1 _25995_ (.A(net3141),
    .B(net5087),
    .Y(_08013_));
 sg13g2_a21oi_1 _25996_ (.A1(net5633),
    .A2(net5087),
    .Y(_01699_),
    .B1(_08013_));
 sg13g2_nor2_1 _25997_ (.A(net5258),
    .B(_03124_),
    .Y(_08014_));
 sg13g2_nor2_1 _25998_ (.A(net3485),
    .B(net5086),
    .Y(_08015_));
 sg13g2_a21oi_1 _25999_ (.A1(net5775),
    .A2(net5086),
    .Y(_01700_),
    .B1(_08015_));
 sg13g2_nor2_1 _26000_ (.A(net4200),
    .B(net5086),
    .Y(_08016_));
 sg13g2_a21oi_1 _26001_ (.A1(net5792),
    .A2(net5085),
    .Y(_01701_),
    .B1(_08016_));
 sg13g2_nor2_1 _26002_ (.A(net3956),
    .B(net5085),
    .Y(_08017_));
 sg13g2_a21oi_1 _26003_ (.A1(net5722),
    .A2(net5085),
    .Y(_01702_),
    .B1(_08017_));
 sg13g2_nor2_1 _26004_ (.A(net3754),
    .B(net5085),
    .Y(_08018_));
 sg13g2_a21oi_1 _26005_ (.A1(net5702),
    .A2(net5085),
    .Y(_01703_),
    .B1(_08018_));
 sg13g2_nor2_1 _26006_ (.A(net4367),
    .B(net5086),
    .Y(_08019_));
 sg13g2_a21oi_1 _26007_ (.A1(net5680),
    .A2(net5085),
    .Y(_01704_),
    .B1(_08019_));
 sg13g2_nor2_1 _26008_ (.A(net3219),
    .B(_08014_),
    .Y(_08020_));
 sg13g2_a21oi_1 _26009_ (.A1(net5602),
    .A2(net5086),
    .Y(_01705_),
    .B1(_08020_));
 sg13g2_nor2_1 _26010_ (.A(net3281),
    .B(net5086),
    .Y(_08021_));
 sg13g2_a21oi_1 _26011_ (.A1(net5662),
    .A2(net5086),
    .Y(_01706_),
    .B1(_08021_));
 sg13g2_nor2_1 _26012_ (.A(net4175),
    .B(net5085),
    .Y(_08022_));
 sg13g2_a21oi_1 _26013_ (.A1(net5633),
    .A2(net5085),
    .Y(_01707_),
    .B1(_08022_));
 sg13g2_nand3_1 _26014_ (.B(_03122_),
    .C(net5251),
    .A(_09105_),
    .Y(_08023_));
 sg13g2_mux2_1 _26015_ (.A0(net5743),
    .A1(net6586),
    .S(_08023_),
    .X(_01708_));
 sg13g2_mux2_1 _26016_ (.A0(net5746),
    .A1(net6673),
    .S(_08023_),
    .X(_01709_));
 sg13g2_mux2_1 _26017_ (.A0(net5618),
    .A1(net7189),
    .S(_08023_),
    .X(_01710_));
 sg13g2_mux2_1 _26018_ (.A0(net5612),
    .A1(net6608),
    .S(_08023_),
    .X(_01711_));
 sg13g2_mux2_1 _26019_ (.A0(net5609),
    .A1(net4551),
    .S(_08023_),
    .X(_01712_));
 sg13g2_mux2_1 _26020_ (.A0(net5584),
    .A1(net6987),
    .S(_08023_),
    .X(_01713_));
 sg13g2_mux2_1 _26021_ (.A0(net5577),
    .A1(net6981),
    .S(_08023_),
    .X(_01714_));
 sg13g2_mux2_1 _26022_ (.A0(net5643),
    .A1(net6715),
    .S(_08023_),
    .X(_01715_));
 sg13g2_nor2_1 _26023_ (.A(net5238),
    .B(_03124_),
    .Y(_08024_));
 sg13g2_nor2_1 _26024_ (.A(net3958),
    .B(net5084),
    .Y(_08025_));
 sg13g2_a21oi_1 _26025_ (.A1(net5775),
    .A2(net5084),
    .Y(_01716_),
    .B1(_08025_));
 sg13g2_nor2_1 _26026_ (.A(net3150),
    .B(net5083),
    .Y(_08026_));
 sg13g2_a21oi_1 _26027_ (.A1(net5794),
    .A2(net5083),
    .Y(_01717_),
    .B1(_08026_));
 sg13g2_nor2_1 _26028_ (.A(net3235),
    .B(net5083),
    .Y(_08027_));
 sg13g2_a21oi_1 _26029_ (.A1(net5725),
    .A2(net5083),
    .Y(_01718_),
    .B1(_08027_));
 sg13g2_nor2_1 _26030_ (.A(net4950),
    .B(net5083),
    .Y(_08028_));
 sg13g2_a21oi_1 _26031_ (.A1(net5701),
    .A2(net5083),
    .Y(_01719_),
    .B1(_08028_));
 sg13g2_nor2_1 _26032_ (.A(net3821),
    .B(net5083),
    .Y(_08029_));
 sg13g2_a21oi_1 _26033_ (.A1(net5680),
    .A2(net5083),
    .Y(_01720_),
    .B1(_08029_));
 sg13g2_nor2_1 _26034_ (.A(net3883),
    .B(net5084),
    .Y(_08030_));
 sg13g2_a21oi_1 _26035_ (.A1(net5602),
    .A2(net5084),
    .Y(_01721_),
    .B1(_08030_));
 sg13g2_nor2_1 _26036_ (.A(net4282),
    .B(net5084),
    .Y(_08031_));
 sg13g2_a21oi_1 _26037_ (.A1(net5663),
    .A2(net5084),
    .Y(_01722_),
    .B1(_08031_));
 sg13g2_nor2_1 _26038_ (.A(net4224),
    .B(net5084),
    .Y(_08032_));
 sg13g2_a21oi_1 _26039_ (.A1(net5638),
    .A2(net5084),
    .Y(_01723_),
    .B1(_08032_));
 sg13g2_nor2_1 _26040_ (.A(net5203),
    .B(net5257),
    .Y(_08033_));
 sg13g2_nor2_1 _26041_ (.A(net4242),
    .B(net5017),
    .Y(_08034_));
 sg13g2_a21oi_1 _26042_ (.A1(net5762),
    .A2(net5017),
    .Y(_01724_),
    .B1(_08034_));
 sg13g2_nor2_1 _26043_ (.A(net3301),
    .B(net5017),
    .Y(_08035_));
 sg13g2_a21oi_1 _26044_ (.A1(net5783),
    .A2(net5017),
    .Y(_01725_),
    .B1(_08035_));
 sg13g2_nor2_1 _26045_ (.A(net3792),
    .B(net5017),
    .Y(_08036_));
 sg13g2_a21oi_1 _26046_ (.A1(net5713),
    .A2(net5017),
    .Y(_01726_),
    .B1(_08036_));
 sg13g2_nor2_1 _26047_ (.A(net3864),
    .B(net5016),
    .Y(_08037_));
 sg13g2_a21oi_1 _26048_ (.A1(net5690),
    .A2(net5016),
    .Y(_01727_),
    .B1(_08037_));
 sg13g2_nor2_1 _26049_ (.A(net4395),
    .B(net5017),
    .Y(_08038_));
 sg13g2_a21oi_1 _26050_ (.A1(net5668),
    .A2(net5017),
    .Y(_01728_),
    .B1(_08038_));
 sg13g2_nor2_1 _26051_ (.A(net3959),
    .B(net5016),
    .Y(_08039_));
 sg13g2_a21oi_1 _26052_ (.A1(net5592),
    .A2(net5016),
    .Y(_01729_),
    .B1(_08039_));
 sg13g2_nor2_1 _26053_ (.A(net4212),
    .B(net5016),
    .Y(_08040_));
 sg13g2_a21oi_1 _26054_ (.A1(net5651),
    .A2(net5016),
    .Y(_01730_),
    .B1(_08040_));
 sg13g2_nor2_1 _26055_ (.A(net4154),
    .B(net5016),
    .Y(_08041_));
 sg13g2_a21oi_1 _26056_ (.A1(net5631),
    .A2(net5016),
    .Y(_01731_),
    .B1(_08041_));
 sg13g2_nor2_1 _26057_ (.A(net5256),
    .B(_03124_),
    .Y(_08042_));
 sg13g2_nor2_1 _26058_ (.A(net3249),
    .B(net5081),
    .Y(_08043_));
 sg13g2_a21oi_1 _26059_ (.A1(net5775),
    .A2(net5081),
    .Y(_01732_),
    .B1(_08043_));
 sg13g2_nor2_1 _26060_ (.A(net3290),
    .B(net5082),
    .Y(_08044_));
 sg13g2_a21oi_1 _26061_ (.A1(net5795),
    .A2(net5082),
    .Y(_01733_),
    .B1(_08044_));
 sg13g2_nor2_1 _26062_ (.A(net3113),
    .B(net5082),
    .Y(_08045_));
 sg13g2_a21oi_1 _26063_ (.A1(net5724),
    .A2(net5082),
    .Y(_01734_),
    .B1(_08045_));
 sg13g2_nor2_1 _26064_ (.A(net3557),
    .B(net5082),
    .Y(_08046_));
 sg13g2_a21oi_1 _26065_ (.A1(net5701),
    .A2(net5082),
    .Y(_01735_),
    .B1(_08046_));
 sg13g2_nor2_1 _26066_ (.A(net3529),
    .B(net5081),
    .Y(_08047_));
 sg13g2_a21oi_1 _26067_ (.A1(net5680),
    .A2(net5081),
    .Y(_01736_),
    .B1(_08047_));
 sg13g2_nor2_1 _26068_ (.A(net4462),
    .B(net5081),
    .Y(_08048_));
 sg13g2_a21oi_1 _26069_ (.A1(net5602),
    .A2(net5081),
    .Y(_01737_),
    .B1(_08048_));
 sg13g2_nor2_1 _26070_ (.A(net3692),
    .B(net5081),
    .Y(_08049_));
 sg13g2_a21oi_1 _26071_ (.A1(net5663),
    .A2(net5081),
    .Y(_01738_),
    .B1(_08049_));
 sg13g2_nor2_1 _26072_ (.A(net3346),
    .B(net5082),
    .Y(_08050_));
 sg13g2_a21oi_1 _26073_ (.A1(net5638),
    .A2(_08042_),
    .Y(_01739_),
    .B1(_08050_));
 sg13g2_nor2_1 _26074_ (.A(net5238),
    .B(_03134_),
    .Y(_08051_));
 sg13g2_nor2_1 _26075_ (.A(net3078),
    .B(net5014),
    .Y(_08052_));
 sg13g2_a21oi_1 _26076_ (.A1(net5769),
    .A2(net5014),
    .Y(_01740_),
    .B1(_08052_));
 sg13g2_nor2_1 _26077_ (.A(net3248),
    .B(net5014),
    .Y(_08053_));
 sg13g2_a21oi_1 _26078_ (.A1(net5789),
    .A2(net5014),
    .Y(_01741_),
    .B1(_08053_));
 sg13g2_nor2_1 _26079_ (.A(net3978),
    .B(net5015),
    .Y(_08054_));
 sg13g2_a21oi_1 _26080_ (.A1(net5719),
    .A2(net5015),
    .Y(_01742_),
    .B1(_08054_));
 sg13g2_nor2_1 _26081_ (.A(net3061),
    .B(net5015),
    .Y(_08055_));
 sg13g2_a21oi_1 _26082_ (.A1(net5696),
    .A2(net5015),
    .Y(_01743_),
    .B1(_08055_));
 sg13g2_nor2_1 _26083_ (.A(net3555),
    .B(net5014),
    .Y(_08056_));
 sg13g2_a21oi_1 _26084_ (.A1(net5674),
    .A2(net5014),
    .Y(_01744_),
    .B1(_08056_));
 sg13g2_nor2_1 _26085_ (.A(net3445),
    .B(net5015),
    .Y(_08057_));
 sg13g2_a21oi_1 _26086_ (.A1(net5593),
    .A2(net5015),
    .Y(_01745_),
    .B1(_08057_));
 sg13g2_nor2_1 _26087_ (.A(net3880),
    .B(net5014),
    .Y(_08058_));
 sg13g2_a21oi_1 _26088_ (.A1(net5655),
    .A2(net5014),
    .Y(_01746_),
    .B1(_08058_));
 sg13g2_nor2_1 _26089_ (.A(net3195),
    .B(net5015),
    .Y(_08059_));
 sg13g2_a21oi_1 _26090_ (.A1(net5630),
    .A2(net5015),
    .Y(_01747_),
    .B1(_08059_));
 sg13g2_nor2_1 _26091_ (.A(net5203),
    .B(net5237),
    .Y(_08060_));
 sg13g2_nor2_1 _26092_ (.A(net3088),
    .B(net5013),
    .Y(_08061_));
 sg13g2_a21oi_1 _26093_ (.A1(net5762),
    .A2(net5013),
    .Y(_01748_),
    .B1(_08061_));
 sg13g2_nor2_1 _26094_ (.A(net3961),
    .B(_08060_),
    .Y(_08062_));
 sg13g2_a21oi_1 _26095_ (.A1(net5782),
    .A2(net5013),
    .Y(_01749_),
    .B1(_08062_));
 sg13g2_nor2_1 _26096_ (.A(net3140),
    .B(net5013),
    .Y(_08063_));
 sg13g2_a21oi_1 _26097_ (.A1(net5712),
    .A2(net5012),
    .Y(_01750_),
    .B1(_08063_));
 sg13g2_nor2_1 _26098_ (.A(net3179),
    .B(net5013),
    .Y(_08064_));
 sg13g2_a21oi_1 _26099_ (.A1(net5690),
    .A2(net5012),
    .Y(_01751_),
    .B1(_08064_));
 sg13g2_nor2_1 _26100_ (.A(net3040),
    .B(net5013),
    .Y(_08065_));
 sg13g2_a21oi_1 _26101_ (.A1(net5668),
    .A2(net5013),
    .Y(_01752_),
    .B1(_08065_));
 sg13g2_nor2_1 _26102_ (.A(net3776),
    .B(net5012),
    .Y(_08066_));
 sg13g2_a21oi_1 _26103_ (.A1(net5591),
    .A2(net5012),
    .Y(_01753_),
    .B1(_08066_));
 sg13g2_nor2_1 _26104_ (.A(net4358),
    .B(net5012),
    .Y(_08067_));
 sg13g2_a21oi_1 _26105_ (.A1(net5650),
    .A2(net5012),
    .Y(_01754_),
    .B1(_08067_));
 sg13g2_nor2_1 _26106_ (.A(net4335),
    .B(net5012),
    .Y(_08068_));
 sg13g2_a21oi_1 _26107_ (.A1(net5629),
    .A2(net5012),
    .Y(_01755_),
    .B1(_08068_));
 sg13g2_nor2_1 _26108_ (.A(net5259),
    .B(_03134_),
    .Y(_08069_));
 sg13g2_nor2_1 _26109_ (.A(net3184),
    .B(_08069_),
    .Y(_08070_));
 sg13g2_a21oi_1 _26110_ (.A1(net5769),
    .A2(net5010),
    .Y(_01756_),
    .B1(_08070_));
 sg13g2_nor2_1 _26111_ (.A(net4322),
    .B(net5011),
    .Y(_08071_));
 sg13g2_a21oi_1 _26112_ (.A1(net5789),
    .A2(net5011),
    .Y(_01757_),
    .B1(_08071_));
 sg13g2_nor2_1 _26113_ (.A(net3389),
    .B(net5010),
    .Y(_08072_));
 sg13g2_a21oi_1 _26114_ (.A1(net5719),
    .A2(net5011),
    .Y(_01758_),
    .B1(_08072_));
 sg13g2_nor2_1 _26115_ (.A(net4318),
    .B(net5010),
    .Y(_08073_));
 sg13g2_a21oi_1 _26116_ (.A1(net5696),
    .A2(net5010),
    .Y(_01759_),
    .B1(_08073_));
 sg13g2_nor2_1 _26117_ (.A(net3544),
    .B(net5011),
    .Y(_08074_));
 sg13g2_a21oi_1 _26118_ (.A1(net5674),
    .A2(net5011),
    .Y(_01760_),
    .B1(_08074_));
 sg13g2_nor2_1 _26119_ (.A(net4723),
    .B(net5010),
    .Y(_08075_));
 sg13g2_a21oi_1 _26120_ (.A1(net5594),
    .A2(net5010),
    .Y(_01761_),
    .B1(_08075_));
 sg13g2_nor2_1 _26121_ (.A(net4234),
    .B(net5011),
    .Y(_08076_));
 sg13g2_a21oi_1 _26122_ (.A1(net5655),
    .A2(net5011),
    .Y(_01762_),
    .B1(_08076_));
 sg13g2_nor2_1 _26123_ (.A(net3510),
    .B(net5010),
    .Y(_08077_));
 sg13g2_a21oi_1 _26124_ (.A1(net5630),
    .A2(net5010),
    .Y(_01763_),
    .B1(_08077_));
 sg13g2_nor2_1 _26125_ (.A(_03134_),
    .B(net5237),
    .Y(_08078_));
 sg13g2_nor2_1 _26126_ (.A(net3079),
    .B(net5009),
    .Y(_08079_));
 sg13g2_a21oi_1 _26127_ (.A1(net5769),
    .A2(net5009),
    .Y(_01764_),
    .B1(_08079_));
 sg13g2_nor2_1 _26128_ (.A(net3099),
    .B(net5008),
    .Y(_08080_));
 sg13g2_a21oi_1 _26129_ (.A1(net5789),
    .A2(net5008),
    .Y(_01765_),
    .B1(_08080_));
 sg13g2_nor2_1 _26130_ (.A(net3713),
    .B(net5009),
    .Y(_08081_));
 sg13g2_a21oi_1 _26131_ (.A1(net5719),
    .A2(net5008),
    .Y(_01766_),
    .B1(_08081_));
 sg13g2_nor2_1 _26132_ (.A(net3637),
    .B(net5009),
    .Y(_08082_));
 sg13g2_a21oi_1 _26133_ (.A1(net5696),
    .A2(net5009),
    .Y(_01767_),
    .B1(_08082_));
 sg13g2_nor2_1 _26134_ (.A(net3370),
    .B(net5008),
    .Y(_08083_));
 sg13g2_a21oi_1 _26135_ (.A1(net5674),
    .A2(net5008),
    .Y(_01768_),
    .B1(_08083_));
 sg13g2_nor2_1 _26136_ (.A(net3259),
    .B(net5009),
    .Y(_08084_));
 sg13g2_a21oi_1 _26137_ (.A1(net5594),
    .A2(net5008),
    .Y(_01769_),
    .B1(_08084_));
 sg13g2_nor2_1 _26138_ (.A(net3980),
    .B(net5008),
    .Y(_08085_));
 sg13g2_a21oi_1 _26139_ (.A1(net5655),
    .A2(net5008),
    .Y(_01770_),
    .B1(_08085_));
 sg13g2_nor2_1 _26140_ (.A(net3379),
    .B(net5009),
    .Y(_08086_));
 sg13g2_a21oi_1 _26141_ (.A1(net5630),
    .A2(net5009),
    .Y(_01771_),
    .B1(_08086_));
 sg13g2_nor2_1 _26142_ (.A(net6522),
    .B(net5532),
    .Y(_01772_));
 sg13g2_and2_1 _26143_ (.A(net6543),
    .B(net5564),
    .X(_01773_));
 sg13g2_nor2_1 _26144_ (.A(net6522),
    .B(net5560),
    .Y(_01774_));
 sg13g2_nor2_1 _26145_ (.A(net6524),
    .B(net5548),
    .Y(_01775_));
 sg13g2_nor2_1 _26146_ (.A(net6524),
    .B(net5279),
    .Y(_01776_));
 sg13g2_nor2_1 _26147_ (.A(net6524),
    .B(net5569),
    .Y(_01777_));
 sg13g2_nor2_1 _26148_ (.A(net6524),
    .B(net5543),
    .Y(_01778_));
 sg13g2_and2_1 _26149_ (.A(net6543),
    .B(net5514),
    .X(_01779_));
 sg13g2_nor2_1 _26150_ (.A(net6522),
    .B(_09272_),
    .Y(_01780_));
 sg13g2_nor2_1 _26151_ (.A(net6522),
    .B(_09278_),
    .Y(_01781_));
 sg13g2_nor2_1 _26152_ (.A(net6522),
    .B(_09283_),
    .Y(_01782_));
 sg13g2_and2_1 _26153_ (.A(net6543),
    .B(net5541),
    .X(_01783_));
 sg13g2_nor2_1 _26154_ (.A(net6522),
    .B(net5536),
    .Y(_01784_));
 sg13g2_nor2_1 _26155_ (.A(_03134_),
    .B(net5249),
    .Y(_08087_));
 sg13g2_nor2_1 _26156_ (.A(net3009),
    .B(net5007),
    .Y(_08088_));
 sg13g2_a21oi_1 _26157_ (.A1(net5769),
    .A2(net5007),
    .Y(_01785_),
    .B1(_08088_));
 sg13g2_nor2_1 _26158_ (.A(net4449),
    .B(net5006),
    .Y(_08089_));
 sg13g2_a21oi_1 _26159_ (.A1(net5789),
    .A2(net5006),
    .Y(_01786_),
    .B1(_08089_));
 sg13g2_nor2_1 _26160_ (.A(net3069),
    .B(net5007),
    .Y(_08090_));
 sg13g2_a21oi_1 _26161_ (.A1(net5719),
    .A2(net5007),
    .Y(_01787_),
    .B1(_08090_));
 sg13g2_nor2_1 _26162_ (.A(net3401),
    .B(net5007),
    .Y(_08091_));
 sg13g2_a21oi_1 _26163_ (.A1(net5696),
    .A2(net5007),
    .Y(_01788_),
    .B1(_08091_));
 sg13g2_nor2_1 _26164_ (.A(net3277),
    .B(net5006),
    .Y(_08092_));
 sg13g2_a21oi_1 _26165_ (.A1(net5674),
    .A2(net5006),
    .Y(_01789_),
    .B1(_08092_));
 sg13g2_nor2_1 _26166_ (.A(net3218),
    .B(net5006),
    .Y(_08093_));
 sg13g2_a21oi_1 _26167_ (.A1(net5594),
    .A2(net5006),
    .Y(_01790_),
    .B1(_08093_));
 sg13g2_nor2_1 _26168_ (.A(net4060),
    .B(net5006),
    .Y(_08094_));
 sg13g2_a21oi_1 _26169_ (.A1(net5655),
    .A2(net5006),
    .Y(_01791_),
    .B1(_08094_));
 sg13g2_nor2_1 _26170_ (.A(net3201),
    .B(net5007),
    .Y(_08095_));
 sg13g2_a21oi_1 _26171_ (.A1(net5630),
    .A2(net5007),
    .Y(_01792_),
    .B1(_08095_));
 sg13g2_nand3_1 _26172_ (.B(_09329_),
    .C(net5252),
    .A(net5556),
    .Y(_08096_));
 sg13g2_mux2_1 _26173_ (.A0(net5740),
    .A1(net4852),
    .S(_08096_),
    .X(_01793_));
 sg13g2_mux2_1 _26174_ (.A0(net5745),
    .A1(net4663),
    .S(_08096_),
    .X(_01794_));
 sg13g2_mux2_1 _26175_ (.A0(net5621),
    .A1(net4619),
    .S(_08096_),
    .X(_01795_));
 sg13g2_mux2_1 _26176_ (.A0(net5615),
    .A1(net7033),
    .S(_08096_),
    .X(_01796_));
 sg13g2_mux2_1 _26177_ (.A0(net5607),
    .A1(net4620),
    .S(_08096_),
    .X(_01797_));
 sg13g2_mux2_1 _26178_ (.A0(net5582),
    .A1(net6666),
    .S(_08096_),
    .X(_01798_));
 sg13g2_mux2_1 _26179_ (.A0(net5575),
    .A1(net6697),
    .S(_08096_),
    .X(_01799_));
 sg13g2_mux2_1 _26180_ (.A0(net5641),
    .A1(net6633),
    .S(_08096_),
    .X(_01800_));
 sg13g2_nor2_1 _26181_ (.A(_09331_),
    .B(net5257),
    .Y(_08097_));
 sg13g2_nor2_1 _26182_ (.A(net4366),
    .B(net5005),
    .Y(_08098_));
 sg13g2_a21oi_1 _26183_ (.A1(net5762),
    .A2(net5005),
    .Y(_01801_),
    .B1(_08098_));
 sg13g2_nor2_1 _26184_ (.A(net3654),
    .B(net5005),
    .Y(_08099_));
 sg13g2_a21oi_1 _26185_ (.A1(net5782),
    .A2(net5005),
    .Y(_01802_),
    .B1(_08099_));
 sg13g2_nor2_1 _26186_ (.A(net3996),
    .B(net5004),
    .Y(_08100_));
 sg13g2_a21oi_1 _26187_ (.A1(net5712),
    .A2(net5004),
    .Y(_01803_),
    .B1(_08100_));
 sg13g2_nor2_1 _26188_ (.A(net3564),
    .B(net5005),
    .Y(_08101_));
 sg13g2_a21oi_1 _26189_ (.A1(net5690),
    .A2(net5005),
    .Y(_01804_),
    .B1(_08101_));
 sg13g2_nor2_1 _26190_ (.A(net3188),
    .B(net5004),
    .Y(_08102_));
 sg13g2_a21oi_1 _26191_ (.A1(net5669),
    .A2(net5004),
    .Y(_01805_),
    .B1(_08102_));
 sg13g2_nor2_1 _26192_ (.A(net4285),
    .B(net5005),
    .Y(_08103_));
 sg13g2_a21oi_1 _26193_ (.A1(net5591),
    .A2(net5005),
    .Y(_01806_),
    .B1(_08103_));
 sg13g2_nor2_1 _26194_ (.A(net3387),
    .B(net5004),
    .Y(_08104_));
 sg13g2_a21oi_1 _26195_ (.A1(net5650),
    .A2(net5004),
    .Y(_01807_),
    .B1(_08104_));
 sg13g2_nor2_1 _26196_ (.A(net4027),
    .B(net5004),
    .Y(_08105_));
 sg13g2_a21oi_1 _26197_ (.A1(net5629),
    .A2(net5004),
    .Y(_01808_),
    .B1(_08105_));
 sg13g2_and2_1 _26198_ (.A(\flash_rom.spi_select ),
    .B(_03203_),
    .X(_08106_));
 sg13g2_or2_1 _26199_ (.X(_08107_),
    .B(_08106_),
    .A(_07827_));
 sg13g2_nor2_2 _26200_ (.A(\flash_rom.spi_select ),
    .B(_07827_),
    .Y(_08108_));
 sg13g2_inv_1 _26201_ (.Y(_08109_),
    .A(_08108_));
 sg13g2_nor2_1 _26202_ (.A(_00112_),
    .B(\flash_rom.spi_select ),
    .Y(_08110_));
 sg13g2_xnor2_1 _26203_ (.Y(_08111_),
    .A(net6245),
    .B(\flash_rom.fsm_state[1] ));
 sg13g2_nand4_1 _26204_ (.B(_07829_),
    .C(_08110_),
    .A(_11057_),
    .Y(_08112_),
    .D(_08111_));
 sg13g2_o21ai_1 _26205_ (.B1(_08112_),
    .Y(_08113_),
    .A1(\flash_rom.spi_clk_out ),
    .A2(_08109_));
 sg13g2_nor2_1 _26206_ (.A(_08107_),
    .B(_08113_),
    .Y(_08114_));
 sg13g2_and3_1 _26207_ (.X(_08115_),
    .A(\flash_rom.spi_clk_out ),
    .B(_08108_),
    .C(_08112_));
 sg13g2_o21ai_1 _26208_ (.B1(_07826_),
    .Y(_08116_),
    .A1(net7393),
    .A2(_08114_));
 sg13g2_a21oi_1 _26209_ (.A1(net7393),
    .A2(_08115_),
    .Y(_01809_),
    .B1(_08116_));
 sg13g2_nand2_1 _26210_ (.Y(_08117_),
    .A(\flash_rom.fsm_state[1] ),
    .B(net7562));
 sg13g2_nor2_1 _26211_ (.A(net6245),
    .B(_08117_),
    .Y(_08118_));
 sg13g2_o21ai_1 _26212_ (.B1(_07829_),
    .Y(_08119_),
    .A1(net6245),
    .A2(_08117_));
 sg13g2_xnor2_1 _26213_ (.Y(_08120_),
    .A(net7475),
    .B(net7393));
 sg13g2_nand2_1 _26214_ (.Y(_08121_),
    .A(_08119_),
    .B(_08120_));
 sg13g2_o21ai_1 _26215_ (.B1(_07826_),
    .Y(_08122_),
    .A1(net7475),
    .A2(_08114_));
 sg13g2_a21oi_1 _26216_ (.A1(_08115_),
    .A2(_08121_),
    .Y(_01810_),
    .B1(_08122_));
 sg13g2_nand3_1 _26217_ (.B(_11056_),
    .C(_07829_),
    .A(net7303),
    .Y(_08123_));
 sg13g2_nand3_1 _26218_ (.B(_08115_),
    .C(_08123_),
    .A(_11058_),
    .Y(_08124_));
 sg13g2_o21ai_1 _26219_ (.B1(_08124_),
    .Y(_08125_),
    .A1(net7444),
    .A2(_08114_));
 sg13g2_nor2_1 _26220_ (.A(_07825_),
    .B(_08125_),
    .Y(_01811_));
 sg13g2_nor3_1 _26221_ (.A(\flash_rom.stall_read ),
    .B(_07828_),
    .C(_07830_),
    .Y(_08126_));
 sg13g2_a221oi_1 _26222_ (.B2(_08108_),
    .C1(_08126_),
    .B1(_07830_),
    .A1(\flash_rom.stall_read ),
    .Y(_08127_),
    .A2(_07827_));
 sg13g2_nand2b_2 _26223_ (.Y(_08128_),
    .B(_08127_),
    .A_N(_08106_));
 sg13g2_inv_1 _26224_ (.Y(_08129_),
    .A(_08128_));
 sg13g2_a21oi_1 _26225_ (.A1(net4155),
    .A2(_07828_),
    .Y(_08130_),
    .B1(_08128_));
 sg13g2_a221oi_1 _26226_ (.B2(_08108_),
    .C1(_07825_),
    .B1(_08130_),
    .A1(_08473_),
    .Y(_01812_),
    .A2(_08128_));
 sg13g2_nor3_1 _26227_ (.A(_11055_),
    .B(_11056_),
    .C(_08128_),
    .Y(_08131_));
 sg13g2_nor2_1 _26228_ (.A(net7509),
    .B(_08129_),
    .Y(_08132_));
 sg13g2_nor3_1 _26229_ (.A(_07825_),
    .B(_08131_),
    .C(_08132_),
    .Y(_01813_));
 sg13g2_o21ai_1 _26230_ (.B1(net6245),
    .Y(_08133_),
    .A1(_08117_),
    .A2(_08128_));
 sg13g2_o21ai_1 _26231_ (.B1(_08129_),
    .Y(_08134_),
    .A1(_07827_),
    .A2(_08118_));
 sg13g2_a21oi_1 _26232_ (.A1(_08133_),
    .A2(_08134_),
    .Y(_01814_),
    .B1(_07825_));
 sg13g2_nor2_2 _26233_ (.A(_00112_),
    .B(_07828_),
    .Y(_08135_));
 sg13g2_mux2_1 _26234_ (.A0(net4793),
    .A1(net9),
    .S(net5941),
    .X(_01815_));
 sg13g2_mux2_1 _26235_ (.A0(net7402),
    .A1(net10),
    .S(_08135_),
    .X(_01816_));
 sg13g2_mux2_1 _26236_ (.A0(net4846),
    .A1(net11),
    .S(net5941),
    .X(_01817_));
 sg13g2_mux2_1 _26237_ (.A0(net4903),
    .A1(net12),
    .S(net5941),
    .X(_01818_));
 sg13g2_mux2_1 _26238_ (.A0(net3488),
    .A1(\external_rom_data[0] ),
    .S(net5941),
    .X(_01819_));
 sg13g2_mux2_1 _26239_ (.A0(net3356),
    .A1(\external_rom_data[1] ),
    .S(net5941),
    .X(_01820_));
 sg13g2_mux2_1 _26240_ (.A0(net4165),
    .A1(\external_rom_data[2] ),
    .S(net5941),
    .X(_01821_));
 sg13g2_mux2_1 _26241_ (.A0(net4380),
    .A1(\external_rom_data[3] ),
    .S(net5941),
    .X(_01822_));
 sg13g2_a22oi_1 _26242_ (.Y(_08136_),
    .B1(_08108_),
    .B2(net7428),
    .A2(_08107_),
    .A1(\flash_rom.spi_clk_out ));
 sg13g2_nand2_1 _26243_ (.Y(_01823_),
    .A(_07826_),
    .B(net7429));
 sg13g2_mux2_1 _26244_ (.A0(_00132_),
    .A1(\flash_rom.fsm_state[2] ),
    .S(\flash_rom.fsm_state[1] ),
    .X(_08137_));
 sg13g2_nand3_1 _26245_ (.B(_09038_),
    .C(_08137_),
    .A(\flash_rom.spi_clk_out ),
    .Y(_08138_));
 sg13g2_nor2_1 _26246_ (.A(net5976),
    .B(net5941),
    .Y(_08139_));
 sg13g2_nand2_1 _26247_ (.Y(_08140_),
    .A(_08138_),
    .B(_08139_));
 sg13g2_a221oi_1 _26248_ (.B2(_07829_),
    .C1(_08107_),
    .B1(_08140_),
    .A1(_09038_),
    .Y(_08141_),
    .A2(_07830_));
 sg13g2_o21ai_1 _26249_ (.B1(_08141_),
    .Y(_08142_),
    .A1(net6245),
    .A2(\flash_rom.fsm_state[1] ));
 sg13g2_o21ai_1 _26250_ (.B1(_07826_),
    .Y(_08143_),
    .A1(net7297),
    .A2(_08141_));
 sg13g2_nor2b_1 _26251_ (.A(_08143_),
    .B_N(_08142_),
    .Y(_01824_));
 sg13g2_o21ai_1 _26252_ (.B1(_07826_),
    .Y(_08144_),
    .A1(uio_oe[5]),
    .A2(_08141_));
 sg13g2_a21oi_1 _26253_ (.A1(net7304),
    .A2(_08141_),
    .Y(_01825_),
    .B1(_08144_));
 sg13g2_o21ai_1 _26254_ (.B1(_09173_),
    .Y(_08145_),
    .A1(_09202_),
    .A2(_09203_));
 sg13g2_nand3_1 _26255_ (.B(net6563),
    .C(_08145_),
    .A(net7368),
    .Y(_08146_));
 sg13g2_o21ai_1 _26256_ (.B1(_08146_),
    .Y(_01826_),
    .A1(net5080),
    .A2(_09201_));
 sg13g2_a22oi_1 _26257_ (.Y(_08147_),
    .B1(_08145_),
    .B2(net7335),
    .A2(_09203_),
    .A1(_09173_));
 sg13g2_nor2_1 _26258_ (.A(net6533),
    .B(_08147_),
    .Y(_01827_));
 sg13g2_nand3_1 _26259_ (.B(net6561),
    .C(_08145_),
    .A(net7361),
    .Y(_08148_));
 sg13g2_o21ai_1 _26260_ (.B1(_08148_),
    .Y(_01828_),
    .A1(net5080),
    .A2(_05513_));
 sg13g2_nor2_1 _26261_ (.A(net5259),
    .B(_07321_),
    .Y(_08149_));
 sg13g2_nor2_1 _26262_ (.A(net4420),
    .B(net5002),
    .Y(_08150_));
 sg13g2_a21oi_1 _26263_ (.A1(net5760),
    .A2(net5002),
    .Y(_01829_),
    .B1(_08150_));
 sg13g2_nor2_1 _26264_ (.A(net4032),
    .B(net5002),
    .Y(_08151_));
 sg13g2_a21oi_1 _26265_ (.A1(net5781),
    .A2(net5002),
    .Y(_01830_),
    .B1(_08151_));
 sg13g2_nor2_1 _26266_ (.A(net3380),
    .B(net5002),
    .Y(_08152_));
 sg13g2_a21oi_1 _26267_ (.A1(net5711),
    .A2(net5002),
    .Y(_01831_),
    .B1(_08152_));
 sg13g2_nor2_1 _26268_ (.A(net3321),
    .B(net5003),
    .Y(_08153_));
 sg13g2_a21oi_1 _26269_ (.A1(net5689),
    .A2(net5003),
    .Y(_01832_),
    .B1(_08153_));
 sg13g2_nor2_1 _26270_ (.A(net4217),
    .B(net5002),
    .Y(_08154_));
 sg13g2_a21oi_1 _26271_ (.A1(net5666),
    .A2(net5002),
    .Y(_01833_),
    .B1(_08154_));
 sg13g2_nor2_1 _26272_ (.A(net3416),
    .B(net5003),
    .Y(_08155_));
 sg13g2_a21oi_1 _26273_ (.A1(net5588),
    .A2(net5003),
    .Y(_01834_),
    .B1(_08155_));
 sg13g2_nor2_1 _26274_ (.A(net3482),
    .B(net5003),
    .Y(_08156_));
 sg13g2_a21oi_1 _26275_ (.A1(net5648),
    .A2(net5003),
    .Y(_01835_),
    .B1(_08156_));
 sg13g2_nor2_1 _26276_ (.A(net4771),
    .B(net5003),
    .Y(_08157_));
 sg13g2_a21oi_1 _26277_ (.A1(net5625),
    .A2(net5003),
    .Y(_01836_),
    .B1(_08157_));
 sg13g2_nand2_2 _26278_ (.Y(_08158_),
    .A(net5250),
    .B(_07320_));
 sg13g2_mux2_1 _26279_ (.A0(net5740),
    .A1(net4761),
    .S(_08158_),
    .X(_01837_));
 sg13g2_mux2_1 _26280_ (.A0(net5745),
    .A1(net4455),
    .S(_08158_),
    .X(_01838_));
 sg13g2_mux2_1 _26281_ (.A0(net5616),
    .A1(net4458),
    .S(_08158_),
    .X(_01839_));
 sg13g2_mux2_1 _26282_ (.A0(net5611),
    .A1(net7013),
    .S(_08158_),
    .X(_01840_));
 sg13g2_mux2_1 _26283_ (.A0(net5607),
    .A1(net6640),
    .S(_08158_),
    .X(_01841_));
 sg13g2_mux2_1 _26284_ (.A0(net5580),
    .A1(net4469),
    .S(_08158_),
    .X(_01842_));
 sg13g2_mux2_1 _26285_ (.A0(net5575),
    .A1(net4682),
    .S(_08158_),
    .X(_01843_));
 sg13g2_mux2_1 _26286_ (.A0(net5641),
    .A1(net6779),
    .S(_08158_),
    .X(_01844_));
 sg13g2_nor2_1 _26287_ (.A(net5237),
    .B(_07321_),
    .Y(_08159_));
 sg13g2_nor2_1 _26288_ (.A(net3001),
    .B(net5000),
    .Y(_08160_));
 sg13g2_a21oi_1 _26289_ (.A1(net5760),
    .A2(net5000),
    .Y(_01845_),
    .B1(_08160_));
 sg13g2_nor2_1 _26290_ (.A(net3724),
    .B(net5000),
    .Y(_08161_));
 sg13g2_a21oi_1 _26291_ (.A1(net5781),
    .A2(net5000),
    .Y(_01846_),
    .B1(_08161_));
 sg13g2_nor2_1 _26292_ (.A(net3058),
    .B(net5000),
    .Y(_08162_));
 sg13g2_a21oi_1 _26293_ (.A1(net5709),
    .A2(net5000),
    .Y(_01847_),
    .B1(_08162_));
 sg13g2_nor2_1 _26294_ (.A(net3124),
    .B(net5001),
    .Y(_08163_));
 sg13g2_a21oi_1 _26295_ (.A1(net5689),
    .A2(net5001),
    .Y(_01848_),
    .B1(_08163_));
 sg13g2_nor2_1 _26296_ (.A(net4440),
    .B(net5000),
    .Y(_08164_));
 sg13g2_a21oi_1 _26297_ (.A1(net5666),
    .A2(net5000),
    .Y(_01849_),
    .B1(_08164_));
 sg13g2_nor2_1 _26298_ (.A(net3034),
    .B(net5001),
    .Y(_08165_));
 sg13g2_a21oi_1 _26299_ (.A1(net5587),
    .A2(net5001),
    .Y(_01850_),
    .B1(_08165_));
 sg13g2_nor2_1 _26300_ (.A(net3522),
    .B(net5001),
    .Y(_08166_));
 sg13g2_a21oi_1 _26301_ (.A1(net5648),
    .A2(net5001),
    .Y(_01851_),
    .B1(_08166_));
 sg13g2_nor2_1 _26302_ (.A(net3132),
    .B(net5001),
    .Y(_08167_));
 sg13g2_a21oi_1 _26303_ (.A1(net5625),
    .A2(net5001),
    .Y(_01852_),
    .B1(_08167_));
 sg13g2_nor2_1 _26304_ (.A(net5249),
    .B(_07321_),
    .Y(_08168_));
 sg13g2_nor2_1 _26305_ (.A(net3193),
    .B(net4998),
    .Y(_08169_));
 sg13g2_a21oi_1 _26306_ (.A1(net5760),
    .A2(net4998),
    .Y(_01853_),
    .B1(_08169_));
 sg13g2_nor2_1 _26307_ (.A(net3318),
    .B(net4998),
    .Y(_08170_));
 sg13g2_a21oi_1 _26308_ (.A1(net5781),
    .A2(net4998),
    .Y(_01854_),
    .B1(_08170_));
 sg13g2_nor2_1 _26309_ (.A(net3323),
    .B(net4998),
    .Y(_08171_));
 sg13g2_a21oi_1 _26310_ (.A1(net5709),
    .A2(net4998),
    .Y(_01855_),
    .B1(_08171_));
 sg13g2_nor2_1 _26311_ (.A(net3046),
    .B(net4999),
    .Y(_08172_));
 sg13g2_a21oi_1 _26312_ (.A1(net5689),
    .A2(net4999),
    .Y(_01856_),
    .B1(_08172_));
 sg13g2_nor2_1 _26313_ (.A(net3377),
    .B(net4998),
    .Y(_08173_));
 sg13g2_a21oi_1 _26314_ (.A1(net5666),
    .A2(net4998),
    .Y(_01857_),
    .B1(_08173_));
 sg13g2_nor2_1 _26315_ (.A(net4553),
    .B(net4999),
    .Y(_08174_));
 sg13g2_a21oi_1 _26316_ (.A1(net5587),
    .A2(net4999),
    .Y(_01858_),
    .B1(_08174_));
 sg13g2_nor2_1 _26317_ (.A(net4048),
    .B(net4999),
    .Y(_08175_));
 sg13g2_a21oi_1 _26318_ (.A1(net5648),
    .A2(net4999),
    .Y(_01859_),
    .B1(_08175_));
 sg13g2_nor2_1 _26319_ (.A(net3023),
    .B(net4999),
    .Y(_08176_));
 sg13g2_a21oi_1 _26320_ (.A1(net5625),
    .A2(net4999),
    .Y(_01860_),
    .B1(_08176_));
 sg13g2_and2_2 _26321_ (.A(_09413_),
    .B(net5250),
    .X(_08177_));
 sg13g2_nor2_1 _26322_ (.A(net3647),
    .B(net4997),
    .Y(_08178_));
 sg13g2_a21oi_1 _26323_ (.A1(net5762),
    .A2(net4997),
    .Y(_01861_),
    .B1(_08178_));
 sg13g2_nor2_1 _26324_ (.A(net6908),
    .B(net4997),
    .Y(_08179_));
 sg13g2_a21oi_1 _26325_ (.A1(net5782),
    .A2(net4997),
    .Y(_01862_),
    .B1(_08179_));
 sg13g2_nor2_1 _26326_ (.A(net3675),
    .B(net4996),
    .Y(_08180_));
 sg13g2_a21oi_1 _26327_ (.A1(net5712),
    .A2(net4996),
    .Y(_01863_),
    .B1(_08180_));
 sg13g2_nor2_1 _26328_ (.A(net4302),
    .B(net4997),
    .Y(_08181_));
 sg13g2_a21oi_1 _26329_ (.A1(net5690),
    .A2(net4997),
    .Y(_01864_),
    .B1(_08181_));
 sg13g2_nor2_1 _26330_ (.A(net3174),
    .B(net4996),
    .Y(_08182_));
 sg13g2_a21oi_1 _26331_ (.A1(net5668),
    .A2(net4996),
    .Y(_01865_),
    .B1(_08182_));
 sg13g2_nor2_1 _26332_ (.A(net3807),
    .B(net4997),
    .Y(_08183_));
 sg13g2_a21oi_1 _26333_ (.A1(net5591),
    .A2(net4997),
    .Y(_01866_),
    .B1(_08183_));
 sg13g2_nor2_1 _26334_ (.A(net3425),
    .B(net4996),
    .Y(_08184_));
 sg13g2_a21oi_1 _26335_ (.A1(net5650),
    .A2(net4996),
    .Y(_01867_),
    .B1(_08184_));
 sg13g2_nor2_1 _26336_ (.A(net3816),
    .B(net4996),
    .Y(_08185_));
 sg13g2_a21oi_1 _26337_ (.A1(net5629),
    .A2(net4996),
    .Y(_01868_),
    .B1(_08185_));
 sg13g2_nor2_1 _26338_ (.A(_09422_),
    .B(net5257),
    .Y(_08186_));
 sg13g2_nor2_1 _26339_ (.A(net4196),
    .B(net4995),
    .Y(_08187_));
 sg13g2_a21oi_1 _26340_ (.A1(net5759),
    .A2(net4994),
    .Y(_01869_),
    .B1(_08187_));
 sg13g2_nor2_1 _26341_ (.A(net3552),
    .B(net4994),
    .Y(_08188_));
 sg13g2_a21oi_1 _26342_ (.A1(net5780),
    .A2(net4994),
    .Y(_01870_),
    .B1(_08188_));
 sg13g2_nor2_1 _26343_ (.A(net4255),
    .B(_08186_),
    .Y(_08189_));
 sg13g2_a21oi_1 _26344_ (.A1(net5709),
    .A2(net4995),
    .Y(_01871_),
    .B1(_08189_));
 sg13g2_nor2_1 _26345_ (.A(net4742),
    .B(net4995),
    .Y(_08190_));
 sg13g2_a21oi_1 _26346_ (.A1(net5686),
    .A2(net4995),
    .Y(_01872_),
    .B1(_08190_));
 sg13g2_nor2_1 _26347_ (.A(net3223),
    .B(net4994),
    .Y(_08191_));
 sg13g2_a21oi_1 _26348_ (.A1(net5666),
    .A2(net4994),
    .Y(_01873_),
    .B1(_08191_));
 sg13g2_nor2_1 _26349_ (.A(net3554),
    .B(net4995),
    .Y(_08192_));
 sg13g2_a21oi_1 _26350_ (.A1(net5585),
    .A2(net4995),
    .Y(_01874_),
    .B1(_08192_));
 sg13g2_nor2_1 _26351_ (.A(net3372),
    .B(net4994),
    .Y(_08193_));
 sg13g2_a21oi_1 _26352_ (.A1(net5649),
    .A2(net4994),
    .Y(_01875_),
    .B1(_08193_));
 sg13g2_nor2_1 _26353_ (.A(net4049),
    .B(net4995),
    .Y(_08194_));
 sg13g2_a21oi_1 _26354_ (.A1(net5622),
    .A2(net4994),
    .Y(_01876_),
    .B1(_08194_));
 sg13g2_nor2_1 _26355_ (.A(net5939),
    .B(net5814),
    .Y(_08195_));
 sg13g2_a221oi_1 _26356_ (.B2(net6249),
    .C1(net5750),
    .B1(net5948),
    .A1(\atari2600.cpu.DIMUX[5] ),
    .Y(_08196_),
    .A2(net5927));
 sg13g2_a21oi_1 _26357_ (.A1(_08658_),
    .A2(_09082_),
    .Y(_08197_),
    .B1(_08196_));
 sg13g2_mux2_1 _26358_ (.A0(net7125),
    .A1(_08197_),
    .S(_08195_),
    .X(_01877_));
 sg13g2_o21ai_1 _26359_ (.B1(net4386),
    .Y(_08198_),
    .A1(net5939),
    .A2(net5814));
 sg13g2_a221oi_1 _26360_ (.B2(net6248),
    .C1(net5750),
    .B1(net5948),
    .A1(net5825),
    .Y(_08199_),
    .A2(net5927));
 sg13g2_nor2_1 _26361_ (.A(\atari2600.cpu.PC[14] ),
    .B(_09083_),
    .Y(_08200_));
 sg13g2_nand2b_1 _26362_ (.Y(_08201_),
    .B(_08195_),
    .A_N(_08199_));
 sg13g2_o21ai_1 _26363_ (.B1(_08198_),
    .Y(_01878_),
    .A1(_08200_),
    .A2(_08201_));
 sg13g2_o21ai_1 _26364_ (.B1(net4452),
    .Y(_08202_),
    .A1(net5939),
    .A2(net5814));
 sg13g2_a221oi_1 _26365_ (.B2(\atari2600.cpu.ADD[7] ),
    .C1(net5750),
    .B1(net5948),
    .A1(\atari2600.cpu.DIMUX[7] ),
    .Y(_08203_),
    .A2(net5927));
 sg13g2_o21ai_1 _26366_ (.B1(_08195_),
    .Y(_08204_),
    .A1(\atari2600.cpu.PC[15] ),
    .A2(_09083_));
 sg13g2_o21ai_1 _26367_ (.B1(_08202_),
    .Y(_01879_),
    .A1(_08203_),
    .A2(_08204_));
 sg13g2_o21ai_1 _26368_ (.B1(net6582),
    .Y(_08205_),
    .A1(net6208),
    .A2(_03191_));
 sg13g2_a21oi_1 _26369_ (.A1(net6208),
    .A2(_03191_),
    .Y(_01880_),
    .B1(_08205_));
 sg13g2_a21oi_1 _26370_ (.A1(net6209),
    .A2(_03191_),
    .Y(_08206_),
    .B1(net6153));
 sg13g2_nand2_1 _26371_ (.Y(_08207_),
    .A(net6582),
    .B(_03192_));
 sg13g2_nor2_1 _26372_ (.A(_08206_),
    .B(_08207_),
    .Y(_01881_));
 sg13g2_xor2_1 _26373_ (.B(_03192_),
    .A(net6134),
    .X(_08208_));
 sg13g2_nor2_1 _26374_ (.A(_03199_),
    .B(_08208_),
    .Y(_01882_));
 sg13g2_nor2_1 _26375_ (.A(net3016),
    .B(_03192_),
    .Y(_08209_));
 sg13g2_xnor2_1 _26376_ (.Y(_08210_),
    .A(net6133),
    .B(_08209_));
 sg13g2_nor2_1 _26377_ (.A(_03199_),
    .B(net3017),
    .Y(_01883_));
 sg13g2_nor2_1 _26378_ (.A(net6092),
    .B(_03192_),
    .Y(_08211_));
 sg13g2_xnor2_1 _26379_ (.Y(_08212_),
    .A(net6128),
    .B(_08211_));
 sg13g2_nor2_1 _26380_ (.A(_03199_),
    .B(_08212_),
    .Y(_01884_));
 sg13g2_nor3_1 _26381_ (.A(net3144),
    .B(net6092),
    .C(_03192_),
    .Y(_08213_));
 sg13g2_xnor2_1 _26382_ (.Y(_08214_),
    .A(\hvsync_gen.hpos[7] ),
    .B(_08213_));
 sg13g2_nor2_1 _26383_ (.A(_03199_),
    .B(net3145),
    .Y(_01885_));
 sg13g2_nor2_1 _26384_ (.A(_09224_),
    .B(_03192_),
    .Y(_08215_));
 sg13g2_xnor2_1 _26385_ (.Y(_08216_),
    .A(net6126),
    .B(_08215_));
 sg13g2_nor2_1 _26386_ (.A(_03199_),
    .B(_08216_),
    .Y(_01886_));
 sg13g2_nor3_1 _26387_ (.A(net7254),
    .B(_09224_),
    .C(_03192_),
    .Y(_08217_));
 sg13g2_o21ai_1 _26388_ (.B1(_03198_),
    .Y(_08218_),
    .A1(net6125),
    .A2(_08217_));
 sg13g2_a21oi_1 _26389_ (.A1(net6125),
    .A2(_08217_),
    .Y(_01887_),
    .B1(_08218_));
 sg13g2_nor2_1 _26390_ (.A(_09331_),
    .B(net5237),
    .Y(_08219_));
 sg13g2_nor2_1 _26391_ (.A(net3569),
    .B(net4992),
    .Y(_08220_));
 sg13g2_a21oi_1 _26392_ (.A1(net5761),
    .A2(net4992),
    .Y(_01888_),
    .B1(_08220_));
 sg13g2_nor2_1 _26393_ (.A(net3072),
    .B(net4992),
    .Y(_08221_));
 sg13g2_a21oi_1 _26394_ (.A1(net5781),
    .A2(net4992),
    .Y(_01889_),
    .B1(_08221_));
 sg13g2_nor2_1 _26395_ (.A(net3732),
    .B(net4992),
    .Y(_08222_));
 sg13g2_a21oi_1 _26396_ (.A1(net5710),
    .A2(net4992),
    .Y(_01890_),
    .B1(_08222_));
 sg13g2_nor2_1 _26397_ (.A(net4398),
    .B(net4993),
    .Y(_08223_));
 sg13g2_a21oi_1 _26398_ (.A1(net5686),
    .A2(net4993),
    .Y(_01891_),
    .B1(_08223_));
 sg13g2_nor2_1 _26399_ (.A(net3744),
    .B(_08219_),
    .Y(_08224_));
 sg13g2_a21oi_1 _26400_ (.A1(net5667),
    .A2(net4992),
    .Y(_01892_),
    .B1(_08224_));
 sg13g2_nor2_1 _26401_ (.A(net3018),
    .B(net4993),
    .Y(_08225_));
 sg13g2_a21oi_1 _26402_ (.A1(net5587),
    .A2(net4993),
    .Y(_01893_),
    .B1(_08225_));
 sg13g2_nor2_1 _26403_ (.A(net3102),
    .B(net4993),
    .Y(_08226_));
 sg13g2_a21oi_1 _26404_ (.A1(net5649),
    .A2(net4993),
    .Y(_01894_),
    .B1(_08226_));
 sg13g2_nor2_1 _26405_ (.A(net4187),
    .B(net4993),
    .Y(_08227_));
 sg13g2_a21oi_1 _26406_ (.A1(net5624),
    .A2(net4992),
    .Y(_01895_),
    .B1(_08227_));
 sg13g2_nor2_2 _26407_ (.A(_10069_),
    .B(net6067),
    .Y(_08228_));
 sg13g2_and2_1 _26408_ (.A(_10013_),
    .B(net6072),
    .X(_08229_));
 sg13g2_nand2_2 _26409_ (.Y(_08230_),
    .A(_10013_),
    .B(net6072));
 sg13g2_nand2_2 _26410_ (.Y(_08231_),
    .A(net5968),
    .B(net5966));
 sg13g2_mux2_1 _26411_ (.A0(net6466),
    .A1(net7056),
    .S(_08231_),
    .X(_01896_));
 sg13g2_mux2_1 _26412_ (.A0(net6437),
    .A1(net4863),
    .S(_08231_),
    .X(_01897_));
 sg13g2_mux2_1 _26413_ (.A0(net6405),
    .A1(net7177),
    .S(_08231_),
    .X(_01898_));
 sg13g2_mux2_1 _26414_ (.A0(net6378),
    .A1(net7069),
    .S(_08231_),
    .X(_01899_));
 sg13g2_mux2_1 _26415_ (.A0(net6350),
    .A1(net7101),
    .S(_08231_),
    .X(_01900_));
 sg13g2_mux2_1 _26416_ (.A0(net6319),
    .A1(net7052),
    .S(_08231_),
    .X(_01901_));
 sg13g2_mux2_1 _26417_ (.A0(net6290),
    .A1(net4586),
    .S(_08231_),
    .X(_01902_));
 sg13g2_or2_2 _26418_ (.X(_08232_),
    .B(_10136_),
    .A(_10124_));
 sg13g2_nor2_2 _26419_ (.A(_08230_),
    .B(net5965),
    .Y(_08233_));
 sg13g2_mux2_1 _26420_ (.A0(net3414),
    .A1(net6463),
    .S(_08233_),
    .X(_01903_));
 sg13g2_mux2_1 _26421_ (.A0(net3476),
    .A1(net6435),
    .S(_08233_),
    .X(_01904_));
 sg13g2_mux2_1 _26422_ (.A0(net4470),
    .A1(net6406),
    .S(_08233_),
    .X(_01905_));
 sg13g2_mux2_1 _26423_ (.A0(net3442),
    .A1(net6380),
    .S(_08233_),
    .X(_01906_));
 sg13g2_mux2_1 _26424_ (.A0(net4246),
    .A1(net6349),
    .S(_08233_),
    .X(_01907_));
 sg13g2_mux2_1 _26425_ (.A0(net4257),
    .A1(net6323),
    .S(_08233_),
    .X(_01908_));
 sg13g2_mux2_1 _26426_ (.A0(net4063),
    .A1(net6289),
    .S(_08233_),
    .X(_01909_));
 sg13g2_nor2_2 _26427_ (.A(net6501),
    .B(net6124),
    .Y(_08234_));
 sg13g2_nand2_2 _26428_ (.Y(_08235_),
    .A(_08626_),
    .B(net6503));
 sg13g2_nor2_2 _26429_ (.A(net6067),
    .B(_08235_),
    .Y(_08236_));
 sg13g2_nand2_2 _26430_ (.Y(_08237_),
    .A(_10070_),
    .B(_08234_));
 sg13g2_and2_1 _26431_ (.A(_10012_),
    .B(net6072),
    .X(_08238_));
 sg13g2_nand2_2 _26432_ (.Y(_08239_),
    .A(_10012_),
    .B(net6072));
 sg13g2_nand2_2 _26433_ (.Y(_08240_),
    .A(_08236_),
    .B(net5963));
 sg13g2_mux2_1 _26434_ (.A0(net6463),
    .A1(net4570),
    .S(_08240_),
    .X(_01910_));
 sg13g2_mux2_1 _26435_ (.A0(net6437),
    .A1(net6700),
    .S(_08240_),
    .X(_01911_));
 sg13g2_mux2_1 _26436_ (.A0(net6405),
    .A1(net6857),
    .S(_08240_),
    .X(_01912_));
 sg13g2_mux2_1 _26437_ (.A0(net6377),
    .A1(net6940),
    .S(_08240_),
    .X(_01913_));
 sg13g2_mux2_1 _26438_ (.A0(net6350),
    .A1(net4959),
    .S(_08240_),
    .X(_01914_));
 sg13g2_mux2_1 _26439_ (.A0(net6318),
    .A1(net6854),
    .S(_08240_),
    .X(_01915_));
 sg13g2_mux2_1 _26440_ (.A0(net6288),
    .A1(net7001),
    .S(_08240_),
    .X(_01916_));
 sg13g2_nor2_2 _26441_ (.A(_10069_),
    .B(_10124_),
    .Y(_08241_));
 sg13g2_nor2b_2 _26442_ (.A(_10014_),
    .B_N(_10019_),
    .Y(_08242_));
 sg13g2_nand2b_1 _26443_ (.Y(_08243_),
    .B(net6072),
    .A_N(_10014_));
 sg13g2_nand2_2 _26444_ (.Y(_08244_),
    .A(net5962),
    .B(_08242_));
 sg13g2_mux2_1 _26445_ (.A0(net6457),
    .A1(net4855),
    .S(_08244_),
    .X(_01917_));
 sg13g2_mux2_1 _26446_ (.A0(net6428),
    .A1(net4642),
    .S(_08244_),
    .X(_01918_));
 sg13g2_mux2_1 _26447_ (.A0(net6399),
    .A1(net4895),
    .S(_08244_),
    .X(_01919_));
 sg13g2_mux2_1 _26448_ (.A0(net6370),
    .A1(net4856),
    .S(_08244_),
    .X(_01920_));
 sg13g2_mux2_1 _26449_ (.A0(net6342),
    .A1(net4816),
    .S(_08244_),
    .X(_01921_));
 sg13g2_mux2_1 _26450_ (.A0(net6311),
    .A1(net6933),
    .S(_08244_),
    .X(_01922_));
 sg13g2_mux2_1 _26451_ (.A0(net6280),
    .A1(net6758),
    .S(_08244_),
    .X(_01923_));
 sg13g2_nor2_2 _26452_ (.A(net6067),
    .B(_03130_),
    .Y(_08245_));
 sg13g2_nand2_2 _26453_ (.Y(_08246_),
    .A(_10070_),
    .B(_03129_));
 sg13g2_nor2_2 _26454_ (.A(net6000),
    .B(_08246_),
    .Y(_08247_));
 sg13g2_mux2_1 _26455_ (.A0(net4174),
    .A1(net6458),
    .S(_08247_),
    .X(_01924_));
 sg13g2_mux2_1 _26456_ (.A0(net3981),
    .A1(net6427),
    .S(_08247_),
    .X(_01925_));
 sg13g2_mux2_1 _26457_ (.A0(net4316),
    .A1(net6403),
    .S(_08247_),
    .X(_01926_));
 sg13g2_mux2_1 _26458_ (.A0(net3825),
    .A1(net6375),
    .S(_08247_),
    .X(_01927_));
 sg13g2_mux2_1 _26459_ (.A0(net4079),
    .A1(net6346),
    .S(_08247_),
    .X(_01928_));
 sg13g2_mux2_1 _26460_ (.A0(net4311),
    .A1(net6312),
    .S(_08247_),
    .X(_01929_));
 sg13g2_mux2_1 _26461_ (.A0(net3628),
    .A1(net6280),
    .S(_08247_),
    .X(_01930_));
 sg13g2_nor2_2 _26462_ (.A(net6118),
    .B(net6481),
    .Y(_08248_));
 sg13g2_nand2_2 _26463_ (.Y(_08249_),
    .A(net6489),
    .B(_08633_));
 sg13g2_nor2_1 _26464_ (.A(_10002_),
    .B(_08249_),
    .Y(_08250_));
 sg13g2_nor2_2 _26465_ (.A(_10124_),
    .B(_08235_),
    .Y(_08251_));
 sg13g2_nand2_2 _26466_ (.Y(_08252_),
    .A(_10123_),
    .B(_08234_));
 sg13g2_nand2_2 _26467_ (.Y(_08253_),
    .A(net5960),
    .B(_08251_));
 sg13g2_mux2_1 _26468_ (.A0(net6471),
    .A1(net4623),
    .S(_08253_),
    .X(_01931_));
 sg13g2_mux2_1 _26469_ (.A0(net6439),
    .A1(net4549),
    .S(_08253_),
    .X(_01932_));
 sg13g2_mux2_1 _26470_ (.A0(net6412),
    .A1(net7051),
    .S(_08253_),
    .X(_01933_));
 sg13g2_mux2_1 _26471_ (.A0(net6382),
    .A1(net4581),
    .S(_08253_),
    .X(_01934_));
 sg13g2_mux2_1 _26472_ (.A0(net6352),
    .A1(net6953),
    .S(_08253_),
    .X(_01935_));
 sg13g2_mux2_1 _26473_ (.A0(net6324),
    .A1(net4870),
    .S(_08253_),
    .X(_01936_));
 sg13g2_mux2_1 _26474_ (.A0(net6292),
    .A1(net4665),
    .S(_08253_),
    .X(_01937_));
 sg13g2_nor3_2 _26475_ (.A(_10002_),
    .B(net6030),
    .C(_08249_),
    .Y(_08254_));
 sg13g2_mux2_1 _26476_ (.A0(net4076),
    .A1(net6469),
    .S(_08254_),
    .X(_01938_));
 sg13g2_mux2_1 _26477_ (.A0(net3876),
    .A1(net6441),
    .S(_08254_),
    .X(_01939_));
 sg13g2_mux2_1 _26478_ (.A0(net3739),
    .A1(net6409),
    .S(_08254_),
    .X(_01940_));
 sg13g2_mux2_1 _26479_ (.A0(net3848),
    .A1(net6383),
    .S(_08254_),
    .X(_01941_));
 sg13g2_mux2_1 _26480_ (.A0(net3623),
    .A1(net6353),
    .S(_08254_),
    .X(_01942_));
 sg13g2_mux2_1 _26481_ (.A0(net3577),
    .A1(net6325),
    .S(_08254_),
    .X(_01943_));
 sg13g2_mux2_1 _26482_ (.A0(net4274),
    .A1(net6293),
    .S(_08254_),
    .X(_01944_));
 sg13g2_and2_2 _26483_ (.A(_10013_),
    .B(_08248_),
    .X(_08255_));
 sg13g2_nand2_2 _26484_ (.Y(_08256_),
    .A(_10013_),
    .B(_08248_));
 sg13g2_nor2_2 _26485_ (.A(_03132_),
    .B(net5959),
    .Y(_08257_));
 sg13g2_mux2_1 _26486_ (.A0(net3809),
    .A1(net6475),
    .S(_08257_),
    .X(_01945_));
 sg13g2_mux2_1 _26487_ (.A0(net3712),
    .A1(net6449),
    .S(_08257_),
    .X(_01946_));
 sg13g2_mux2_1 _26488_ (.A0(net4333),
    .A1(net6420),
    .S(_08257_),
    .X(_01947_));
 sg13g2_mux2_1 _26489_ (.A0(net3823),
    .A1(net6390),
    .S(_08257_),
    .X(_01948_));
 sg13g2_mux2_1 _26490_ (.A0(net4087),
    .A1(net6361),
    .S(_08257_),
    .X(_01949_));
 sg13g2_mux2_1 _26491_ (.A0(net3704),
    .A1(net6331),
    .S(_08257_),
    .X(_01950_));
 sg13g2_mux2_1 _26492_ (.A0(net3492),
    .A1(net6303),
    .S(_08257_),
    .X(_01951_));
 sg13g2_and2_2 _26493_ (.A(_10012_),
    .B(_08248_),
    .X(_08258_));
 sg13g2_nand2_2 _26494_ (.Y(_08259_),
    .A(_10012_),
    .B(_08248_));
 sg13g2_nand2_2 _26495_ (.Y(_08260_),
    .A(net5968),
    .B(_08258_));
 sg13g2_mux2_1 _26496_ (.A0(net6477),
    .A1(net4818),
    .S(_08260_),
    .X(_01952_));
 sg13g2_mux2_1 _26497_ (.A0(net6446),
    .A1(net6741),
    .S(_08260_),
    .X(_01953_));
 sg13g2_mux2_1 _26498_ (.A0(net6417),
    .A1(net6849),
    .S(_08260_),
    .X(_01954_));
 sg13g2_mux2_1 _26499_ (.A0(net6388),
    .A1(net4905),
    .S(_08260_),
    .X(_01955_));
 sg13g2_mux2_1 _26500_ (.A0(net6359),
    .A1(net4909),
    .S(_08260_),
    .X(_01956_));
 sg13g2_mux2_1 _26501_ (.A0(net6329),
    .A1(net6776),
    .S(_08260_),
    .X(_01957_));
 sg13g2_mux2_1 _26502_ (.A0(net6299),
    .A1(net6639),
    .S(_08260_),
    .X(_01958_));
 sg13g2_nor2_2 _26503_ (.A(net5965),
    .B(_08259_),
    .Y(_08261_));
 sg13g2_mux2_1 _26504_ (.A0(net3484),
    .A1(net6473),
    .S(_08261_),
    .X(_01959_));
 sg13g2_mux2_1 _26505_ (.A0(net4084),
    .A1(net6447),
    .S(_08261_),
    .X(_01960_));
 sg13g2_mux2_1 _26506_ (.A0(net3603),
    .A1(net6421),
    .S(_08261_),
    .X(_01961_));
 sg13g2_mux2_1 _26507_ (.A0(net3955),
    .A1(net6386),
    .S(_08261_),
    .X(_01962_));
 sg13g2_mux2_1 _26508_ (.A0(net3596),
    .A1(net6362),
    .S(_08261_),
    .X(_01963_));
 sg13g2_mux2_1 _26509_ (.A0(net3954),
    .A1(net6332),
    .S(_08261_),
    .X(_01964_));
 sg13g2_mux2_1 _26510_ (.A0(net3914),
    .A1(net6301),
    .S(_08261_),
    .X(_01965_));
 sg13g2_nor2_2 _26511_ (.A(_10014_),
    .B(_08249_),
    .Y(_08262_));
 sg13g2_nand2b_2 _26512_ (.Y(_08263_),
    .B(_08248_),
    .A_N(_10014_));
 sg13g2_nor2_2 _26513_ (.A(_08237_),
    .B(_08263_),
    .Y(_08264_));
 sg13g2_mux2_1 _26514_ (.A0(net4291),
    .A1(net6472),
    .S(_08264_),
    .X(_01966_));
 sg13g2_mux2_1 _26515_ (.A0(net4505),
    .A1(net6443),
    .S(_08264_),
    .X(_01967_));
 sg13g2_mux2_1 _26516_ (.A0(net4233),
    .A1(net6414),
    .S(_08264_),
    .X(_01968_));
 sg13g2_mux2_1 _26517_ (.A0(net4427),
    .A1(net6385),
    .S(_08264_),
    .X(_01969_));
 sg13g2_mux2_1 _26518_ (.A0(net3970),
    .A1(net6356),
    .S(_08264_),
    .X(_01970_));
 sg13g2_mux2_1 _26519_ (.A0(net4262),
    .A1(net6326),
    .S(_08264_),
    .X(_01971_));
 sg13g2_mux2_1 _26520_ (.A0(net4003),
    .A1(net6296),
    .S(_08264_),
    .X(_01972_));
 sg13g2_and2_1 _26521_ (.A(_10001_),
    .B(_10025_),
    .X(_08265_));
 sg13g2_nand2_2 _26522_ (.Y(_08266_),
    .A(_10001_),
    .B(_10025_));
 sg13g2_nand2_2 _26523_ (.Y(_08267_),
    .A(net5962),
    .B(net5956));
 sg13g2_mux2_1 _26524_ (.A0(net6457),
    .A1(net4606),
    .S(_08267_),
    .X(_01973_));
 sg13g2_mux2_1 _26525_ (.A0(net6427),
    .A1(net6752),
    .S(_08267_),
    .X(_01974_));
 sg13g2_mux2_1 _26526_ (.A0(net6399),
    .A1(net4757),
    .S(_08267_),
    .X(_01975_));
 sg13g2_mux2_1 _26527_ (.A0(net6367),
    .A1(net4790),
    .S(_08267_),
    .X(_01976_));
 sg13g2_mux2_1 _26528_ (.A0(net6338),
    .A1(net7186),
    .S(_08267_),
    .X(_01977_));
 sg13g2_mux2_1 _26529_ (.A0(net6314),
    .A1(net4692),
    .S(_08267_),
    .X(_01978_));
 sg13g2_mux2_1 _26530_ (.A0(net6282),
    .A1(net4756),
    .S(_08267_),
    .X(_01979_));
 sg13g2_nand2_2 _26531_ (.Y(_08268_),
    .A(_08245_),
    .B(net5955));
 sg13g2_mux2_1 _26532_ (.A0(net6453),
    .A1(net6726),
    .S(_08268_),
    .X(_01980_));
 sg13g2_mux2_1 _26533_ (.A0(net6424),
    .A1(net4700),
    .S(_08268_),
    .X(_01981_));
 sg13g2_mux2_1 _26534_ (.A0(net6394),
    .A1(net4786),
    .S(_08268_),
    .X(_01982_));
 sg13g2_mux2_1 _26535_ (.A0(net6367),
    .A1(net4918),
    .S(_08268_),
    .X(_01983_));
 sg13g2_mux2_1 _26536_ (.A0(net6338),
    .A1(net6906),
    .S(_08268_),
    .X(_01984_));
 sg13g2_mux2_1 _26537_ (.A0(net6308),
    .A1(net4717),
    .S(_08268_),
    .X(_01985_));
 sg13g2_mux2_1 _26538_ (.A0(net6283),
    .A1(net6904),
    .S(_08268_),
    .X(_01986_));
 sg13g2_and2_2 _26539_ (.A(_10013_),
    .B(_10025_),
    .X(_08269_));
 sg13g2_nand2_2 _26540_ (.Y(_08270_),
    .A(_10013_),
    .B(_10025_));
 sg13g2_nor2_2 _26541_ (.A(_08252_),
    .B(_08270_),
    .Y(_08271_));
 sg13g2_mux2_1 _26542_ (.A0(net4402),
    .A1(net6460),
    .S(_08271_),
    .X(_01987_));
 sg13g2_mux2_1 _26543_ (.A0(net4297),
    .A1(net6432),
    .S(_08271_),
    .X(_01988_));
 sg13g2_mux2_1 _26544_ (.A0(net3983),
    .A1(net6404),
    .S(_08271_),
    .X(_01989_));
 sg13g2_mux2_1 _26545_ (.A0(net3993),
    .A1(net6374),
    .S(_08271_),
    .X(_01990_));
 sg13g2_mux2_1 _26546_ (.A0(net3725),
    .A1(net6345),
    .S(_08271_),
    .X(_01991_));
 sg13g2_mux2_1 _26547_ (.A0(net4372),
    .A1(net6315),
    .S(_08271_),
    .X(_01992_));
 sg13g2_mux2_1 _26548_ (.A0(net4361),
    .A1(net6285),
    .S(_08271_),
    .X(_01993_));
 sg13g2_nor2_2 _26549_ (.A(net6029),
    .B(net5954),
    .Y(_08272_));
 sg13g2_mux2_1 _26550_ (.A0(net4430),
    .A1(net6459),
    .S(_08272_),
    .X(_01994_));
 sg13g2_mux2_1 _26551_ (.A0(net4261),
    .A1(net6431),
    .S(_08272_),
    .X(_01995_));
 sg13g2_mux2_1 _26552_ (.A0(net3991),
    .A1(net6401),
    .S(_08272_),
    .X(_01996_));
 sg13g2_mux2_1 _26553_ (.A0(net3860),
    .A1(net6374),
    .S(_08272_),
    .X(_01997_));
 sg13g2_mux2_1 _26554_ (.A0(net4448),
    .A1(net6344),
    .S(_08272_),
    .X(_01998_));
 sg13g2_mux2_1 _26555_ (.A0(net4112),
    .A1(net6316),
    .S(_08272_),
    .X(_01999_));
 sg13g2_mux2_1 _26556_ (.A0(net4265),
    .A1(net6284),
    .S(_08272_),
    .X(_02000_));
 sg13g2_nand2_2 _26557_ (.Y(_08273_),
    .A(_03131_),
    .B(net5966));
 sg13g2_mux2_1 _26558_ (.A0(net6467),
    .A1(net6850),
    .S(_08273_),
    .X(_02001_));
 sg13g2_mux2_1 _26559_ (.A0(net6440),
    .A1(net6728),
    .S(_08273_),
    .X(_02002_));
 sg13g2_mux2_1 _26560_ (.A0(net6411),
    .A1(net4713),
    .S(_08273_),
    .X(_02003_));
 sg13g2_mux2_1 _26561_ (.A0(net6381),
    .A1(net4543),
    .S(_08273_),
    .X(_02004_));
 sg13g2_mux2_1 _26562_ (.A0(net6353),
    .A1(net6727),
    .S(_08273_),
    .X(_02005_));
 sg13g2_mux2_1 _26563_ (.A0(net6322),
    .A1(net6882),
    .S(_08273_),
    .X(_02006_));
 sg13g2_mux2_1 _26564_ (.A0(net6291),
    .A1(net6931),
    .S(_08273_),
    .X(_02007_));
 sg13g2_nor2_2 _26565_ (.A(_10126_),
    .B(_03130_),
    .Y(_08274_));
 sg13g2_nand2_2 _26566_ (.Y(_08275_),
    .A(_10125_),
    .B(_03129_));
 sg13g2_nand2_2 _26567_ (.Y(_08276_),
    .A(net5967),
    .B(_08274_));
 sg13g2_mux2_1 _26568_ (.A0(net6467),
    .A1(net7037),
    .S(_08276_),
    .X(_02008_));
 sg13g2_mux2_1 _26569_ (.A0(net6440),
    .A1(net6615),
    .S(_08276_),
    .X(_02009_));
 sg13g2_mux2_1 _26570_ (.A0(net6409),
    .A1(net6682),
    .S(_08276_),
    .X(_02010_));
 sg13g2_mux2_1 _26571_ (.A0(net6381),
    .A1(net6659),
    .S(_08276_),
    .X(_02011_));
 sg13g2_mux2_1 _26572_ (.A0(net6353),
    .A1(net4822),
    .S(_08276_),
    .X(_02012_));
 sg13g2_mux2_1 _26573_ (.A0(net6322),
    .A1(net6872),
    .S(_08276_),
    .X(_02013_));
 sg13g2_mux2_1 _26574_ (.A0(net6291),
    .A1(net7089),
    .S(_08276_),
    .X(_02014_));
 sg13g2_nand2_2 _26575_ (.Y(_08277_),
    .A(net5966),
    .B(_08245_));
 sg13g2_mux2_1 _26576_ (.A0(net6467),
    .A1(net6860),
    .S(_08277_),
    .X(_02015_));
 sg13g2_mux2_1 _26577_ (.A0(net6440),
    .A1(net7005),
    .S(_08277_),
    .X(_02016_));
 sg13g2_mux2_1 _26578_ (.A0(net6408),
    .A1(net6817),
    .S(_08277_),
    .X(_02017_));
 sg13g2_mux2_1 _26579_ (.A0(net6381),
    .A1(net6885),
    .S(_08277_),
    .X(_02018_));
 sg13g2_mux2_1 _26580_ (.A0(net6353),
    .A1(net6732),
    .S(_08277_),
    .X(_02019_));
 sg13g2_mux2_1 _26581_ (.A0(net6322),
    .A1(net6868),
    .S(_08277_),
    .X(_02020_));
 sg13g2_mux2_1 _26582_ (.A0(net6291),
    .A1(net6909),
    .S(_08277_),
    .X(_02021_));
 sg13g2_nor2b_2 _26583_ (.A(_10136_),
    .B_N(_06549_),
    .Y(_08278_));
 sg13g2_nand2b_2 _26584_ (.Y(_08279_),
    .B(_06549_),
    .A_N(_10136_));
 sg13g2_nand2_2 _26585_ (.Y(_08280_),
    .A(net5966),
    .B(_08278_));
 sg13g2_mux2_1 _26586_ (.A0(net6463),
    .A1(net4610),
    .S(_08280_),
    .X(_02022_));
 sg13g2_mux2_1 _26587_ (.A0(net6440),
    .A1(net6835),
    .S(_08280_),
    .X(_02023_));
 sg13g2_mux2_1 _26588_ (.A0(net6406),
    .A1(net4602),
    .S(_08280_),
    .X(_02024_));
 sg13g2_mux2_1 _26589_ (.A0(net6378),
    .A1(net6652),
    .S(_08280_),
    .X(_02025_));
 sg13g2_mux2_1 _26590_ (.A0(net6349),
    .A1(net4645),
    .S(_08280_),
    .X(_02026_));
 sg13g2_mux2_1 _26591_ (.A0(net6323),
    .A1(net4592),
    .S(_08280_),
    .X(_02027_));
 sg13g2_mux2_1 _26592_ (.A0(net6289),
    .A1(net4540),
    .S(_08280_),
    .X(_02028_));
 sg13g2_nor2_2 _26593_ (.A(_10069_),
    .B(_10126_),
    .Y(_08281_));
 sg13g2_nand2_2 _26594_ (.Y(_08282_),
    .A(net6028),
    .B(net5953));
 sg13g2_mux2_1 _26595_ (.A0(net6455),
    .A1(net4753),
    .S(_08282_),
    .X(_02029_));
 sg13g2_mux2_1 _26596_ (.A0(net6426),
    .A1(net6654),
    .S(_08282_),
    .X(_02030_));
 sg13g2_mux2_1 _26597_ (.A0(net6400),
    .A1(net4651),
    .S(_08282_),
    .X(_02031_));
 sg13g2_mux2_1 _26598_ (.A0(net6368),
    .A1(net4736),
    .S(_08282_),
    .X(_02032_));
 sg13g2_mux2_1 _26599_ (.A0(net6341),
    .A1(net4544),
    .S(_08282_),
    .X(_02033_));
 sg13g2_mux2_1 _26600_ (.A0(net6309),
    .A1(net6855),
    .S(_08282_),
    .X(_02034_));
 sg13g2_mux2_1 _26601_ (.A0(net6279),
    .A1(net6685),
    .S(_08282_),
    .X(_02035_));
 sg13g2_or2_2 _26602_ (.X(_08283_),
    .B(_10136_),
    .A(_10126_));
 sg13g2_nor2_2 _26603_ (.A(_08230_),
    .B(_08283_),
    .Y(_08284_));
 sg13g2_mux2_1 _26604_ (.A0(net3802),
    .A1(net6468),
    .S(_08284_),
    .X(_02036_));
 sg13g2_mux2_1 _26605_ (.A0(net3847),
    .A1(net6435),
    .S(_08284_),
    .X(_02037_));
 sg13g2_mux2_1 _26606_ (.A0(net4270),
    .A1(net6406),
    .S(_08284_),
    .X(_02038_));
 sg13g2_mux2_1 _26607_ (.A0(net4393),
    .A1(net6379),
    .S(_08284_),
    .X(_02039_));
 sg13g2_mux2_1 _26608_ (.A0(net4088),
    .A1(net6349),
    .S(_08284_),
    .X(_02040_));
 sg13g2_mux2_1 _26609_ (.A0(net3595),
    .A1(net6323),
    .S(_08284_),
    .X(_02041_));
 sg13g2_mux2_1 _26610_ (.A0(net4327),
    .A1(net6289),
    .S(_08284_),
    .X(_02042_));
 sg13g2_nor2_2 _26611_ (.A(net6030),
    .B(_08230_),
    .Y(_08285_));
 sg13g2_mux2_1 _26612_ (.A0(net3568),
    .A1(net6468),
    .S(_08285_),
    .X(_02043_));
 sg13g2_mux2_1 _26613_ (.A0(net3559),
    .A1(net6440),
    .S(_08285_),
    .X(_02044_));
 sg13g2_mux2_1 _26614_ (.A0(net4163),
    .A1(net6406),
    .S(_08285_),
    .X(_02045_));
 sg13g2_mux2_1 _26615_ (.A0(net4447),
    .A1(net6379),
    .S(_08285_),
    .X(_02046_));
 sg13g2_mux2_1 _26616_ (.A0(net3836),
    .A1(net6353),
    .S(_08285_),
    .X(_02047_));
 sg13g2_mux2_1 _26617_ (.A0(net4247),
    .A1(net6334),
    .S(_08285_),
    .X(_02048_));
 sg13g2_mux2_1 _26618_ (.A0(net3520),
    .A1(net6289),
    .S(_08285_),
    .X(_02049_));
 sg13g2_nand2_2 _26619_ (.Y(_08286_),
    .A(_06550_),
    .B(net5964));
 sg13g2_mux2_1 _26620_ (.A0(net6464),
    .A1(net4845),
    .S(_08286_),
    .X(_02050_));
 sg13g2_mux2_1 _26621_ (.A0(net6436),
    .A1(net4884),
    .S(_08286_),
    .X(_02051_));
 sg13g2_mux2_1 _26622_ (.A0(net6407),
    .A1(net6753),
    .S(_08286_),
    .X(_02052_));
 sg13g2_mux2_1 _26623_ (.A0(net6379),
    .A1(net4868),
    .S(_08286_),
    .X(_02053_));
 sg13g2_mux2_1 _26624_ (.A0(net6348),
    .A1(net6748),
    .S(_08286_),
    .X(_02054_));
 sg13g2_mux2_1 _26625_ (.A0(net6319),
    .A1(net6806),
    .S(_08286_),
    .X(_02055_));
 sg13g2_mux2_1 _26626_ (.A0(net6290),
    .A1(net6844),
    .S(_08286_),
    .X(_02056_));
 sg13g2_nand2_2 _26627_ (.Y(_08287_),
    .A(net5963),
    .B(_08241_));
 sg13g2_mux2_1 _26628_ (.A0(net6464),
    .A1(net4956),
    .S(_08287_),
    .X(_02057_));
 sg13g2_mux2_1 _26629_ (.A0(net6435),
    .A1(net6881),
    .S(_08287_),
    .X(_02058_));
 sg13g2_mux2_1 _26630_ (.A0(net6407),
    .A1(net4872),
    .S(_08287_),
    .X(_02059_));
 sg13g2_mux2_1 _26631_ (.A0(net6379),
    .A1(net6859),
    .S(_08287_),
    .X(_02060_));
 sg13g2_mux2_1 _26632_ (.A0(net6348),
    .A1(net4802),
    .S(_08287_),
    .X(_02061_));
 sg13g2_mux2_1 _26633_ (.A0(net6320),
    .A1(net4948),
    .S(_08287_),
    .X(_02062_));
 sg13g2_mux2_1 _26634_ (.A0(net6290),
    .A1(net4550),
    .S(_08287_),
    .X(_02063_));
 sg13g2_nand2_2 _26635_ (.Y(_08288_),
    .A(net5963),
    .B(_08281_));
 sg13g2_mux2_1 _26636_ (.A0(net6465),
    .A1(net6772),
    .S(_08288_),
    .X(_02064_));
 sg13g2_mux2_1 _26637_ (.A0(net6436),
    .A1(net6990),
    .S(_08288_),
    .X(_02065_));
 sg13g2_mux2_1 _26638_ (.A0(net6407),
    .A1(net6800),
    .S(_08288_),
    .X(_02066_));
 sg13g2_mux2_1 _26639_ (.A0(net6379),
    .A1(net4849),
    .S(_08288_),
    .X(_02067_));
 sg13g2_mux2_1 _26640_ (.A0(net6348),
    .A1(net6625),
    .S(_08288_),
    .X(_02068_));
 sg13g2_mux2_1 _26641_ (.A0(net6319),
    .A1(net4688),
    .S(_08288_),
    .X(_02069_));
 sg13g2_mux2_1 _26642_ (.A0(net6290),
    .A1(net6982),
    .S(_08288_),
    .X(_02070_));
 sg13g2_nand2_2 _26643_ (.Y(_08289_),
    .A(_08228_),
    .B(net5963));
 sg13g2_mux2_1 _26644_ (.A0(net6465),
    .A1(net4787),
    .S(_08289_),
    .X(_02071_));
 sg13g2_mux2_1 _26645_ (.A0(net6436),
    .A1(net4834),
    .S(_08289_),
    .X(_02072_));
 sg13g2_mux2_1 _26646_ (.A0(net6407),
    .A1(net6672),
    .S(_08289_),
    .X(_02073_));
 sg13g2_mux2_1 _26647_ (.A0(net6379),
    .A1(net4947),
    .S(_08289_),
    .X(_02074_));
 sg13g2_mux2_1 _26648_ (.A0(net6348),
    .A1(net6968),
    .S(_08289_),
    .X(_02075_));
 sg13g2_mux2_1 _26649_ (.A0(net6320),
    .A1(net6942),
    .S(_08289_),
    .X(_02076_));
 sg13g2_mux2_1 _26650_ (.A0(net6290),
    .A1(net4871),
    .S(_08289_),
    .X(_02077_));
 sg13g2_and2_2 _26651_ (.A(_06549_),
    .B(_08234_),
    .X(_08290_));
 sg13g2_nand2_2 _26652_ (.Y(_08291_),
    .A(net5963),
    .B(net5951));
 sg13g2_mux2_1 _26653_ (.A0(net6463),
    .A1(net4792),
    .S(_08291_),
    .X(_02078_));
 sg13g2_mux2_1 _26654_ (.A0(net6434),
    .A1(net6898),
    .S(_08291_),
    .X(_02079_));
 sg13g2_mux2_1 _26655_ (.A0(net6405),
    .A1(net4693),
    .S(_08291_),
    .X(_02080_));
 sg13g2_mux2_1 _26656_ (.A0(net6377),
    .A1(net4902),
    .S(_08291_),
    .X(_02081_));
 sg13g2_mux2_1 _26657_ (.A0(net6340),
    .A1(net4668),
    .S(_08291_),
    .X(_02082_));
 sg13g2_mux2_1 _26658_ (.A0(net6318),
    .A1(net6768),
    .S(_08291_),
    .X(_02083_));
 sg13g2_mux2_1 _26659_ (.A0(net6288),
    .A1(net6888),
    .S(_08291_),
    .X(_02084_));
 sg13g2_nand2_2 _26660_ (.Y(_08292_),
    .A(net5963),
    .B(_08251_));
 sg13g2_mux2_1 _26661_ (.A0(net6463),
    .A1(net6957),
    .S(_08292_),
    .X(_02085_));
 sg13g2_mux2_1 _26662_ (.A0(net6434),
    .A1(net7026),
    .S(_08292_),
    .X(_02086_));
 sg13g2_mux2_1 _26663_ (.A0(net6405),
    .A1(net6617),
    .S(_08292_),
    .X(_02087_));
 sg13g2_mux2_1 _26664_ (.A0(net6377),
    .A1(net4740),
    .S(_08292_),
    .X(_02088_));
 sg13g2_mux2_1 _26665_ (.A0(net6340),
    .A1(net4593),
    .S(_08292_),
    .X(_02089_));
 sg13g2_mux2_1 _26666_ (.A0(net6318),
    .A1(net4880),
    .S(_08292_),
    .X(_02090_));
 sg13g2_mux2_1 _26667_ (.A0(net6288),
    .A1(net6927),
    .S(_08292_),
    .X(_02091_));
 sg13g2_nor2_2 _26668_ (.A(_10126_),
    .B(_08235_),
    .Y(_08293_));
 sg13g2_nand2_2 _26669_ (.Y(_08294_),
    .A(_10125_),
    .B(_08234_));
 sg13g2_nand2_2 _26670_ (.Y(_08295_),
    .A(net5963),
    .B(_08293_));
 sg13g2_mux2_1 _26671_ (.A0(net6463),
    .A1(net6744),
    .S(_08295_),
    .X(_02092_));
 sg13g2_mux2_1 _26672_ (.A0(net6434),
    .A1(net7078),
    .S(_08295_),
    .X(_02093_));
 sg13g2_mux2_1 _26673_ (.A0(net6405),
    .A1(net6959),
    .S(_08295_),
    .X(_02094_));
 sg13g2_mux2_1 _26674_ (.A0(net6377),
    .A1(net6704),
    .S(_08295_),
    .X(_02095_));
 sg13g2_mux2_1 _26675_ (.A0(net6350),
    .A1(net7006),
    .S(_08295_),
    .X(_02096_));
 sg13g2_mux2_1 _26676_ (.A0(net6318),
    .A1(net7098),
    .S(_08295_),
    .X(_02097_));
 sg13g2_mux2_1 _26677_ (.A0(net6288),
    .A1(net4636),
    .S(_08295_),
    .X(_02098_));
 sg13g2_nand2_2 _26678_ (.Y(_08296_),
    .A(net6028),
    .B(net5968));
 sg13g2_mux2_1 _26679_ (.A0(net6455),
    .A1(net6858),
    .S(_08296_),
    .X(_02099_));
 sg13g2_mux2_1 _26680_ (.A0(net6426),
    .A1(net7011),
    .S(_08296_),
    .X(_02100_));
 sg13g2_mux2_1 _26681_ (.A0(net6400),
    .A1(net6693),
    .S(_08296_),
    .X(_02101_));
 sg13g2_mux2_1 _26682_ (.A0(net6369),
    .A1(net6757),
    .S(_08296_),
    .X(_02102_));
 sg13g2_mux2_1 _26683_ (.A0(net6341),
    .A1(net4633),
    .S(_08296_),
    .X(_02103_));
 sg13g2_mux2_1 _26684_ (.A0(net6309),
    .A1(net6905),
    .S(_08296_),
    .X(_02104_));
 sg13g2_mux2_1 _26685_ (.A0(net6279),
    .A1(net4796),
    .S(_08296_),
    .X(_02105_));
 sg13g2_and2_2 _26686_ (.A(_03129_),
    .B(_06549_),
    .X(_08297_));
 sg13g2_nand2_2 _26687_ (.Y(_08298_),
    .A(net5964),
    .B(net5950));
 sg13g2_mux2_1 _26688_ (.A0(net6455),
    .A1(net4637),
    .S(_08298_),
    .X(_02106_));
 sg13g2_mux2_1 _26689_ (.A0(net6430),
    .A1(net4931),
    .S(_08298_),
    .X(_02107_));
 sg13g2_mux2_1 _26690_ (.A0(net6398),
    .A1(net4930),
    .S(_08298_),
    .X(_02108_));
 sg13g2_mux2_1 _26691_ (.A0(net6369),
    .A1(net4759),
    .S(_08298_),
    .X(_02109_));
 sg13g2_mux2_1 _26692_ (.A0(net6340),
    .A1(net4560),
    .S(_08298_),
    .X(_02110_));
 sg13g2_mux2_1 _26693_ (.A0(net6309),
    .A1(net4894),
    .S(_08298_),
    .X(_02111_));
 sg13g2_mux2_1 _26694_ (.A0(net6281),
    .A1(net4388),
    .S(_08298_),
    .X(_02112_));
 sg13g2_nand2_2 _26695_ (.Y(_08299_),
    .A(_03131_),
    .B(net5964));
 sg13g2_mux2_1 _26696_ (.A0(net6455),
    .A1(net4778),
    .S(_08299_),
    .X(_02113_));
 sg13g2_mux2_1 _26697_ (.A0(net6434),
    .A1(net4883),
    .S(_08299_),
    .X(_02114_));
 sg13g2_mux2_1 _26698_ (.A0(net6398),
    .A1(net4934),
    .S(_08299_),
    .X(_02115_));
 sg13g2_mux2_1 _26699_ (.A0(net6369),
    .A1(net6923),
    .S(_08299_),
    .X(_02116_));
 sg13g2_mux2_1 _26700_ (.A0(net6340),
    .A1(net6914),
    .S(_08299_),
    .X(_02117_));
 sg13g2_mux2_1 _26701_ (.A0(net6309),
    .A1(net6667),
    .S(_08299_),
    .X(_02118_));
 sg13g2_mux2_1 _26702_ (.A0(net6281),
    .A1(net6808),
    .S(_08299_),
    .X(_02119_));
 sg13g2_nand2_2 _26703_ (.Y(_08300_),
    .A(net5964),
    .B(_08274_));
 sg13g2_mux2_1 _26704_ (.A0(net6455),
    .A1(net6866),
    .S(_08300_),
    .X(_02120_));
 sg13g2_mux2_1 _26705_ (.A0(net6434),
    .A1(net7010),
    .S(_08300_),
    .X(_02121_));
 sg13g2_mux2_1 _26706_ (.A0(net6398),
    .A1(net4582),
    .S(_08300_),
    .X(_02122_));
 sg13g2_mux2_1 _26707_ (.A0(net6368),
    .A1(net7027),
    .S(_08300_),
    .X(_02123_));
 sg13g2_mux2_1 _26708_ (.A0(net6340),
    .A1(net6830),
    .S(_08300_),
    .X(_02124_));
 sg13g2_mux2_1 _26709_ (.A0(net6309),
    .A1(net4777),
    .S(_08300_),
    .X(_02125_));
 sg13g2_mux2_1 _26710_ (.A0(net6281),
    .A1(net4375),
    .S(_08300_),
    .X(_02126_));
 sg13g2_nand2_2 _26711_ (.Y(_08301_),
    .A(net5964),
    .B(_08245_));
 sg13g2_mux2_1 _26712_ (.A0(net6455),
    .A1(net6730),
    .S(_08301_),
    .X(_02127_));
 sg13g2_mux2_1 _26713_ (.A0(net6434),
    .A1(net6926),
    .S(_08301_),
    .X(_02128_));
 sg13g2_mux2_1 _26714_ (.A0(net6398),
    .A1(net6803),
    .S(_08301_),
    .X(_02129_));
 sg13g2_mux2_1 _26715_ (.A0(net6369),
    .A1(net6848),
    .S(_08301_),
    .X(_02130_));
 sg13g2_mux2_1 _26716_ (.A0(net6340),
    .A1(net4726),
    .S(_08301_),
    .X(_02131_));
 sg13g2_mux2_1 _26717_ (.A0(net6309),
    .A1(net6895),
    .S(_08301_),
    .X(_02132_));
 sg13g2_mux2_1 _26718_ (.A0(net6288),
    .A1(net7062),
    .S(_08301_),
    .X(_02133_));
 sg13g2_nand2_2 _26719_ (.Y(_08302_),
    .A(net5963),
    .B(_08278_));
 sg13g2_mux2_1 _26720_ (.A0(net6464),
    .A1(net6599),
    .S(_08302_),
    .X(_02134_));
 sg13g2_mux2_1 _26721_ (.A0(net6436),
    .A1(net7047),
    .S(_08302_),
    .X(_02135_));
 sg13g2_mux2_1 _26722_ (.A0(net6413),
    .A1(net7042),
    .S(_08302_),
    .X(_02136_));
 sg13g2_mux2_1 _26723_ (.A0(net6377),
    .A1(net4638),
    .S(_08302_),
    .X(_02137_));
 sg13g2_mux2_1 _26724_ (.A0(net6348),
    .A1(net4800),
    .S(_08302_),
    .X(_02138_));
 sg13g2_mux2_1 _26725_ (.A0(net6318),
    .A1(net6600),
    .S(_08302_),
    .X(_02139_));
 sg13g2_mux2_1 _26726_ (.A0(net6288),
    .A1(net6724),
    .S(_08302_),
    .X(_02140_));
 sg13g2_nor2_2 _26727_ (.A(_08232_),
    .B(_08239_),
    .Y(_08303_));
 sg13g2_mux2_1 _26728_ (.A0(net4268),
    .A1(net6464),
    .S(_08303_),
    .X(_02141_));
 sg13g2_mux2_1 _26729_ (.A0(net4405),
    .A1(net6436),
    .S(_08303_),
    .X(_02142_));
 sg13g2_mux2_1 _26730_ (.A0(net3658),
    .A1(net6413),
    .S(_08303_),
    .X(_02143_));
 sg13g2_mux2_1 _26731_ (.A0(net3455),
    .A1(net6377),
    .S(_08303_),
    .X(_02144_));
 sg13g2_mux2_1 _26732_ (.A0(net4145),
    .A1(net6348),
    .S(_08303_),
    .X(_02145_));
 sg13g2_mux2_1 _26733_ (.A0(net3635),
    .A1(net6318),
    .S(_08303_),
    .X(_02146_));
 sg13g2_mux2_1 _26734_ (.A0(net3820),
    .A1(net6289),
    .S(_08303_),
    .X(_02147_));
 sg13g2_nor2_2 _26735_ (.A(_08239_),
    .B(_08283_),
    .Y(_08304_));
 sg13g2_mux2_1 _26736_ (.A0(net3448),
    .A1(net6464),
    .S(_08304_),
    .X(_02148_));
 sg13g2_mux2_1 _26737_ (.A0(net4019),
    .A1(net6436),
    .S(_08304_),
    .X(_02149_));
 sg13g2_mux2_1 _26738_ (.A0(net4225),
    .A1(net6407),
    .S(_08304_),
    .X(_02150_));
 sg13g2_mux2_1 _26739_ (.A0(net3932),
    .A1(net6377),
    .S(_08304_),
    .X(_02151_));
 sg13g2_mux2_1 _26740_ (.A0(net4115),
    .A1(net6348),
    .S(_08304_),
    .X(_02152_));
 sg13g2_mux2_1 _26741_ (.A0(net4150),
    .A1(net6318),
    .S(_08304_),
    .X(_02153_));
 sg13g2_mux2_1 _26742_ (.A0(net3560),
    .A1(net6288),
    .S(_08304_),
    .X(_02154_));
 sg13g2_nor2_2 _26743_ (.A(net6030),
    .B(_08239_),
    .Y(_08305_));
 sg13g2_mux2_1 _26744_ (.A0(net3945),
    .A1(net6464),
    .S(_08305_),
    .X(_02155_));
 sg13g2_mux2_1 _26745_ (.A0(net3877),
    .A1(net6435),
    .S(_08305_),
    .X(_02156_));
 sg13g2_mux2_1 _26746_ (.A0(net3710),
    .A1(net6407),
    .S(_08305_),
    .X(_02157_));
 sg13g2_mux2_1 _26747_ (.A0(net3930),
    .A1(net6377),
    .S(_08305_),
    .X(_02158_));
 sg13g2_mux2_1 _26748_ (.A0(net4357),
    .A1(net6348),
    .S(_08305_),
    .X(_02159_));
 sg13g2_mux2_1 _26749_ (.A0(net3875),
    .A1(net6318),
    .S(_08305_),
    .X(_02160_));
 sg13g2_mux2_1 _26750_ (.A0(net4006),
    .A1(net6288),
    .S(_08305_),
    .X(_02161_));
 sg13g2_nand2_2 _26751_ (.Y(_08306_),
    .A(net5969),
    .B(_08242_));
 sg13g2_mux2_1 _26752_ (.A0(net6457),
    .A1(net6907),
    .S(_08306_),
    .X(_02162_));
 sg13g2_mux2_1 _26753_ (.A0(net6428),
    .A1(net4815),
    .S(_08306_),
    .X(_02163_));
 sg13g2_mux2_1 _26754_ (.A0(net6399),
    .A1(net6819),
    .S(_08306_),
    .X(_02164_));
 sg13g2_mux2_1 _26755_ (.A0(net6370),
    .A1(net6871),
    .S(_08306_),
    .X(_02165_));
 sg13g2_mux2_1 _26756_ (.A0(net6342),
    .A1(net7061),
    .S(_08306_),
    .X(_02166_));
 sg13g2_mux2_1 _26757_ (.A0(net6311),
    .A1(net4739),
    .S(_08306_),
    .X(_02167_));
 sg13g2_mux2_1 _26758_ (.A0(net6280),
    .A1(net6932),
    .S(_08306_),
    .X(_02168_));
 sg13g2_nand2_2 _26759_ (.Y(_08307_),
    .A(net6027),
    .B(net5951));
 sg13g2_mux2_1 _26760_ (.A0(net6454),
    .A1(net4514),
    .S(_08307_),
    .X(_02169_));
 sg13g2_mux2_1 _26761_ (.A0(net6425),
    .A1(net4772),
    .S(_08307_),
    .X(_02170_));
 sg13g2_mux2_1 _26762_ (.A0(net6396),
    .A1(net7230),
    .S(_08307_),
    .X(_02171_));
 sg13g2_mux2_1 _26763_ (.A0(net6366),
    .A1(net6690),
    .S(_08307_),
    .X(_02172_));
 sg13g2_mux2_1 _26764_ (.A0(net6336),
    .A1(net4842),
    .S(_08307_),
    .X(_02173_));
 sg13g2_mux2_1 _26765_ (.A0(net6307),
    .A1(net6759),
    .S(_08307_),
    .X(_02174_));
 sg13g2_mux2_1 _26766_ (.A0(net6277),
    .A1(net6769),
    .S(_08307_),
    .X(_02175_));
 sg13g2_nand2_2 _26767_ (.Y(_08308_),
    .A(_08242_),
    .B(net5953));
 sg13g2_mux2_1 _26768_ (.A0(net6456),
    .A1(net7086),
    .S(_08308_),
    .X(_02176_));
 sg13g2_mux2_1 _26769_ (.A0(net6428),
    .A1(net4888),
    .S(_08308_),
    .X(_02177_));
 sg13g2_mux2_1 _26770_ (.A0(net6399),
    .A1(net4805),
    .S(_08308_),
    .X(_02178_));
 sg13g2_mux2_1 _26771_ (.A0(net6370),
    .A1(net4913),
    .S(_08308_),
    .X(_02179_));
 sg13g2_mux2_1 _26772_ (.A0(net6342),
    .A1(net4598),
    .S(_08308_),
    .X(_02180_));
 sg13g2_mux2_1 _26773_ (.A0(net6311),
    .A1(net4720),
    .S(_08308_),
    .X(_02181_));
 sg13g2_mux2_1 _26774_ (.A0(net6280),
    .A1(net4609),
    .S(_08308_),
    .X(_02182_));
 sg13g2_nor3_2 _26775_ (.A(_10069_),
    .B(net6067),
    .C(net6001),
    .Y(_08309_));
 sg13g2_mux2_1 _26776_ (.A0(net4067),
    .A1(net6457),
    .S(_08309_),
    .X(_02183_));
 sg13g2_mux2_1 _26777_ (.A0(net4147),
    .A1(net6428),
    .S(_08309_),
    .X(_02184_));
 sg13g2_mux2_1 _26778_ (.A0(net3909),
    .A1(net6400),
    .S(_08309_),
    .X(_02185_));
 sg13g2_mux2_1 _26779_ (.A0(net4096),
    .A1(net6370),
    .S(_08309_),
    .X(_02186_));
 sg13g2_mux2_1 _26780_ (.A0(net3499),
    .A1(net6342),
    .S(_08309_),
    .X(_02187_));
 sg13g2_mux2_1 _26781_ (.A0(net4385),
    .A1(net6311),
    .S(_08309_),
    .X(_02188_));
 sg13g2_mux2_1 _26782_ (.A0(net3576),
    .A1(net6280),
    .S(_08309_),
    .X(_02189_));
 sg13g2_nand2_2 _26783_ (.Y(_08310_),
    .A(_08242_),
    .B(net5951));
 sg13g2_mux2_1 _26784_ (.A0(net6465),
    .A1(net6829),
    .S(_08310_),
    .X(_02190_));
 sg13g2_mux2_1 _26785_ (.A0(net6443),
    .A1(net4561),
    .S(_08310_),
    .X(_02191_));
 sg13g2_mux2_1 _26786_ (.A0(net6414),
    .A1(net6595),
    .S(_08310_),
    .X(_02192_));
 sg13g2_mux2_1 _26787_ (.A0(net6371),
    .A1(net6790),
    .S(_08310_),
    .X(_02193_));
 sg13g2_mux2_1 _26788_ (.A0(net6346),
    .A1(net6934),
    .S(_08310_),
    .X(_02194_));
 sg13g2_mux2_1 _26789_ (.A0(net6327),
    .A1(net6747),
    .S(_08310_),
    .X(_02195_));
 sg13g2_mux2_1 _26790_ (.A0(net6296),
    .A1(net6771),
    .S(_08310_),
    .X(_02196_));
 sg13g2_nor2_2 _26791_ (.A(net6000),
    .B(_08252_),
    .Y(_08311_));
 sg13g2_mux2_1 _26792_ (.A0(net4243),
    .A1(net6465),
    .S(_08311_),
    .X(_02197_));
 sg13g2_mux2_1 _26793_ (.A0(net3556),
    .A1(net6443),
    .S(_08311_),
    .X(_02198_));
 sg13g2_mux2_1 _26794_ (.A0(net4000),
    .A1(net6414),
    .S(_08311_),
    .X(_02199_));
 sg13g2_mux2_1 _26795_ (.A0(net4258),
    .A1(net6371),
    .S(_08311_),
    .X(_02200_));
 sg13g2_mux2_1 _26796_ (.A0(net3464),
    .A1(net6346),
    .S(_08311_),
    .X(_02201_));
 sg13g2_mux2_1 _26797_ (.A0(net4052),
    .A1(net6320),
    .S(_08311_),
    .X(_02202_));
 sg13g2_mux2_1 _26798_ (.A0(net4068),
    .A1(net6296),
    .S(_08311_),
    .X(_02203_));
 sg13g2_nor2_2 _26799_ (.A(net6000),
    .B(_08294_),
    .Y(_08312_));
 sg13g2_mux2_1 _26800_ (.A0(net4094),
    .A1(net6464),
    .S(_08312_),
    .X(_02204_));
 sg13g2_mux2_1 _26801_ (.A0(net4406),
    .A1(net6443),
    .S(_08312_),
    .X(_02205_));
 sg13g2_mux2_1 _26802_ (.A0(net4383),
    .A1(net6414),
    .S(_08312_),
    .X(_02206_));
 sg13g2_mux2_1 _26803_ (.A0(net3524),
    .A1(net6371),
    .S(_08312_),
    .X(_02207_));
 sg13g2_mux2_1 _26804_ (.A0(net4314),
    .A1(net6358),
    .S(_08312_),
    .X(_02208_));
 sg13g2_mux2_1 _26805_ (.A0(net3461),
    .A1(net6320),
    .S(_08312_),
    .X(_02209_));
 sg13g2_mux2_1 _26806_ (.A0(net3612),
    .A1(net6296),
    .S(_08312_),
    .X(_02210_));
 sg13g2_nor2_2 _26807_ (.A(_08237_),
    .B(net6000),
    .Y(_08313_));
 sg13g2_mux2_1 _26808_ (.A0(net3795),
    .A1(net6464),
    .S(_08313_),
    .X(_02211_));
 sg13g2_mux2_1 _26809_ (.A0(net3925),
    .A1(net6443),
    .S(_08313_),
    .X(_02212_));
 sg13g2_mux2_1 _26810_ (.A0(net3621),
    .A1(net6414),
    .S(_08313_),
    .X(_02213_));
 sg13g2_mux2_1 _26811_ (.A0(net3916),
    .A1(net6371),
    .S(_08313_),
    .X(_02214_));
 sg13g2_mux2_1 _26812_ (.A0(net4193),
    .A1(net6358),
    .S(_08313_),
    .X(_02215_));
 sg13g2_mux2_1 _26813_ (.A0(net4036),
    .A1(net6320),
    .S(_08313_),
    .X(_02216_));
 sg13g2_mux2_1 _26814_ (.A0(net4178),
    .A1(net6296),
    .S(_08313_),
    .X(_02217_));
 sg13g2_nand2_2 _26815_ (.Y(_08314_),
    .A(_08242_),
    .B(net5950));
 sg13g2_mux2_1 _26816_ (.A0(net6458),
    .A1(net4953),
    .S(_08314_),
    .X(_02218_));
 sg13g2_mux2_1 _26817_ (.A0(net6427),
    .A1(net7031),
    .S(_08314_),
    .X(_02219_));
 sg13g2_mux2_1 _26818_ (.A0(net6403),
    .A1(net6805),
    .S(_08314_),
    .X(_02220_));
 sg13g2_mux2_1 _26819_ (.A0(net6370),
    .A1(net6822),
    .S(_08314_),
    .X(_02221_));
 sg13g2_mux2_1 _26820_ (.A0(net6346),
    .A1(net4776),
    .S(_08314_),
    .X(_02222_));
 sg13g2_mux2_1 _26821_ (.A0(net6311),
    .A1(net4876),
    .S(_08314_),
    .X(_02223_));
 sg13g2_mux2_1 _26822_ (.A0(net6280),
    .A1(net4769),
    .S(_08314_),
    .X(_02224_));
 sg13g2_nor2_2 _26823_ (.A(_03132_),
    .B(net6000),
    .Y(_08315_));
 sg13g2_mux2_1 _26824_ (.A0(net4082),
    .A1(net6458),
    .S(_08315_),
    .X(_02225_));
 sg13g2_mux2_1 _26825_ (.A0(net3783),
    .A1(net6427),
    .S(_08315_),
    .X(_02226_));
 sg13g2_mux2_1 _26826_ (.A0(net4058),
    .A1(net6402),
    .S(_08315_),
    .X(_02227_));
 sg13g2_mux2_1 _26827_ (.A0(net3592),
    .A1(net6370),
    .S(_08315_),
    .X(_02228_));
 sg13g2_mux2_1 _26828_ (.A0(net3933),
    .A1(net6342),
    .S(_08315_),
    .X(_02229_));
 sg13g2_mux2_1 _26829_ (.A0(net4180),
    .A1(net6311),
    .S(_08315_),
    .X(_02230_));
 sg13g2_mux2_1 _26830_ (.A0(net3685),
    .A1(net6280),
    .S(_08315_),
    .X(_02231_));
 sg13g2_nor2_2 _26831_ (.A(net6000),
    .B(_08275_),
    .Y(_08316_));
 sg13g2_mux2_1 _26832_ (.A0(net4377),
    .A1(net6457),
    .S(_08316_),
    .X(_02232_));
 sg13g2_mux2_1 _26833_ (.A0(net3730),
    .A1(net6427),
    .S(_08316_),
    .X(_02233_));
 sg13g2_mux2_1 _26834_ (.A0(net3490),
    .A1(net6402),
    .S(_08316_),
    .X(_02234_));
 sg13g2_mux2_1 _26835_ (.A0(net3790),
    .A1(net6375),
    .S(_08316_),
    .X(_02235_));
 sg13g2_mux2_1 _26836_ (.A0(net3599),
    .A1(net6346),
    .S(_08316_),
    .X(_02236_));
 sg13g2_mux2_1 _26837_ (.A0(net4354),
    .A1(net6312),
    .S(_08316_),
    .X(_02237_));
 sg13g2_mux2_1 _26838_ (.A0(net3830),
    .A1(net6280),
    .S(_08316_),
    .X(_02238_));
 sg13g2_nand2_2 _26839_ (.Y(_08317_),
    .A(net6027),
    .B(_08251_));
 sg13g2_mux2_1 _26840_ (.A0(net6454),
    .A1(net4729),
    .S(_08317_),
    .X(_02239_));
 sg13g2_mux2_1 _26841_ (.A0(net6425),
    .A1(net7000),
    .S(_08317_),
    .X(_02240_));
 sg13g2_mux2_1 _26842_ (.A0(net6397),
    .A1(net7045),
    .S(_08317_),
    .X(_02241_));
 sg13g2_mux2_1 _26843_ (.A0(net6366),
    .A1(net6588),
    .S(_08317_),
    .X(_02242_));
 sg13g2_mux2_1 _26844_ (.A0(net6335),
    .A1(net6750),
    .S(_08317_),
    .X(_02243_));
 sg13g2_mux2_1 _26845_ (.A0(net6307),
    .A1(net6886),
    .S(_08317_),
    .X(_02244_));
 sg13g2_mux2_1 _26846_ (.A0(net6277),
    .A1(net4533),
    .S(_08317_),
    .X(_02245_));
 sg13g2_nor2_2 _26847_ (.A(net6001),
    .B(_08279_),
    .Y(_08318_));
 sg13g2_mux2_1 _26848_ (.A0(net3601),
    .A1(net6456),
    .S(_08318_),
    .X(_02246_));
 sg13g2_mux2_1 _26849_ (.A0(net3687),
    .A1(net6429),
    .S(_08318_),
    .X(_02247_));
 sg13g2_mux2_1 _26850_ (.A0(net4153),
    .A1(net6398),
    .S(_08318_),
    .X(_02248_));
 sg13g2_mux2_1 _26851_ (.A0(net4226),
    .A1(net6371),
    .S(_08318_),
    .X(_02249_));
 sg13g2_mux2_1 _26852_ (.A0(net3518),
    .A1(net6341),
    .S(_08318_),
    .X(_02250_));
 sg13g2_mux2_1 _26853_ (.A0(net4001),
    .A1(net6311),
    .S(_08318_),
    .X(_02251_));
 sg13g2_mux2_1 _26854_ (.A0(net3897),
    .A1(net6281),
    .S(_08318_),
    .X(_02252_));
 sg13g2_nor2_2 _26855_ (.A(_08232_),
    .B(net6001),
    .Y(_08319_));
 sg13g2_mux2_1 _26856_ (.A0(net3734),
    .A1(net6458),
    .S(_08319_),
    .X(_02253_));
 sg13g2_mux2_1 _26857_ (.A0(net3984),
    .A1(net6429),
    .S(_08319_),
    .X(_02254_));
 sg13g2_mux2_1 _26858_ (.A0(net3911),
    .A1(net6399),
    .S(_08319_),
    .X(_02255_));
 sg13g2_mux2_1 _26859_ (.A0(net3512),
    .A1(net6371),
    .S(_08319_),
    .X(_02256_));
 sg13g2_mux2_1 _26860_ (.A0(net3946),
    .A1(net6340),
    .S(_08319_),
    .X(_02257_));
 sg13g2_mux2_1 _26861_ (.A0(net3566),
    .A1(net6320),
    .S(_08319_),
    .X(_02258_));
 sg13g2_mux2_1 _26862_ (.A0(net4040),
    .A1(net6305),
    .S(_08319_),
    .X(_02259_));
 sg13g2_nor2_2 _26863_ (.A(net6000),
    .B(net5952),
    .Y(_08320_));
 sg13g2_mux2_1 _26864_ (.A0(net4035),
    .A1(net6455),
    .S(_08320_),
    .X(_02260_));
 sg13g2_mux2_1 _26865_ (.A0(net3500),
    .A1(net6429),
    .S(_08320_),
    .X(_02261_));
 sg13g2_mux2_1 _26866_ (.A0(net4334),
    .A1(net6398),
    .S(_08320_),
    .X(_02262_));
 sg13g2_mux2_1 _26867_ (.A0(net3803),
    .A1(net6371),
    .S(_08320_),
    .X(_02263_));
 sg13g2_mux2_1 _26868_ (.A0(net4326),
    .A1(net6341),
    .S(_08320_),
    .X(_02264_));
 sg13g2_mux2_1 _26869_ (.A0(net3622),
    .A1(net6311),
    .S(_08320_),
    .X(_02265_));
 sg13g2_mux2_1 _26870_ (.A0(net3467),
    .A1(net6281),
    .S(_08320_),
    .X(_02266_));
 sg13g2_nor2_2 _26871_ (.A(net6030),
    .B(net6000),
    .Y(_08321_));
 sg13g2_mux2_1 _26872_ (.A0(net3742),
    .A1(net6463),
    .S(_08321_),
    .X(_02267_));
 sg13g2_mux2_1 _26873_ (.A0(net3614),
    .A1(net6429),
    .S(_08321_),
    .X(_02268_));
 sg13g2_mux2_1 _26874_ (.A0(net4267),
    .A1(net6399),
    .S(_08321_),
    .X(_02269_));
 sg13g2_mux2_1 _26875_ (.A0(net3917),
    .A1(net6371),
    .S(_08321_),
    .X(_02270_));
 sg13g2_mux2_1 _26876_ (.A0(net3853),
    .A1(net6340),
    .S(_08321_),
    .X(_02271_));
 sg13g2_mux2_1 _26877_ (.A0(net3648),
    .A1(net6320),
    .S(_08321_),
    .X(_02272_));
 sg13g2_mux2_1 _26878_ (.A0(net4138),
    .A1(net6290),
    .S(_08321_),
    .X(_02273_));
 sg13g2_nand2_2 _26879_ (.Y(_08322_),
    .A(_06550_),
    .B(net5961));
 sg13g2_mux2_1 _26880_ (.A0(net6470),
    .A1(net7002),
    .S(_08322_),
    .X(_02274_));
 sg13g2_mux2_1 _26881_ (.A0(net6441),
    .A1(net4765),
    .S(_08322_),
    .X(_02275_));
 sg13g2_mux2_1 _26882_ (.A0(net6410),
    .A1(net6922),
    .S(_08322_),
    .X(_02276_));
 sg13g2_mux2_1 _26883_ (.A0(net6384),
    .A1(net4468),
    .S(_08322_),
    .X(_02277_));
 sg13g2_mux2_1 _26884_ (.A0(net6354),
    .A1(net4500),
    .S(_08322_),
    .X(_02278_));
 sg13g2_mux2_1 _26885_ (.A0(net6330),
    .A1(net6912),
    .S(_08322_),
    .X(_02279_));
 sg13g2_mux2_1 _26886_ (.A0(net6294),
    .A1(net4945),
    .S(_08322_),
    .X(_02280_));
 sg13g2_nand2_2 _26887_ (.Y(_08323_),
    .A(net5962),
    .B(net5961));
 sg13g2_mux2_1 _26888_ (.A0(net6469),
    .A1(net4927),
    .S(_08323_),
    .X(_02281_));
 sg13g2_mux2_1 _26889_ (.A0(net6446),
    .A1(net4912),
    .S(_08323_),
    .X(_02282_));
 sg13g2_mux2_1 _26890_ (.A0(net6410),
    .A1(net6719),
    .S(_08323_),
    .X(_02283_));
 sg13g2_mux2_1 _26891_ (.A0(net6391),
    .A1(net4721),
    .S(_08323_),
    .X(_02284_));
 sg13g2_mux2_1 _26892_ (.A0(net6354),
    .A1(net4725),
    .S(_08323_),
    .X(_02285_));
 sg13g2_mux2_1 _26893_ (.A0(net6330),
    .A1(net7135),
    .S(_08323_),
    .X(_02286_));
 sg13g2_mux2_1 _26894_ (.A0(net6294),
    .A1(net6969),
    .S(_08323_),
    .X(_02287_));
 sg13g2_nand2_2 _26895_ (.Y(_08324_),
    .A(net5961),
    .B(net5953));
 sg13g2_mux2_1 _26896_ (.A0(net6469),
    .A1(net6951),
    .S(_08324_),
    .X(_02288_));
 sg13g2_mux2_1 _26897_ (.A0(net6441),
    .A1(net4951),
    .S(_08324_),
    .X(_02289_));
 sg13g2_mux2_1 _26898_ (.A0(net6410),
    .A1(net4768),
    .S(_08324_),
    .X(_02290_));
 sg13g2_mux2_1 _26899_ (.A0(net6383),
    .A1(net4524),
    .S(_08324_),
    .X(_02291_));
 sg13g2_mux2_1 _26900_ (.A0(net6354),
    .A1(net6614),
    .S(_08324_),
    .X(_02292_));
 sg13g2_mux2_1 _26901_ (.A0(net6325),
    .A1(net6856),
    .S(_08324_),
    .X(_02293_));
 sg13g2_mux2_1 _26902_ (.A0(net6294),
    .A1(net4521),
    .S(_08324_),
    .X(_02294_));
 sg13g2_nand2_2 _26903_ (.Y(_08325_),
    .A(net5968),
    .B(net5961));
 sg13g2_mux2_1 _26904_ (.A0(net6469),
    .A1(net4751),
    .S(_08325_),
    .X(_02295_));
 sg13g2_mux2_1 _26905_ (.A0(net6441),
    .A1(net4597),
    .S(_08325_),
    .X(_02296_));
 sg13g2_mux2_1 _26906_ (.A0(net6410),
    .A1(net4957),
    .S(_08325_),
    .X(_02297_));
 sg13g2_mux2_1 _26907_ (.A0(net6383),
    .A1(net4516),
    .S(_08325_),
    .X(_02298_));
 sg13g2_mux2_1 _26908_ (.A0(net6354),
    .A1(net6836),
    .S(_08325_),
    .X(_02299_));
 sg13g2_mux2_1 _26909_ (.A0(net6325),
    .A1(net6609),
    .S(_08325_),
    .X(_02300_));
 sg13g2_mux2_1 _26910_ (.A0(net6294),
    .A1(net6689),
    .S(_08325_),
    .X(_02301_));
 sg13g2_nand2_2 _26911_ (.Y(_08326_),
    .A(net5960),
    .B(_08290_));
 sg13g2_mux2_1 _26912_ (.A0(net6471),
    .A1(net6892),
    .S(_08326_),
    .X(_02302_));
 sg13g2_mux2_1 _26913_ (.A0(net6439),
    .A1(net6899),
    .S(_08326_),
    .X(_02303_));
 sg13g2_mux2_1 _26914_ (.A0(net6412),
    .A1(net4708),
    .S(_08326_),
    .X(_02304_));
 sg13g2_mux2_1 _26915_ (.A0(net6382),
    .A1(net4890),
    .S(_08326_),
    .X(_02305_));
 sg13g2_mux2_1 _26916_ (.A0(net6352),
    .A1(net6611),
    .S(_08326_),
    .X(_02306_));
 sg13g2_mux2_1 _26917_ (.A0(net6324),
    .A1(net4541),
    .S(_08326_),
    .X(_02307_));
 sg13g2_mux2_1 _26918_ (.A0(net6292),
    .A1(net4803),
    .S(_08326_),
    .X(_02308_));
 sg13g2_nand2_2 _26919_ (.Y(_08327_),
    .A(net6027),
    .B(_08293_));
 sg13g2_mux2_1 _26920_ (.A0(net6454),
    .A1(net6751),
    .S(_08327_),
    .X(_02309_));
 sg13g2_mux2_1 _26921_ (.A0(net6425),
    .A1(net6723),
    .S(_08327_),
    .X(_02310_));
 sg13g2_mux2_1 _26922_ (.A0(net6397),
    .A1(net4605),
    .S(_08327_),
    .X(_02311_));
 sg13g2_mux2_1 _26923_ (.A0(net6366),
    .A1(net6714),
    .S(_08327_),
    .X(_02312_));
 sg13g2_mux2_1 _26924_ (.A0(net6335),
    .A1(net7066),
    .S(_08327_),
    .X(_02313_));
 sg13g2_mux2_1 _26925_ (.A0(net6307),
    .A1(net4896),
    .S(_08327_),
    .X(_02314_));
 sg13g2_mux2_1 _26926_ (.A0(net6277),
    .A1(net4621),
    .S(_08327_),
    .X(_02315_));
 sg13g2_nand2_2 _26927_ (.Y(_08328_),
    .A(net5960),
    .B(_08293_));
 sg13g2_mux2_1 _26928_ (.A0(net6468),
    .A1(net6936),
    .S(_08328_),
    .X(_02316_));
 sg13g2_mux2_1 _26929_ (.A0(net6439),
    .A1(net4774),
    .S(_08328_),
    .X(_02317_));
 sg13g2_mux2_1 _26930_ (.A0(net6408),
    .A1(net6584),
    .S(_08328_),
    .X(_02318_));
 sg13g2_mux2_1 _26931_ (.A0(net6382),
    .A1(net6703),
    .S(_08328_),
    .X(_02319_));
 sg13g2_mux2_1 _26932_ (.A0(net6352),
    .A1(net6683),
    .S(_08328_),
    .X(_02320_));
 sg13g2_mux2_1 _26933_ (.A0(net6324),
    .A1(net4943),
    .S(_08328_),
    .X(_02321_));
 sg13g2_mux2_1 _26934_ (.A0(net6292),
    .A1(net6756),
    .S(_08328_),
    .X(_02322_));
 sg13g2_nand2_2 _26935_ (.Y(_08329_),
    .A(_08236_),
    .B(net5960));
 sg13g2_mux2_1 _26936_ (.A0(net6468),
    .A1(net6828),
    .S(_08329_),
    .X(_02323_));
 sg13g2_mux2_1 _26937_ (.A0(net6439),
    .A1(net6862),
    .S(_08329_),
    .X(_02324_));
 sg13g2_mux2_1 _26938_ (.A0(net6408),
    .A1(net4781),
    .S(_08329_),
    .X(_02325_));
 sg13g2_mux2_1 _26939_ (.A0(net6382),
    .A1(net4650),
    .S(_08329_),
    .X(_02326_));
 sg13g2_mux2_1 _26940_ (.A0(net6351),
    .A1(net4684),
    .S(_08329_),
    .X(_02327_));
 sg13g2_mux2_1 _26941_ (.A0(net6324),
    .A1(net6986),
    .S(_08329_),
    .X(_02328_));
 sg13g2_mux2_1 _26942_ (.A0(net6292),
    .A1(net4583),
    .S(_08329_),
    .X(_02329_));
 sg13g2_nand2_2 _26943_ (.Y(_08330_),
    .A(net5960),
    .B(_08297_));
 sg13g2_mux2_1 _26944_ (.A0(net6468),
    .A1(net6736),
    .S(_08330_),
    .X(_02330_));
 sg13g2_mux2_1 _26945_ (.A0(net6438),
    .A1(net6738),
    .S(_08330_),
    .X(_02331_));
 sg13g2_mux2_1 _26946_ (.A0(net6409),
    .A1(net4589),
    .S(_08330_),
    .X(_02332_));
 sg13g2_mux2_1 _26947_ (.A0(net6382),
    .A1(net6602),
    .S(_08330_),
    .X(_02333_));
 sg13g2_mux2_1 _26948_ (.A0(net6352),
    .A1(net6722),
    .S(_08330_),
    .X(_02334_));
 sg13g2_mux2_1 _26949_ (.A0(net6323),
    .A1(net4675),
    .S(_08330_),
    .X(_02335_));
 sg13g2_mux2_1 _26950_ (.A0(net6294),
    .A1(net6623),
    .S(_08330_),
    .X(_02336_));
 sg13g2_nand2_2 _26951_ (.Y(_08331_),
    .A(_03131_),
    .B(net5960));
 sg13g2_mux2_1 _26952_ (.A0(net6469),
    .A1(net6875),
    .S(_08331_),
    .X(_02337_));
 sg13g2_mux2_1 _26953_ (.A0(net6438),
    .A1(net4928),
    .S(_08331_),
    .X(_02338_));
 sg13g2_mux2_1 _26954_ (.A0(net6409),
    .A1(net6869),
    .S(_08331_),
    .X(_02339_));
 sg13g2_mux2_1 _26955_ (.A0(net6382),
    .A1(net7017),
    .S(_08331_),
    .X(_02340_));
 sg13g2_mux2_1 _26956_ (.A0(net6351),
    .A1(net4892),
    .S(_08331_),
    .X(_02341_));
 sg13g2_mux2_1 _26957_ (.A0(net6323),
    .A1(net6777),
    .S(_08331_),
    .X(_02342_));
 sg13g2_mux2_1 _26958_ (.A0(net6294),
    .A1(net4564),
    .S(_08331_),
    .X(_02343_));
 sg13g2_nand2_2 _26959_ (.Y(_08332_),
    .A(net5960),
    .B(_08274_));
 sg13g2_mux2_1 _26960_ (.A0(net6468),
    .A1(net6870),
    .S(_08332_),
    .X(_02344_));
 sg13g2_mux2_1 _26961_ (.A0(net6438),
    .A1(net6658),
    .S(_08332_),
    .X(_02345_));
 sg13g2_mux2_1 _26962_ (.A0(net6409),
    .A1(net7082),
    .S(_08332_),
    .X(_02346_));
 sg13g2_mux2_1 _26963_ (.A0(net6382),
    .A1(net6787),
    .S(_08332_),
    .X(_02347_));
 sg13g2_mux2_1 _26964_ (.A0(net6351),
    .A1(net4577),
    .S(_08332_),
    .X(_02348_));
 sg13g2_mux2_1 _26965_ (.A0(net6323),
    .A1(net6811),
    .S(_08332_),
    .X(_02349_));
 sg13g2_mux2_1 _26966_ (.A0(net6294),
    .A1(net6976),
    .S(_08332_),
    .X(_02350_));
 sg13g2_nand2_2 _26967_ (.Y(_08333_),
    .A(_08245_),
    .B(net5960));
 sg13g2_mux2_1 _26968_ (.A0(net6468),
    .A1(net6742),
    .S(_08333_),
    .X(_02351_));
 sg13g2_mux2_1 _26969_ (.A0(net6438),
    .A1(net4851),
    .S(_08333_),
    .X(_02352_));
 sg13g2_mux2_1 _26970_ (.A0(net6410),
    .A1(net6720),
    .S(_08333_),
    .X(_02353_));
 sg13g2_mux2_1 _26971_ (.A0(net6382),
    .A1(net4714),
    .S(_08333_),
    .X(_02354_));
 sg13g2_mux2_1 _26972_ (.A0(net6351),
    .A1(net4659),
    .S(_08333_),
    .X(_02355_));
 sg13g2_mux2_1 _26973_ (.A0(net6323),
    .A1(net6943),
    .S(_08333_),
    .X(_02356_));
 sg13g2_mux2_1 _26974_ (.A0(net6294),
    .A1(net6863),
    .S(_08333_),
    .X(_02357_));
 sg13g2_nand2_2 _26975_ (.Y(_08334_),
    .A(net5961),
    .B(_08278_));
 sg13g2_mux2_1 _26976_ (.A0(net6469),
    .A1(net6960),
    .S(_08334_),
    .X(_02358_));
 sg13g2_mux2_1 _26977_ (.A0(net6440),
    .A1(net4567),
    .S(_08334_),
    .X(_02359_));
 sg13g2_mux2_1 _26978_ (.A0(net6409),
    .A1(net4502),
    .S(_08334_),
    .X(_02360_));
 sg13g2_mux2_1 _26979_ (.A0(net6383),
    .A1(net4755),
    .S(_08334_),
    .X(_02361_));
 sg13g2_mux2_1 _26980_ (.A0(net6353),
    .A1(net4475),
    .S(_08334_),
    .X(_02362_));
 sg13g2_mux2_1 _26981_ (.A0(net6325),
    .A1(net4555),
    .S(_08334_),
    .X(_02363_));
 sg13g2_mux2_1 _26982_ (.A0(net6293),
    .A1(net6733),
    .S(_08334_),
    .X(_02364_));
 sg13g2_nor2b_2 _26983_ (.A(net5965),
    .B_N(net5961),
    .Y(_08335_));
 sg13g2_mux2_1 _26984_ (.A0(net3838),
    .A1(net6469),
    .S(_08335_),
    .X(_02365_));
 sg13g2_mux2_1 _26985_ (.A0(net3796),
    .A1(net6440),
    .S(_08335_),
    .X(_02366_));
 sg13g2_mux2_1 _26986_ (.A0(net3454),
    .A1(net6409),
    .S(_08335_),
    .X(_02367_));
 sg13g2_mux2_1 _26987_ (.A0(net3937),
    .A1(net6383),
    .S(_08335_),
    .X(_02368_));
 sg13g2_mux2_1 _26988_ (.A0(net4097),
    .A1(net6353),
    .S(_08335_),
    .X(_02369_));
 sg13g2_mux2_1 _26989_ (.A0(net3494),
    .A1(net6325),
    .S(_08335_),
    .X(_02370_));
 sg13g2_mux2_1 _26990_ (.A0(net4389),
    .A1(net6293),
    .S(_08335_),
    .X(_02371_));
 sg13g2_nor3_2 _26991_ (.A(_10002_),
    .B(_08249_),
    .C(net5952),
    .Y(_08336_));
 sg13g2_mux2_1 _26992_ (.A0(net3766),
    .A1(net6469),
    .S(_08336_),
    .X(_02372_));
 sg13g2_mux2_1 _26993_ (.A0(net4044),
    .A1(net6441),
    .S(_08336_),
    .X(_02373_));
 sg13g2_mux2_1 _26994_ (.A0(net3468),
    .A1(net6409),
    .S(_08336_),
    .X(_02374_));
 sg13g2_mux2_1 _26995_ (.A0(net3570),
    .A1(net6383),
    .S(_08336_),
    .X(_02375_));
 sg13g2_mux2_1 _26996_ (.A0(net3625),
    .A1(net6354),
    .S(_08336_),
    .X(_02376_));
 sg13g2_mux2_1 _26997_ (.A0(net3833),
    .A1(net6325),
    .S(_08336_),
    .X(_02377_));
 sg13g2_mux2_1 _26998_ (.A0(net4013),
    .A1(net6293),
    .S(_08336_),
    .X(_02378_));
 sg13g2_nand2_2 _26999_ (.Y(_08337_),
    .A(net6027),
    .B(_08236_));
 sg13g2_mux2_1 _27000_ (.A0(net6454),
    .A1(net4615),
    .S(_08337_),
    .X(_02379_));
 sg13g2_mux2_1 _27001_ (.A0(net6425),
    .A1(net4661),
    .S(_08337_),
    .X(_02380_));
 sg13g2_mux2_1 _27002_ (.A0(net6397),
    .A1(net6783),
    .S(_08337_),
    .X(_02381_));
 sg13g2_mux2_1 _27003_ (.A0(net6366),
    .A1(net6766),
    .S(_08337_),
    .X(_02382_));
 sg13g2_mux2_1 _27004_ (.A0(net6335),
    .A1(net7134),
    .S(_08337_),
    .X(_02383_));
 sg13g2_mux2_1 _27005_ (.A0(net6306),
    .A1(net4578),
    .S(_08337_),
    .X(_02384_));
 sg13g2_mux2_1 _27006_ (.A0(net6277),
    .A1(net4862),
    .S(_08337_),
    .X(_02385_));
 sg13g2_nand2_2 _27007_ (.Y(_08338_),
    .A(_06550_),
    .B(_08255_));
 sg13g2_mux2_1 _27008_ (.A0(net6477),
    .A1(net6616),
    .S(_08338_),
    .X(_02386_));
 sg13g2_mux2_1 _27009_ (.A0(net6448),
    .A1(net6827),
    .S(_08338_),
    .X(_02387_));
 sg13g2_mux2_1 _27010_ (.A0(net6418),
    .A1(net4485),
    .S(_08338_),
    .X(_02388_));
 sg13g2_mux2_1 _27011_ (.A0(net6388),
    .A1(net4861),
    .S(_08338_),
    .X(_02389_));
 sg13g2_mux2_1 _27012_ (.A0(net6360),
    .A1(net4881),
    .S(_08338_),
    .X(_02390_));
 sg13g2_mux2_1 _27013_ (.A0(net6330),
    .A1(net4612),
    .S(_08338_),
    .X(_02391_));
 sg13g2_mux2_1 _27014_ (.A0(net6300),
    .A1(net4932),
    .S(_08338_),
    .X(_02392_));
 sg13g2_nand2_2 _27015_ (.Y(_08339_),
    .A(net5962),
    .B(_08255_));
 sg13g2_mux2_1 _27016_ (.A0(net6477),
    .A1(net4594),
    .S(_08339_),
    .X(_02393_));
 sg13g2_mux2_1 _27017_ (.A0(net6448),
    .A1(net4914),
    .S(_08339_),
    .X(_02394_));
 sg13g2_mux2_1 _27018_ (.A0(net6418),
    .A1(net6799),
    .S(_08339_),
    .X(_02395_));
 sg13g2_mux2_1 _27019_ (.A0(net6388),
    .A1(net4797),
    .S(_08339_),
    .X(_02396_));
 sg13g2_mux2_1 _27020_ (.A0(net6360),
    .A1(net4719),
    .S(_08339_),
    .X(_02397_));
 sg13g2_mux2_1 _27021_ (.A0(net6330),
    .A1(net6688),
    .S(_08339_),
    .X(_02398_));
 sg13g2_mux2_1 _27022_ (.A0(net6300),
    .A1(net7020),
    .S(_08339_),
    .X(_02399_));
 sg13g2_nand2_2 _27023_ (.Y(_08340_),
    .A(_08255_),
    .B(net5953));
 sg13g2_mux2_1 _27024_ (.A0(net6477),
    .A1(net6937),
    .S(_08340_),
    .X(_02400_));
 sg13g2_mux2_1 _27025_ (.A0(net6448),
    .A1(net4794),
    .S(_08340_),
    .X(_02401_));
 sg13g2_mux2_1 _27026_ (.A0(net6418),
    .A1(net4529),
    .S(_08340_),
    .X(_02402_));
 sg13g2_mux2_1 _27027_ (.A0(net6388),
    .A1(net4552),
    .S(_08340_),
    .X(_02403_));
 sg13g2_mux2_1 _27028_ (.A0(net6360),
    .A1(net6883),
    .S(_08340_),
    .X(_02404_));
 sg13g2_mux2_1 _27029_ (.A0(net6330),
    .A1(net4507),
    .S(_08340_),
    .X(_02405_));
 sg13g2_mux2_1 _27030_ (.A0(net6300),
    .A1(net6833),
    .S(_08340_),
    .X(_02406_));
 sg13g2_nand2_2 _27031_ (.Y(_08341_),
    .A(net5968),
    .B(_08255_));
 sg13g2_mux2_1 _27032_ (.A0(net6477),
    .A1(net7106),
    .S(_08341_),
    .X(_02407_));
 sg13g2_mux2_1 _27033_ (.A0(net6446),
    .A1(net4562),
    .S(_08341_),
    .X(_02408_));
 sg13g2_mux2_1 _27034_ (.A0(net6418),
    .A1(net4806),
    .S(_08341_),
    .X(_02409_));
 sg13g2_mux2_1 _27035_ (.A0(net6388),
    .A1(net4559),
    .S(_08341_),
    .X(_02410_));
 sg13g2_mux2_1 _27036_ (.A0(net6359),
    .A1(net4604),
    .S(_08341_),
    .X(_02411_));
 sg13g2_mux2_1 _27037_ (.A0(net6330),
    .A1(net4939),
    .S(_08341_),
    .X(_02412_));
 sg13g2_mux2_1 _27038_ (.A0(net6300),
    .A1(net6798),
    .S(_08341_),
    .X(_02413_));
 sg13g2_nand2_2 _27039_ (.Y(_08342_),
    .A(_08255_),
    .B(net5951));
 sg13g2_mux2_1 _27040_ (.A0(net6476),
    .A1(net6665),
    .S(_08342_),
    .X(_02414_));
 sg13g2_mux2_1 _27041_ (.A0(net6449),
    .A1(net6884),
    .S(_08342_),
    .X(_02415_));
 sg13g2_mux2_1 _27042_ (.A0(net6420),
    .A1(net6711),
    .S(_08342_),
    .X(_02416_));
 sg13g2_mux2_1 _27043_ (.A0(net6389),
    .A1(net6978),
    .S(_08342_),
    .X(_02417_));
 sg13g2_mux2_1 _27044_ (.A0(net6362),
    .A1(net4622),
    .S(_08342_),
    .X(_02418_));
 sg13g2_mux2_1 _27045_ (.A0(net6332),
    .A1(net6972),
    .S(_08342_),
    .X(_02419_));
 sg13g2_mux2_1 _27046_ (.A0(net6302),
    .A1(net4694),
    .S(_08342_),
    .X(_02420_));
 sg13g2_nor2_2 _27047_ (.A(_08252_),
    .B(net5959),
    .Y(_08343_));
 sg13g2_mux2_1 _27048_ (.A0(net4349),
    .A1(net6476),
    .S(_08343_),
    .X(_02421_));
 sg13g2_mux2_1 _27049_ (.A0(net4018),
    .A1(net6449),
    .S(_08343_),
    .X(_02422_));
 sg13g2_mux2_1 _27050_ (.A0(net4331),
    .A1(net6419),
    .S(_08343_),
    .X(_02423_));
 sg13g2_mux2_1 _27051_ (.A0(net3850),
    .A1(net6389),
    .S(_08343_),
    .X(_02424_));
 sg13g2_mux2_1 _27052_ (.A0(net3691),
    .A1(net6362),
    .S(_08343_),
    .X(_02425_));
 sg13g2_mux2_1 _27053_ (.A0(net3677),
    .A1(net6332),
    .S(_08343_),
    .X(_02426_));
 sg13g2_mux2_1 _27054_ (.A0(net4248),
    .A1(net6302),
    .S(_08343_),
    .X(_02427_));
 sg13g2_nor2_2 _27055_ (.A(net5959),
    .B(_08294_),
    .Y(_08344_));
 sg13g2_mux2_1 _27056_ (.A0(net4169),
    .A1(net6476),
    .S(_08344_),
    .X(_02428_));
 sg13g2_mux2_1 _27057_ (.A0(net4005),
    .A1(net6449),
    .S(_08344_),
    .X(_02429_));
 sg13g2_mux2_1 _27058_ (.A0(net4134),
    .A1(net6419),
    .S(_08344_),
    .X(_02430_));
 sg13g2_mux2_1 _27059_ (.A0(net4204),
    .A1(net6389),
    .S(_08344_),
    .X(_02431_));
 sg13g2_mux2_1 _27060_ (.A0(net4266),
    .A1(net6362),
    .S(_08344_),
    .X(_02432_));
 sg13g2_mux2_1 _27061_ (.A0(net3935),
    .A1(net6332),
    .S(_08344_),
    .X(_02433_));
 sg13g2_mux2_1 _27062_ (.A0(net4050),
    .A1(net6302),
    .S(_08344_),
    .X(_02434_));
 sg13g2_nor2_2 _27063_ (.A(_08237_),
    .B(net5959),
    .Y(_08345_));
 sg13g2_mux2_1 _27064_ (.A0(net4162),
    .A1(net6476),
    .S(_08345_),
    .X(_02435_));
 sg13g2_mux2_1 _27065_ (.A0(net4120),
    .A1(net6449),
    .S(_08345_),
    .X(_02436_));
 sg13g2_mux2_1 _27066_ (.A0(net4348),
    .A1(net6419),
    .S(_08345_),
    .X(_02437_));
 sg13g2_mux2_1 _27067_ (.A0(net4240),
    .A1(net6389),
    .S(_08345_),
    .X(_02438_));
 sg13g2_mux2_1 _27068_ (.A0(net3867),
    .A1(net6361),
    .S(_08345_),
    .X(_02439_));
 sg13g2_mux2_1 _27069_ (.A0(net3998),
    .A1(net6332),
    .S(_08345_),
    .X(_02440_));
 sg13g2_mux2_1 _27070_ (.A0(net3632),
    .A1(net6302),
    .S(_08345_),
    .X(_02441_));
 sg13g2_nand2_2 _27071_ (.Y(_08346_),
    .A(_08255_),
    .B(_08297_));
 sg13g2_mux2_1 _27072_ (.A0(net6475),
    .A1(net6603),
    .S(_08346_),
    .X(_02442_));
 sg13g2_mux2_1 _27073_ (.A0(net6449),
    .A1(net4528),
    .S(_08346_),
    .X(_02443_));
 sg13g2_mux2_1 _27074_ (.A0(net6420),
    .A1(net6893),
    .S(_08346_),
    .X(_02444_));
 sg13g2_mux2_1 _27075_ (.A0(net6390),
    .A1(net4585),
    .S(_08346_),
    .X(_02445_));
 sg13g2_mux2_1 _27076_ (.A0(net6361),
    .A1(net4812),
    .S(_08346_),
    .X(_02446_));
 sg13g2_mux2_1 _27077_ (.A0(net6331),
    .A1(net4785),
    .S(_08346_),
    .X(_02447_));
 sg13g2_mux2_1 _27078_ (.A0(net6303),
    .A1(net4491),
    .S(_08346_),
    .X(_02448_));
 sg13g2_nand2_2 _27079_ (.Y(_08347_),
    .A(net6028),
    .B(net5950));
 sg13g2_mux2_1 _27080_ (.A0(net6456),
    .A1(net4687),
    .S(_08347_),
    .X(_02449_));
 sg13g2_mux2_1 _27081_ (.A0(net6426),
    .A1(net4489),
    .S(_08347_),
    .X(_02450_));
 sg13g2_mux2_1 _27082_ (.A0(net6397),
    .A1(net4958),
    .S(_08347_),
    .X(_02451_));
 sg13g2_mux2_1 _27083_ (.A0(net6368),
    .A1(net6948),
    .S(_08347_),
    .X(_02452_));
 sg13g2_mux2_1 _27084_ (.A0(net6336),
    .A1(net4904),
    .S(_08347_),
    .X(_02453_));
 sg13g2_mux2_1 _27085_ (.A0(net6310),
    .A1(net4949),
    .S(_08347_),
    .X(_02454_));
 sg13g2_mux2_1 _27086_ (.A0(net6279),
    .A1(net7067),
    .S(_08347_),
    .X(_02455_));
 sg13g2_nor2_2 _27087_ (.A(net5959),
    .B(_08275_),
    .Y(_08348_));
 sg13g2_mux2_1 _27088_ (.A0(net3822),
    .A1(net6475),
    .S(_08348_),
    .X(_02456_));
 sg13g2_mux2_1 _27089_ (.A0(net3609),
    .A1(net6449),
    .S(_08348_),
    .X(_02457_));
 sg13g2_mux2_1 _27090_ (.A0(net3755),
    .A1(net6420),
    .S(_08348_),
    .X(_02458_));
 sg13g2_mux2_1 _27091_ (.A0(net4077),
    .A1(net6390),
    .S(_08348_),
    .X(_02459_));
 sg13g2_mux2_1 _27092_ (.A0(net3913),
    .A1(net6361),
    .S(_08348_),
    .X(_02460_));
 sg13g2_mux2_1 _27093_ (.A0(net4232),
    .A1(net6331),
    .S(_08348_),
    .X(_02461_));
 sg13g2_mux2_1 _27094_ (.A0(net4043),
    .A1(net6303),
    .S(_08348_),
    .X(_02462_));
 sg13g2_nor2_2 _27095_ (.A(_08246_),
    .B(net5959),
    .Y(_08349_));
 sg13g2_mux2_1 _27096_ (.A0(net4369),
    .A1(net6475),
    .S(_08349_),
    .X(_02463_));
 sg13g2_mux2_1 _27097_ (.A0(net3443),
    .A1(net6449),
    .S(_08349_),
    .X(_02464_));
 sg13g2_mux2_1 _27098_ (.A0(net3661),
    .A1(net6419),
    .S(_08349_),
    .X(_02465_));
 sg13g2_mux2_1 _27099_ (.A0(net4157),
    .A1(net6390),
    .S(_08349_),
    .X(_02466_));
 sg13g2_mux2_1 _27100_ (.A0(net4206),
    .A1(net6361),
    .S(_08349_),
    .X(_02467_));
 sg13g2_mux2_1 _27101_ (.A0(net3519),
    .A1(net6331),
    .S(_08349_),
    .X(_02468_));
 sg13g2_mux2_1 _27102_ (.A0(net4231),
    .A1(net6303),
    .S(_08349_),
    .X(_02469_));
 sg13g2_nor2_2 _27103_ (.A(_08256_),
    .B(_08279_),
    .Y(_08350_));
 sg13g2_mux2_1 _27104_ (.A0(net4008),
    .A1(net6475),
    .S(_08350_),
    .X(_02470_));
 sg13g2_mux2_1 _27105_ (.A0(net3837),
    .A1(net6446),
    .S(_08350_),
    .X(_02471_));
 sg13g2_mux2_1 _27106_ (.A0(net3339),
    .A1(net6419),
    .S(_08350_),
    .X(_02472_));
 sg13g2_mux2_1 _27107_ (.A0(net3594),
    .A1(net6389),
    .S(_08350_),
    .X(_02473_));
 sg13g2_mux2_1 _27108_ (.A0(net3697),
    .A1(net6361),
    .S(_08350_),
    .X(_02474_));
 sg13g2_mux2_1 _27109_ (.A0(net3953),
    .A1(net6331),
    .S(_08350_),
    .X(_02475_));
 sg13g2_mux2_1 _27110_ (.A0(net3698),
    .A1(net6301),
    .S(_08350_),
    .X(_02476_));
 sg13g2_nor2_2 _27111_ (.A(net5965),
    .B(_08256_),
    .Y(_08351_));
 sg13g2_mux2_1 _27112_ (.A0(net3700),
    .A1(net6475),
    .S(_08351_),
    .X(_02477_));
 sg13g2_mux2_1 _27113_ (.A0(net4055),
    .A1(net6450),
    .S(_08351_),
    .X(_02478_));
 sg13g2_mux2_1 _27114_ (.A0(net3928),
    .A1(net6419),
    .S(_08351_),
    .X(_02479_));
 sg13g2_mux2_1 _27115_ (.A0(net3633),
    .A1(net6389),
    .S(_08351_),
    .X(_02480_));
 sg13g2_mux2_1 _27116_ (.A0(net3690),
    .A1(net6361),
    .S(_08351_),
    .X(_02481_));
 sg13g2_mux2_1 _27117_ (.A0(net3968),
    .A1(net6331),
    .S(_08351_),
    .X(_02482_));
 sg13g2_mux2_1 _27118_ (.A0(net4011),
    .A1(net6301),
    .S(_08351_),
    .X(_02483_));
 sg13g2_nor2_2 _27119_ (.A(net5959),
    .B(net5952),
    .Y(_08352_));
 sg13g2_mux2_1 _27120_ (.A0(net4051),
    .A1(net6475),
    .S(_08352_),
    .X(_02484_));
 sg13g2_mux2_1 _27121_ (.A0(net3764),
    .A1(net6446),
    .S(_08352_),
    .X(_02485_));
 sg13g2_mux2_1 _27122_ (.A0(net3670),
    .A1(net6419),
    .S(_08352_),
    .X(_02486_));
 sg13g2_mux2_1 _27123_ (.A0(net3506),
    .A1(net6389),
    .S(_08352_),
    .X(_02487_));
 sg13g2_mux2_1 _27124_ (.A0(net4074),
    .A1(net6363),
    .S(_08352_),
    .X(_02488_));
 sg13g2_mux2_1 _27125_ (.A0(net4092),
    .A1(net6331),
    .S(_08352_),
    .X(_02489_));
 sg13g2_mux2_1 _27126_ (.A0(net3470),
    .A1(net6301),
    .S(_08352_),
    .X(_02490_));
 sg13g2_nor2_2 _27127_ (.A(net6030),
    .B(net5959),
    .Y(_08353_));
 sg13g2_mux2_1 _27128_ (.A0(net3729),
    .A1(net6475),
    .S(_08353_),
    .X(_02491_));
 sg13g2_mux2_1 _27129_ (.A0(net4201),
    .A1(net6450),
    .S(_08353_),
    .X(_02492_));
 sg13g2_mux2_1 _27130_ (.A0(net3962),
    .A1(net6419),
    .S(_08353_),
    .X(_02493_));
 sg13g2_mux2_1 _27131_ (.A0(net4132),
    .A1(net6389),
    .S(_08353_),
    .X(_02494_));
 sg13g2_mux2_1 _27132_ (.A0(net4047),
    .A1(net6361),
    .S(_08353_),
    .X(_02495_));
 sg13g2_mux2_1 _27133_ (.A0(net4416),
    .A1(net6331),
    .S(_08353_),
    .X(_02496_));
 sg13g2_mux2_1 _27134_ (.A0(net3749),
    .A1(net6301),
    .S(_08353_),
    .X(_02497_));
 sg13g2_nand2_2 _27135_ (.Y(_08354_),
    .A(net5969),
    .B(_08258_));
 sg13g2_mux2_1 _27136_ (.A0(net6470),
    .A1(net6773),
    .S(_08354_),
    .X(_02498_));
 sg13g2_mux2_1 _27137_ (.A0(net6446),
    .A1(net4935),
    .S(_08354_),
    .X(_02499_));
 sg13g2_mux2_1 _27138_ (.A0(net6417),
    .A1(net6961),
    .S(_08354_),
    .X(_02500_));
 sg13g2_mux2_1 _27139_ (.A0(net6388),
    .A1(net6918),
    .S(_08354_),
    .X(_02501_));
 sg13g2_mux2_1 _27140_ (.A0(net6359),
    .A1(net6755),
    .S(_08354_),
    .X(_02502_));
 sg13g2_mux2_1 _27141_ (.A0(net6329),
    .A1(net7046),
    .S(_08354_),
    .X(_02503_));
 sg13g2_mux2_1 _27142_ (.A0(net6299),
    .A1(net6929),
    .S(_08354_),
    .X(_02504_));
 sg13g2_nand2_2 _27143_ (.Y(_08355_),
    .A(net5962),
    .B(_08258_));
 sg13g2_mux2_1 _27144_ (.A0(net6477),
    .A1(net6789),
    .S(_08355_),
    .X(_02505_));
 sg13g2_mux2_1 _27145_ (.A0(net6446),
    .A1(net4767),
    .S(_08355_),
    .X(_02506_));
 sg13g2_mux2_1 _27146_ (.A0(net6417),
    .A1(net4773),
    .S(_08355_),
    .X(_02507_));
 sg13g2_mux2_1 _27147_ (.A0(net6388),
    .A1(net6713),
    .S(_08355_),
    .X(_02508_));
 sg13g2_mux2_1 _27148_ (.A0(net6359),
    .A1(net4672),
    .S(_08355_),
    .X(_02509_));
 sg13g2_mux2_1 _27149_ (.A0(net6329),
    .A1(net4608),
    .S(_08355_),
    .X(_02510_));
 sg13g2_mux2_1 _27150_ (.A0(net6299),
    .A1(net4547),
    .S(_08355_),
    .X(_02511_));
 sg13g2_nand2_2 _27151_ (.Y(_08356_),
    .A(_08258_),
    .B(net5953));
 sg13g2_mux2_1 _27152_ (.A0(net6470),
    .A1(net6737),
    .S(_08356_),
    .X(_02512_));
 sg13g2_mux2_1 _27153_ (.A0(net6446),
    .A1(net6847),
    .S(_08356_),
    .X(_02513_));
 sg13g2_mux2_1 _27154_ (.A0(net6417),
    .A1(net4836),
    .S(_08356_),
    .X(_02514_));
 sg13g2_mux2_1 _27155_ (.A0(net6388),
    .A1(net4766),
    .S(_08356_),
    .X(_02515_));
 sg13g2_mux2_1 _27156_ (.A0(net6360),
    .A1(net6935),
    .S(_08356_),
    .X(_02516_));
 sg13g2_mux2_1 _27157_ (.A0(net6329),
    .A1(net4760),
    .S(_08356_),
    .X(_02517_));
 sg13g2_mux2_1 _27158_ (.A0(net6299),
    .A1(net6746),
    .S(_08356_),
    .X(_02518_));
 sg13g2_nand2_2 _27159_ (.Y(_08357_),
    .A(net6028),
    .B(net5969));
 sg13g2_mux2_1 _27160_ (.A0(net6456),
    .A1(net4658),
    .S(_08357_),
    .X(_02519_));
 sg13g2_mux2_1 _27161_ (.A0(net6426),
    .A1(net6629),
    .S(_08357_),
    .X(_02520_));
 sg13g2_mux2_1 _27162_ (.A0(net6397),
    .A1(net4809),
    .S(_08357_),
    .X(_02521_));
 sg13g2_mux2_1 _27163_ (.A0(net6368),
    .A1(net4548),
    .S(_08357_),
    .X(_02522_));
 sg13g2_mux2_1 _27164_ (.A0(net6341),
    .A1(net6891),
    .S(_08357_),
    .X(_02523_));
 sg13g2_mux2_1 _27165_ (.A0(net6309),
    .A1(net4882),
    .S(_08357_),
    .X(_02524_));
 sg13g2_mux2_1 _27166_ (.A0(net6279),
    .A1(net4752),
    .S(_08357_),
    .X(_02525_));
 sg13g2_nand2_2 _27167_ (.Y(_08358_),
    .A(_08258_),
    .B(net5951));
 sg13g2_mux2_1 _27168_ (.A0(net6477),
    .A1(net4724),
    .S(_08358_),
    .X(_02526_));
 sg13g2_mux2_1 _27169_ (.A0(net6447),
    .A1(net6605),
    .S(_08358_),
    .X(_02527_));
 sg13g2_mux2_1 _27170_ (.A0(net6417),
    .A1(net4664),
    .S(_08358_),
    .X(_02528_));
 sg13g2_mux2_1 _27171_ (.A0(net6387),
    .A1(net6590),
    .S(_08358_),
    .X(_02529_));
 sg13g2_mux2_1 _27172_ (.A0(net6359),
    .A1(net6620),
    .S(_08358_),
    .X(_02530_));
 sg13g2_mux2_1 _27173_ (.A0(net6327),
    .A1(net4365),
    .S(_08358_),
    .X(_02531_));
 sg13g2_mux2_1 _27174_ (.A0(net6299),
    .A1(net4865),
    .S(_08358_),
    .X(_02532_));
 sg13g2_nor2_2 _27175_ (.A(_08252_),
    .B(_08259_),
    .Y(_08359_));
 sg13g2_mux2_1 _27176_ (.A0(net4167),
    .A1(net6477),
    .S(_08359_),
    .X(_02533_));
 sg13g2_mux2_1 _27177_ (.A0(net3736),
    .A1(net6447),
    .S(_08359_),
    .X(_02534_));
 sg13g2_mux2_1 _27178_ (.A0(net4320),
    .A1(net6417),
    .S(_08359_),
    .X(_02535_));
 sg13g2_mux2_1 _27179_ (.A0(net4140),
    .A1(net6387),
    .S(_08359_),
    .X(_02536_));
 sg13g2_mux2_1 _27180_ (.A0(net4143),
    .A1(net6359),
    .S(_08359_),
    .X(_02537_));
 sg13g2_mux2_1 _27181_ (.A0(net3772),
    .A1(net6327),
    .S(_08359_),
    .X(_02538_));
 sg13g2_mux2_1 _27182_ (.A0(net3817),
    .A1(net6299),
    .S(_08359_),
    .X(_02539_));
 sg13g2_nor2_2 _27183_ (.A(net5958),
    .B(_08294_),
    .Y(_08360_));
 sg13g2_mux2_1 _27184_ (.A0(net4148),
    .A1(net6470),
    .S(_08360_),
    .X(_02540_));
 sg13g2_mux2_1 _27185_ (.A0(net3927),
    .A1(net6447),
    .S(_08360_),
    .X(_02541_));
 sg13g2_mux2_1 _27186_ (.A0(net4149),
    .A1(net6417),
    .S(_08360_),
    .X(_02542_));
 sg13g2_mux2_1 _27187_ (.A0(net4202),
    .A1(net6387),
    .S(_08360_),
    .X(_02543_));
 sg13g2_mux2_1 _27188_ (.A0(net3511),
    .A1(net6359),
    .S(_08360_),
    .X(_02544_));
 sg13g2_mux2_1 _27189_ (.A0(net3161),
    .A1(net6329),
    .S(_08360_),
    .X(_02545_));
 sg13g2_mux2_1 _27190_ (.A0(net3893),
    .A1(net6299),
    .S(_08360_),
    .X(_02546_));
 sg13g2_nor2_2 _27191_ (.A(_08237_),
    .B(net5958),
    .Y(_08361_));
 sg13g2_mux2_1 _27192_ (.A0(net4057),
    .A1(net6470),
    .S(_08361_),
    .X(_02547_));
 sg13g2_mux2_1 _27193_ (.A0(net3898),
    .A1(net6447),
    .S(_08361_),
    .X(_02548_));
 sg13g2_mux2_1 _27194_ (.A0(net3681),
    .A1(net6417),
    .S(_08361_),
    .X(_02549_));
 sg13g2_mux2_1 _27195_ (.A0(net3668),
    .A1(net6387),
    .S(_08361_),
    .X(_02550_));
 sg13g2_mux2_1 _27196_ (.A0(net3517),
    .A1(net6359),
    .S(_08361_),
    .X(_02551_));
 sg13g2_mux2_1 _27197_ (.A0(net4144),
    .A1(net6329),
    .S(_08361_),
    .X(_02552_));
 sg13g2_mux2_1 _27198_ (.A0(net3849),
    .A1(net6299),
    .S(_08361_),
    .X(_02553_));
 sg13g2_nand2_2 _27199_ (.Y(_08362_),
    .A(_08258_),
    .B(net5950));
 sg13g2_mux2_1 _27200_ (.A0(net6473),
    .A1(net6813),
    .S(_08362_),
    .X(_02554_));
 sg13g2_mux2_1 _27201_ (.A0(net6444),
    .A1(net6583),
    .S(_08362_),
    .X(_02555_));
 sg13g2_mux2_1 _27202_ (.A0(net6415),
    .A1(net6594),
    .S(_08362_),
    .X(_02556_));
 sg13g2_mux2_1 _27203_ (.A0(net6386),
    .A1(net4626),
    .S(_08362_),
    .X(_02557_));
 sg13g2_mux2_1 _27204_ (.A0(net6357),
    .A1(net6876),
    .S(_08362_),
    .X(_02558_));
 sg13g2_mux2_1 _27205_ (.A0(net6327),
    .A1(net7100),
    .S(_08362_),
    .X(_02559_));
 sg13g2_mux2_1 _27206_ (.A0(net6298),
    .A1(net6954),
    .S(_08362_),
    .X(_02560_));
 sg13g2_nor2_2 _27207_ (.A(_03132_),
    .B(net5958),
    .Y(_08363_));
 sg13g2_mux2_1 _27208_ (.A0(net3417),
    .A1(net6473),
    .S(_08363_),
    .X(_02561_));
 sg13g2_mux2_1 _27209_ (.A0(net3678),
    .A1(net6451),
    .S(_08363_),
    .X(_02562_));
 sg13g2_mux2_1 _27210_ (.A0(net3429),
    .A1(net6415),
    .S(_08363_),
    .X(_02563_));
 sg13g2_mux2_1 _27211_ (.A0(net4025),
    .A1(net6386),
    .S(_08363_),
    .X(_02564_));
 sg13g2_mux2_1 _27212_ (.A0(net3539),
    .A1(net6357),
    .S(_08363_),
    .X(_02565_));
 sg13g2_mux2_1 _27213_ (.A0(net3824),
    .A1(net6326),
    .S(_08363_),
    .X(_02566_));
 sg13g2_mux2_1 _27214_ (.A0(net3548),
    .A1(net6298),
    .S(_08363_),
    .X(_02567_));
 sg13g2_nor2_2 _27215_ (.A(net5958),
    .B(_08275_),
    .Y(_08364_));
 sg13g2_mux2_1 _27216_ (.A0(net3684),
    .A1(net6473),
    .S(_08364_),
    .X(_02568_));
 sg13g2_mux2_1 _27217_ (.A0(net3498),
    .A1(net6445),
    .S(_08364_),
    .X(_02569_));
 sg13g2_mux2_1 _27218_ (.A0(net4053),
    .A1(net6415),
    .S(_08364_),
    .X(_02570_));
 sg13g2_mux2_1 _27219_ (.A0(net3997),
    .A1(net6386),
    .S(_08364_),
    .X(_02571_));
 sg13g2_mux2_1 _27220_ (.A0(net3839),
    .A1(net6357),
    .S(_08364_),
    .X(_02572_));
 sg13g2_mux2_1 _27221_ (.A0(net4099),
    .A1(net6328),
    .S(_08364_),
    .X(_02573_));
 sg13g2_mux2_1 _27222_ (.A0(net3673),
    .A1(net6298),
    .S(_08364_),
    .X(_02574_));
 sg13g2_nor2_2 _27223_ (.A(_08246_),
    .B(net5958),
    .Y(_08365_));
 sg13g2_mux2_1 _27224_ (.A0(net4026),
    .A1(net6473),
    .S(_08365_),
    .X(_02575_));
 sg13g2_mux2_1 _27225_ (.A0(net3502),
    .A1(net6445),
    .S(_08365_),
    .X(_02576_));
 sg13g2_mux2_1 _27226_ (.A0(net3701),
    .A1(net6415),
    .S(_08365_),
    .X(_02577_));
 sg13g2_mux2_1 _27227_ (.A0(net3579),
    .A1(net6386),
    .S(_08365_),
    .X(_02578_));
 sg13g2_mux2_1 _27228_ (.A0(net3969),
    .A1(net6357),
    .S(_08365_),
    .X(_02579_));
 sg13g2_mux2_1 _27229_ (.A0(net4042),
    .A1(net6326),
    .S(_08365_),
    .X(_02580_));
 sg13g2_mux2_1 _27230_ (.A0(net3865),
    .A1(net6298),
    .S(_08365_),
    .X(_02581_));
 sg13g2_nor2_2 _27231_ (.A(net5958),
    .B(_08279_),
    .Y(_08366_));
 sg13g2_mux2_1 _27232_ (.A0(net3550),
    .A1(net6473),
    .S(_08366_),
    .X(_02582_));
 sg13g2_mux2_1 _27233_ (.A0(net3679),
    .A1(net6447),
    .S(_08366_),
    .X(_02583_));
 sg13g2_mux2_1 _27234_ (.A0(net3907),
    .A1(net6421),
    .S(_08366_),
    .X(_02584_));
 sg13g2_mux2_1 _27235_ (.A0(net3659),
    .A1(net6386),
    .S(_08366_),
    .X(_02585_));
 sg13g2_mux2_1 _27236_ (.A0(net3832),
    .A1(net6362),
    .S(_08366_),
    .X(_02586_));
 sg13g2_mux2_1 _27237_ (.A0(net3515),
    .A1(net6329),
    .S(_08366_),
    .X(_02587_));
 sg13g2_mux2_1 _27238_ (.A0(net3789),
    .A1(net6301),
    .S(_08366_),
    .X(_02588_));
 sg13g2_nand2_2 _27239_ (.Y(_08367_),
    .A(net6027),
    .B(_08274_));
 sg13g2_mux2_1 _27240_ (.A0(net6456),
    .A1(net4854),
    .S(_08367_),
    .X(_02589_));
 sg13g2_mux2_1 _27241_ (.A0(net6426),
    .A1(net4891),
    .S(_08367_),
    .X(_02590_));
 sg13g2_mux2_1 _27242_ (.A0(net6397),
    .A1(net4864),
    .S(_08367_),
    .X(_02591_));
 sg13g2_mux2_1 _27243_ (.A0(net6368),
    .A1(net4611),
    .S(_08367_),
    .X(_02592_));
 sg13g2_mux2_1 _27244_ (.A0(net6336),
    .A1(net6878),
    .S(_08367_),
    .X(_02593_));
 sg13g2_mux2_1 _27245_ (.A0(net6310),
    .A1(net6778),
    .S(_08367_),
    .X(_02594_));
 sg13g2_mux2_1 _27246_ (.A0(net6279),
    .A1(net6837),
    .S(_08367_),
    .X(_02595_));
 sg13g2_nor2_2 _27247_ (.A(net5958),
    .B(net5952),
    .Y(_08368_));
 sg13g2_mux2_1 _27248_ (.A0(net3751),
    .A1(net6472),
    .S(_08368_),
    .X(_02596_));
 sg13g2_mux2_1 _27249_ (.A0(net4127),
    .A1(net6447),
    .S(_08368_),
    .X(_02597_));
 sg13g2_mux2_1 _27250_ (.A0(net4125),
    .A1(net6421),
    .S(_08368_),
    .X(_02598_));
 sg13g2_mux2_1 _27251_ (.A0(net3591),
    .A1(net6386),
    .S(_08368_),
    .X(_02599_));
 sg13g2_mux2_1 _27252_ (.A0(net3504),
    .A1(net6362),
    .S(_08368_),
    .X(_02600_));
 sg13g2_mux2_1 _27253_ (.A0(net4363),
    .A1(net6332),
    .S(_08368_),
    .X(_02601_));
 sg13g2_mux2_1 _27254_ (.A0(net3479),
    .A1(net6301),
    .S(_08368_),
    .X(_02602_));
 sg13g2_nor2_2 _27255_ (.A(net6029),
    .B(net5958),
    .Y(_08369_));
 sg13g2_mux2_1 _27256_ (.A0(net4086),
    .A1(net6476),
    .S(_08369_),
    .X(_02603_));
 sg13g2_mux2_1 _27257_ (.A0(net3923),
    .A1(net6447),
    .S(_08369_),
    .X(_02604_));
 sg13g2_mux2_1 _27258_ (.A0(net3926),
    .A1(net6421),
    .S(_08369_),
    .X(_02605_));
 sg13g2_mux2_1 _27259_ (.A0(net3881),
    .A1(net6386),
    .S(_08369_),
    .X(_02606_));
 sg13g2_mux2_1 _27260_ (.A0(net3852),
    .A1(net6362),
    .S(_08369_),
    .X(_02607_));
 sg13g2_mux2_1 _27261_ (.A0(net3793),
    .A1(net6329),
    .S(_08369_),
    .X(_02608_));
 sg13g2_mux2_1 _27262_ (.A0(net3551),
    .A1(net6301),
    .S(_08369_),
    .X(_02609_));
 sg13g2_nand2_2 _27263_ (.Y(_08370_),
    .A(net5969),
    .B(_08262_));
 sg13g2_mux2_1 _27264_ (.A0(net6474),
    .A1(net4584),
    .S(_08370_),
    .X(_02610_));
 sg13g2_mux2_1 _27265_ (.A0(net6444),
    .A1(net6901),
    .S(_08370_),
    .X(_02611_));
 sg13g2_mux2_1 _27266_ (.A0(net6416),
    .A1(net4698),
    .S(_08370_),
    .X(_02612_));
 sg13g2_mux2_1 _27267_ (.A0(net6387),
    .A1(net4599),
    .S(_08370_),
    .X(_02613_));
 sg13g2_mux2_1 _27268_ (.A0(net6358),
    .A1(net6974),
    .S(_08370_),
    .X(_02614_));
 sg13g2_mux2_1 _27269_ (.A0(net6327),
    .A1(net6843),
    .S(_08370_),
    .X(_02615_));
 sg13g2_mux2_1 _27270_ (.A0(net6297),
    .A1(net7072),
    .S(_08370_),
    .X(_02616_));
 sg13g2_and2_2 _27271_ (.A(_08241_),
    .B(_08262_),
    .X(_08371_));
 sg13g2_mux2_1 _27272_ (.A0(net4020),
    .A1(net6474),
    .S(_08371_),
    .X(_02617_));
 sg13g2_mux2_1 _27273_ (.A0(net4307),
    .A1(net6444),
    .S(_08371_),
    .X(_02618_));
 sg13g2_mux2_1 _27274_ (.A0(net3974),
    .A1(net6416),
    .S(_08371_),
    .X(_02619_));
 sg13g2_mux2_1 _27275_ (.A0(net4016),
    .A1(net6387),
    .S(_08371_),
    .X(_02620_));
 sg13g2_mux2_1 _27276_ (.A0(net3686),
    .A1(net6358),
    .S(_08371_),
    .X(_02621_));
 sg13g2_mux2_1 _27277_ (.A0(net3901),
    .A1(net6327),
    .S(_08371_),
    .X(_02622_));
 sg13g2_mux2_1 _27278_ (.A0(net4222),
    .A1(net6297),
    .S(_08371_),
    .X(_02623_));
 sg13g2_and2_2 _27279_ (.A(_08262_),
    .B(_08281_),
    .X(_08372_));
 sg13g2_mux2_1 _27280_ (.A0(net4183),
    .A1(net6474),
    .S(_08372_),
    .X(_02624_));
 sg13g2_mux2_1 _27281_ (.A0(net3874),
    .A1(net6444),
    .S(_08372_),
    .X(_02625_));
 sg13g2_mux2_1 _27282_ (.A0(net3763),
    .A1(net6414),
    .S(_08372_),
    .X(_02626_));
 sg13g2_mux2_1 _27283_ (.A0(net4093),
    .A1(net6387),
    .S(_08372_),
    .X(_02627_));
 sg13g2_mux2_1 _27284_ (.A0(net4182),
    .A1(net6358),
    .S(_08372_),
    .X(_02628_));
 sg13g2_mux2_1 _27285_ (.A0(net3472),
    .A1(net6327),
    .S(_08372_),
    .X(_02629_));
 sg13g2_mux2_1 _27286_ (.A0(net4239),
    .A1(net6297),
    .S(_08372_),
    .X(_02630_));
 sg13g2_and2_2 _27287_ (.A(net5968),
    .B(_08262_),
    .X(_08373_));
 sg13g2_mux2_1 _27288_ (.A0(net3889),
    .A1(net6474),
    .S(_08373_),
    .X(_02631_));
 sg13g2_mux2_1 _27289_ (.A0(net3995),
    .A1(net6444),
    .S(_08373_),
    .X(_02632_));
 sg13g2_mux2_1 _27290_ (.A0(net3808),
    .A1(net6416),
    .S(_08373_),
    .X(_02633_));
 sg13g2_mux2_1 _27291_ (.A0(net3581),
    .A1(net6387),
    .S(_08373_),
    .X(_02634_));
 sg13g2_mux2_1 _27292_ (.A0(net4205),
    .A1(net6358),
    .S(_08373_),
    .X(_02635_));
 sg13g2_mux2_1 _27293_ (.A0(net4159),
    .A1(net6327),
    .S(_08373_),
    .X(_02636_));
 sg13g2_mux2_1 _27294_ (.A0(net3863),
    .A1(net6297),
    .S(_08373_),
    .X(_02637_));
 sg13g2_nand2_2 _27295_ (.Y(_08374_),
    .A(_08262_),
    .B(_08290_));
 sg13g2_mux2_1 _27296_ (.A0(net6472),
    .A1(net4712),
    .S(_08374_),
    .X(_02638_));
 sg13g2_mux2_1 _27297_ (.A0(net6443),
    .A1(net7199),
    .S(_08374_),
    .X(_02639_));
 sg13g2_mux2_1 _27298_ (.A0(net6414),
    .A1(net6648),
    .S(_08374_),
    .X(_02640_));
 sg13g2_mux2_1 _27299_ (.A0(net6385),
    .A1(net6604),
    .S(_08374_),
    .X(_02641_));
 sg13g2_mux2_1 _27300_ (.A0(net6356),
    .A1(net4730),
    .S(_08374_),
    .X(_02642_));
 sg13g2_mux2_1 _27301_ (.A0(net6326),
    .A1(net4686),
    .S(_08374_),
    .X(_02643_));
 sg13g2_mux2_1 _27302_ (.A0(net6296),
    .A1(net6660),
    .S(_08374_),
    .X(_02644_));
 sg13g2_nor2_2 _27303_ (.A(_08252_),
    .B(_08263_),
    .Y(_08375_));
 sg13g2_mux2_1 _27304_ (.A0(net4428),
    .A1(net6472),
    .S(_08375_),
    .X(_02645_));
 sg13g2_mux2_1 _27305_ (.A0(net3740),
    .A1(net6443),
    .S(_08375_),
    .X(_02646_));
 sg13g2_mux2_1 _27306_ (.A0(net3458),
    .A1(net6414),
    .S(_08375_),
    .X(_02647_));
 sg13g2_mux2_1 _27307_ (.A0(net3478),
    .A1(net6385),
    .S(_08375_),
    .X(_02648_));
 sg13g2_mux2_1 _27308_ (.A0(net3765),
    .A1(net6356),
    .S(_08375_),
    .X(_02649_));
 sg13g2_mux2_1 _27309_ (.A0(net4355),
    .A1(net6326),
    .S(_08375_),
    .X(_02650_));
 sg13g2_mux2_1 _27310_ (.A0(net4007),
    .A1(net6296),
    .S(_08375_),
    .X(_02651_));
 sg13g2_nor2_2 _27311_ (.A(net5957),
    .B(_08294_),
    .Y(_08376_));
 sg13g2_mux2_1 _27312_ (.A0(net4221),
    .A1(net6472),
    .S(_08376_),
    .X(_02652_));
 sg13g2_mux2_1 _27313_ (.A0(net3760),
    .A1(net6443),
    .S(_08376_),
    .X(_02653_));
 sg13g2_mux2_1 _27314_ (.A0(net4130),
    .A1(net6415),
    .S(_08376_),
    .X(_02654_));
 sg13g2_mux2_1 _27315_ (.A0(net4100),
    .A1(net6385),
    .S(_08376_),
    .X(_02655_));
 sg13g2_mux2_1 _27316_ (.A0(net4054),
    .A1(net6356),
    .S(_08376_),
    .X(_02656_));
 sg13g2_mux2_1 _27317_ (.A0(net4463),
    .A1(net6326),
    .S(_08376_),
    .X(_02657_));
 sg13g2_mux2_1 _27318_ (.A0(net4022),
    .A1(net6296),
    .S(_08376_),
    .X(_02658_));
 sg13g2_nand2_2 _27319_ (.Y(_08377_),
    .A(net6027),
    .B(_08245_));
 sg13g2_mux2_1 _27320_ (.A0(net6456),
    .A1(net4754),
    .S(_08377_),
    .X(_02659_));
 sg13g2_mux2_1 _27321_ (.A0(net6426),
    .A1(net4653),
    .S(_08377_),
    .X(_02660_));
 sg13g2_mux2_1 _27322_ (.A0(net6397),
    .A1(net6705),
    .S(_08377_),
    .X(_02661_));
 sg13g2_mux2_1 _27323_ (.A0(net6368),
    .A1(net6636),
    .S(_08377_),
    .X(_02662_));
 sg13g2_mux2_1 _27324_ (.A0(net6341),
    .A1(net7103),
    .S(_08377_),
    .X(_02663_));
 sg13g2_mux2_1 _27325_ (.A0(net6310),
    .A1(net7074),
    .S(_08377_),
    .X(_02664_));
 sg13g2_mux2_1 _27326_ (.A0(net6279),
    .A1(net6956),
    .S(_08377_),
    .X(_02665_));
 sg13g2_nand2_2 _27327_ (.Y(_08378_),
    .A(_08262_),
    .B(net5950));
 sg13g2_mux2_1 _27328_ (.A0(net6474),
    .A1(net4789),
    .S(_08378_),
    .X(_02666_));
 sg13g2_mux2_1 _27329_ (.A0(net6445),
    .A1(net6788),
    .S(_08378_),
    .X(_02667_));
 sg13g2_mux2_1 _27330_ (.A0(net6415),
    .A1(net6826),
    .S(_08378_),
    .X(_02668_));
 sg13g2_mux2_1 _27331_ (.A0(net6385),
    .A1(net4617),
    .S(_08378_),
    .X(_02669_));
 sg13g2_mux2_1 _27332_ (.A0(net6356),
    .A1(net4508),
    .S(_08378_),
    .X(_02670_));
 sg13g2_mux2_1 _27333_ (.A0(net6326),
    .A1(net6731),
    .S(_08378_),
    .X(_02671_));
 sg13g2_mux2_1 _27334_ (.A0(net6304),
    .A1(net6698),
    .S(_08378_),
    .X(_02672_));
 sg13g2_nor2_2 _27335_ (.A(_03132_),
    .B(net5957),
    .Y(_08379_));
 sg13g2_mux2_1 _27336_ (.A0(net3563),
    .A1(net6472),
    .S(_08379_),
    .X(_02673_));
 sg13g2_mux2_1 _27337_ (.A0(net3818),
    .A1(net6445),
    .S(_08379_),
    .X(_02674_));
 sg13g2_mux2_1 _27338_ (.A0(net4124),
    .A1(net6416),
    .S(_08379_),
    .X(_02675_));
 sg13g2_mux2_1 _27339_ (.A0(net3846),
    .A1(net6385),
    .S(_08379_),
    .X(_02676_));
 sg13g2_mux2_1 _27340_ (.A0(net4046),
    .A1(net6356),
    .S(_08379_),
    .X(_02677_));
 sg13g2_mux2_1 _27341_ (.A0(net3890),
    .A1(net6326),
    .S(_08379_),
    .X(_02678_));
 sg13g2_mux2_1 _27342_ (.A0(net3631),
    .A1(net6304),
    .S(_08379_),
    .X(_02679_));
 sg13g2_nor2_2 _27343_ (.A(net5957),
    .B(_08275_),
    .Y(_08380_));
 sg13g2_mux2_1 _27344_ (.A0(net3748),
    .A1(net6472),
    .S(_08380_),
    .X(_02680_));
 sg13g2_mux2_1 _27345_ (.A0(net3721),
    .A1(net6445),
    .S(_08380_),
    .X(_02681_));
 sg13g2_mux2_1 _27346_ (.A0(net3509),
    .A1(net6415),
    .S(_08380_),
    .X(_02682_));
 sg13g2_mux2_1 _27347_ (.A0(net3590),
    .A1(net6385),
    .S(_08380_),
    .X(_02683_));
 sg13g2_mux2_1 _27348_ (.A0(net4344),
    .A1(net6356),
    .S(_08380_),
    .X(_02684_));
 sg13g2_mux2_1 _27349_ (.A0(net4286),
    .A1(net6328),
    .S(_08380_),
    .X(_02685_));
 sg13g2_mux2_1 _27350_ (.A0(net4045),
    .A1(net6298),
    .S(_08380_),
    .X(_02686_));
 sg13g2_nor2_2 _27351_ (.A(_08246_),
    .B(net5957),
    .Y(_08381_));
 sg13g2_mux2_1 _27352_ (.A0(net3801),
    .A1(net6472),
    .S(_08381_),
    .X(_02687_));
 sg13g2_mux2_1 _27353_ (.A0(net3960),
    .A1(net6445),
    .S(_08381_),
    .X(_02688_));
 sg13g2_mux2_1 _27354_ (.A0(net4028),
    .A1(net6415),
    .S(_08381_),
    .X(_02689_));
 sg13g2_mux2_1 _27355_ (.A0(net3785),
    .A1(net6385),
    .S(_08381_),
    .X(_02690_));
 sg13g2_mux2_1 _27356_ (.A0(net3541),
    .A1(net6356),
    .S(_08381_),
    .X(_02691_));
 sg13g2_mux2_1 _27357_ (.A0(net4269),
    .A1(net6328),
    .S(_08381_),
    .X(_02692_));
 sg13g2_mux2_1 _27358_ (.A0(net3780),
    .A1(net6298),
    .S(_08381_),
    .X(_02693_));
 sg13g2_nor2_2 _27359_ (.A(net5957),
    .B(_08279_),
    .Y(_08382_));
 sg13g2_mux2_1 _27360_ (.A0(net4080),
    .A1(net6466),
    .S(_08382_),
    .X(_02694_));
 sg13g2_mux2_1 _27361_ (.A0(net4017),
    .A1(net6435),
    .S(_08382_),
    .X(_02695_));
 sg13g2_mux2_1 _27362_ (.A0(net3774),
    .A1(net6411),
    .S(_08382_),
    .X(_02696_));
 sg13g2_mux2_1 _27363_ (.A0(net3587),
    .A1(net6383),
    .S(_08382_),
    .X(_02697_));
 sg13g2_mux2_1 _27364_ (.A0(net3694),
    .A1(net6349),
    .S(_08382_),
    .X(_02698_));
 sg13g2_mux2_1 _27365_ (.A0(net3987),
    .A1(net6321),
    .S(_08382_),
    .X(_02699_));
 sg13g2_mux2_1 _27366_ (.A0(net3977),
    .A1(net6293),
    .S(_08382_),
    .X(_02700_));
 sg13g2_nor2_2 _27367_ (.A(net5965),
    .B(net5957),
    .Y(_08383_));
 sg13g2_mux2_1 _27368_ (.A0(net3447),
    .A1(net6465),
    .S(_08383_),
    .X(_02701_));
 sg13g2_mux2_1 _27369_ (.A0(net3892),
    .A1(net6435),
    .S(_08383_),
    .X(_02702_));
 sg13g2_mux2_1 _27370_ (.A0(net3858),
    .A1(net6411),
    .S(_08383_),
    .X(_02703_));
 sg13g2_mux2_1 _27371_ (.A0(net3578),
    .A1(net6383),
    .S(_08383_),
    .X(_02704_));
 sg13g2_mux2_1 _27372_ (.A0(net4056),
    .A1(net6349),
    .S(_08383_),
    .X(_02705_));
 sg13g2_mux2_1 _27373_ (.A0(net3624),
    .A1(net6321),
    .S(_08383_),
    .X(_02706_));
 sg13g2_mux2_1 _27374_ (.A0(net3924),
    .A1(net6293),
    .S(_08383_),
    .X(_02707_));
 sg13g2_nor2_2 _27375_ (.A(net5957),
    .B(net5952),
    .Y(_08384_));
 sg13g2_mux2_1 _27376_ (.A0(net3936),
    .A1(net6465),
    .S(_08384_),
    .X(_02708_));
 sg13g2_mux2_1 _27377_ (.A0(net4179),
    .A1(net6435),
    .S(_08384_),
    .X(_02709_));
 sg13g2_mux2_1 _27378_ (.A0(net4241),
    .A1(net6411),
    .S(_08384_),
    .X(_02710_));
 sg13g2_mux2_1 _27379_ (.A0(net3815),
    .A1(net6379),
    .S(_08384_),
    .X(_02711_));
 sg13g2_mux2_1 _27380_ (.A0(net3707),
    .A1(net6349),
    .S(_08384_),
    .X(_02712_));
 sg13g2_mux2_1 _27381_ (.A0(net3756),
    .A1(net6321),
    .S(_08384_),
    .X(_02713_));
 sg13g2_mux2_1 _27382_ (.A0(net4118),
    .A1(net6293),
    .S(_08384_),
    .X(_02714_));
 sg13g2_nor2_2 _27383_ (.A(net6030),
    .B(net5957),
    .Y(_08385_));
 sg13g2_mux2_1 _27384_ (.A0(net4235),
    .A1(net6465),
    .S(_08385_),
    .X(_02715_));
 sg13g2_mux2_1 _27385_ (.A0(net3699),
    .A1(net6435),
    .S(_08385_),
    .X(_02716_));
 sg13g2_mux2_1 _27386_ (.A0(net3944),
    .A1(net6411),
    .S(_08385_),
    .X(_02717_));
 sg13g2_mux2_1 _27387_ (.A0(net3483),
    .A1(net6379),
    .S(_08385_),
    .X(_02718_));
 sg13g2_mux2_1 _27388_ (.A0(net4033),
    .A1(net6349),
    .S(_08385_),
    .X(_02719_));
 sg13g2_mux2_1 _27389_ (.A0(net4473),
    .A1(net6320),
    .S(_08385_),
    .X(_02720_));
 sg13g2_mux2_1 _27390_ (.A0(net3767),
    .A1(net6293),
    .S(_08385_),
    .X(_02721_));
 sg13g2_nand2_2 _27391_ (.Y(_08386_),
    .A(net5969),
    .B(net5956));
 sg13g2_mux2_1 _27392_ (.A0(net6457),
    .A1(net4844),
    .S(_08386_),
    .X(_02722_));
 sg13g2_mux2_1 _27393_ (.A0(net6427),
    .A1(net4603),
    .S(_08386_),
    .X(_02723_));
 sg13g2_mux2_1 _27394_ (.A0(net6394),
    .A1(net6650),
    .S(_08386_),
    .X(_02724_));
 sg13g2_mux2_1 _27395_ (.A0(net6367),
    .A1(net4503),
    .S(_08386_),
    .X(_02725_));
 sg13g2_mux2_1 _27396_ (.A0(net6337),
    .A1(net4588),
    .S(_08386_),
    .X(_02726_));
 sg13g2_mux2_1 _27397_ (.A0(net6313),
    .A1(net4631),
    .S(_08386_),
    .X(_02727_));
 sg13g2_mux2_1 _27398_ (.A0(net6282),
    .A1(net6587),
    .S(_08386_),
    .X(_02728_));
 sg13g2_nand2_2 _27399_ (.Y(_08387_),
    .A(net6027),
    .B(_08278_));
 sg13g2_mux2_1 _27400_ (.A0(net6454),
    .A1(net4901),
    .S(_08387_),
    .X(_02729_));
 sg13g2_mux2_1 _27401_ (.A0(net6425),
    .A1(net4886),
    .S(_08387_),
    .X(_02730_));
 sg13g2_mux2_1 _27402_ (.A0(net6396),
    .A1(net4654),
    .S(_08387_),
    .X(_02731_));
 sg13g2_mux2_1 _27403_ (.A0(net6365),
    .A1(net4691),
    .S(_08387_),
    .X(_02732_));
 sg13g2_mux2_1 _27404_ (.A0(net6335),
    .A1(net6621),
    .S(_08387_),
    .X(_02733_));
 sg13g2_mux2_1 _27405_ (.A0(net6306),
    .A1(net6832),
    .S(_08387_),
    .X(_02734_));
 sg13g2_mux2_1 _27406_ (.A0(net6277),
    .A1(net6645),
    .S(_08387_),
    .X(_02735_));
 sg13g2_nand2_2 _27407_ (.Y(_08388_),
    .A(net5956),
    .B(net5953));
 sg13g2_mux2_1 _27408_ (.A0(net6457),
    .A1(net6734),
    .S(_08388_),
    .X(_02736_));
 sg13g2_mux2_1 _27409_ (.A0(net6427),
    .A1(net6782),
    .S(_08388_),
    .X(_02737_));
 sg13g2_mux2_1 _27410_ (.A0(net6399),
    .A1(net4858),
    .S(_08388_),
    .X(_02738_));
 sg13g2_mux2_1 _27411_ (.A0(net6370),
    .A1(net6801),
    .S(_08388_),
    .X(_02739_));
 sg13g2_mux2_1 _27412_ (.A0(net6337),
    .A1(net4744),
    .S(_08388_),
    .X(_02740_));
 sg13g2_mux2_1 _27413_ (.A0(net6312),
    .A1(net6687),
    .S(_08388_),
    .X(_02741_));
 sg13g2_mux2_1 _27414_ (.A0(net6278),
    .A1(net7035),
    .S(_08388_),
    .X(_02742_));
 sg13g2_nand2_2 _27415_ (.Y(_08389_),
    .A(net5968),
    .B(net5956));
 sg13g2_mux2_1 _27416_ (.A0(net6457),
    .A1(net4840),
    .S(_08389_),
    .X(_02743_));
 sg13g2_mux2_1 _27417_ (.A0(net6427),
    .A1(net6647),
    .S(_08389_),
    .X(_02744_));
 sg13g2_mux2_1 _27418_ (.A0(net6399),
    .A1(net4613),
    .S(_08389_),
    .X(_02745_));
 sg13g2_mux2_1 _27419_ (.A0(net6370),
    .A1(net4747),
    .S(_08389_),
    .X(_02746_));
 sg13g2_mux2_1 _27420_ (.A0(net6337),
    .A1(net6880),
    .S(_08389_),
    .X(_02747_));
 sg13g2_mux2_1 _27421_ (.A0(net6312),
    .A1(net7142),
    .S(_08389_),
    .X(_02748_));
 sg13g2_mux2_1 _27422_ (.A0(net6278),
    .A1(net6995),
    .S(_08389_),
    .X(_02749_));
 sg13g2_nand2_2 _27423_ (.Y(_08390_),
    .A(net5955),
    .B(net5951));
 sg13g2_mux2_1 _27424_ (.A0(net6452),
    .A1(net6917),
    .S(_08390_),
    .X(_02750_));
 sg13g2_mux2_1 _27425_ (.A0(net6423),
    .A1(net6996),
    .S(_08390_),
    .X(_02751_));
 sg13g2_mux2_1 _27426_ (.A0(net6394),
    .A1(net6717),
    .S(_08390_),
    .X(_02752_));
 sg13g2_mux2_1 _27427_ (.A0(net6365),
    .A1(net4733),
    .S(_08390_),
    .X(_02753_));
 sg13g2_mux2_1 _27428_ (.A0(net6337),
    .A1(net6977),
    .S(_08390_),
    .X(_02754_));
 sg13g2_mux2_1 _27429_ (.A0(net6306),
    .A1(net4799),
    .S(_08390_),
    .X(_02755_));
 sg13g2_mux2_1 _27430_ (.A0(net6278),
    .A1(net4710),
    .S(_08390_),
    .X(_02756_));
 sg13g2_nand2_2 _27431_ (.Y(_08391_),
    .A(_08251_),
    .B(net5955));
 sg13g2_mux2_1 _27432_ (.A0(net6452),
    .A1(net6975),
    .S(_08391_),
    .X(_02757_));
 sg13g2_mux2_1 _27433_ (.A0(net6423),
    .A1(net4874),
    .S(_08391_),
    .X(_02758_));
 sg13g2_mux2_1 _27434_ (.A0(net6394),
    .A1(net4591),
    .S(_08391_),
    .X(_02759_));
 sg13g2_mux2_1 _27435_ (.A0(net6365),
    .A1(net6920),
    .S(_08391_),
    .X(_02760_));
 sg13g2_mux2_1 _27436_ (.A0(net6337),
    .A1(net4827),
    .S(_08391_),
    .X(_02761_));
 sg13g2_mux2_1 _27437_ (.A0(net6306),
    .A1(net4624),
    .S(_08391_),
    .X(_02762_));
 sg13g2_mux2_1 _27438_ (.A0(net6278),
    .A1(net6792),
    .S(_08391_),
    .X(_02763_));
 sg13g2_nand2_2 _27439_ (.Y(_08392_),
    .A(net5955),
    .B(_08293_));
 sg13g2_mux2_1 _27440_ (.A0(net6452),
    .A1(net4657),
    .S(_08392_),
    .X(_02764_));
 sg13g2_mux2_1 _27441_ (.A0(net6423),
    .A1(net7007),
    .S(_08392_),
    .X(_02765_));
 sg13g2_mux2_1 _27442_ (.A0(net6394),
    .A1(net6680),
    .S(_08392_),
    .X(_02766_));
 sg13g2_mux2_1 _27443_ (.A0(net6365),
    .A1(net4614),
    .S(_08392_),
    .X(_02767_));
 sg13g2_mux2_1 _27444_ (.A0(net6335),
    .A1(net6634),
    .S(_08392_),
    .X(_02768_));
 sg13g2_mux2_1 _27445_ (.A0(net6306),
    .A1(net6740),
    .S(_08392_),
    .X(_02769_));
 sg13g2_mux2_1 _27446_ (.A0(net6278),
    .A1(net6944),
    .S(_08392_),
    .X(_02770_));
 sg13g2_nand2_2 _27447_ (.Y(_08393_),
    .A(_08236_),
    .B(net5955));
 sg13g2_mux2_1 _27448_ (.A0(net6452),
    .A1(net6760),
    .S(_08393_),
    .X(_02771_));
 sg13g2_mux2_1 _27449_ (.A0(net6423),
    .A1(net7092),
    .S(_08393_),
    .X(_02772_));
 sg13g2_mux2_1 _27450_ (.A0(net6394),
    .A1(net6632),
    .S(_08393_),
    .X(_02773_));
 sg13g2_mux2_1 _27451_ (.A0(net6365),
    .A1(net4703),
    .S(_08393_),
    .X(_02774_));
 sg13g2_mux2_1 _27452_ (.A0(net6337),
    .A1(net6653),
    .S(_08393_),
    .X(_02775_));
 sg13g2_mux2_1 _27453_ (.A0(net6306),
    .A1(net6966),
    .S(_08393_),
    .X(_02776_));
 sg13g2_mux2_1 _27454_ (.A0(net6278),
    .A1(net4542),
    .S(_08393_),
    .X(_02777_));
 sg13g2_nand2_2 _27455_ (.Y(_08394_),
    .A(net5956),
    .B(net5950));
 sg13g2_mux2_1 _27456_ (.A0(net6453),
    .A1(net4685),
    .S(_08394_),
    .X(_02778_));
 sg13g2_mux2_1 _27457_ (.A0(net6424),
    .A1(net4922),
    .S(_08394_),
    .X(_02779_));
 sg13g2_mux2_1 _27458_ (.A0(net6395),
    .A1(net7054),
    .S(_08394_),
    .X(_02780_));
 sg13g2_mux2_1 _27459_ (.A0(net6367),
    .A1(net4558),
    .S(_08394_),
    .X(_02781_));
 sg13g2_mux2_1 _27460_ (.A0(net6338),
    .A1(net6842),
    .S(_08394_),
    .X(_02782_));
 sg13g2_mux2_1 _27461_ (.A0(net6308),
    .A1(net6992),
    .S(_08394_),
    .X(_02783_));
 sg13g2_mux2_1 _27462_ (.A0(net6283),
    .A1(net4731),
    .S(_08394_),
    .X(_02784_));
 sg13g2_nand2_2 _27463_ (.Y(_08395_),
    .A(_03131_),
    .B(net5955));
 sg13g2_mux2_1 _27464_ (.A0(net6453),
    .A1(net4824),
    .S(_08395_),
    .X(_02785_));
 sg13g2_mux2_1 _27465_ (.A0(net6424),
    .A1(net6637),
    .S(_08395_),
    .X(_02786_));
 sg13g2_mux2_1 _27466_ (.A0(net6394),
    .A1(net4889),
    .S(_08395_),
    .X(_02787_));
 sg13g2_mux2_1 _27467_ (.A0(net6367),
    .A1(net4618),
    .S(_08395_),
    .X(_02788_));
 sg13g2_mux2_1 _27468_ (.A0(net6337),
    .A1(net4923),
    .S(_08395_),
    .X(_02789_));
 sg13g2_mux2_1 _27469_ (.A0(net6308),
    .A1(net4926),
    .S(_08395_),
    .X(_02790_));
 sg13g2_mux2_1 _27470_ (.A0(net6283),
    .A1(net6994),
    .S(_08395_),
    .X(_02791_));
 sg13g2_nand2_2 _27471_ (.Y(_08396_),
    .A(net5955),
    .B(_08274_));
 sg13g2_mux2_1 _27472_ (.A0(net6453),
    .A1(net4666),
    .S(_08396_),
    .X(_02792_));
 sg13g2_mux2_1 _27473_ (.A0(net6424),
    .A1(net6823),
    .S(_08396_),
    .X(_02793_));
 sg13g2_mux2_1 _27474_ (.A0(net6394),
    .A1(net6785),
    .S(_08396_),
    .X(_02794_));
 sg13g2_mux2_1 _27475_ (.A0(net6367),
    .A1(net6903),
    .S(_08396_),
    .X(_02795_));
 sg13g2_mux2_1 _27476_ (.A0(net6338),
    .A1(net6677),
    .S(_08396_),
    .X(_02796_));
 sg13g2_mux2_1 _27477_ (.A0(net6308),
    .A1(net6921),
    .S(_08396_),
    .X(_02797_));
 sg13g2_mux2_1 _27478_ (.A0(net6283),
    .A1(net6997),
    .S(_08396_),
    .X(_02798_));
 sg13g2_nor2_2 _27479_ (.A(_03128_),
    .B(net5965),
    .Y(_08397_));
 sg13g2_mux2_1 _27480_ (.A0(net4223),
    .A1(net6454),
    .S(_08397_),
    .X(_02799_));
 sg13g2_mux2_1 _27481_ (.A0(net3915),
    .A1(net6425),
    .S(_08397_),
    .X(_02800_));
 sg13g2_mux2_1 _27482_ (.A0(net3516),
    .A1(net6396),
    .S(_08397_),
    .X(_02801_));
 sg13g2_mux2_1 _27483_ (.A0(net3735),
    .A1(net6365),
    .S(_08397_),
    .X(_02802_));
 sg13g2_mux2_1 _27484_ (.A0(net3542),
    .A1(net6335),
    .S(_08397_),
    .X(_02803_));
 sg13g2_mux2_1 _27485_ (.A0(net3804),
    .A1(net6306),
    .S(_08397_),
    .X(_02804_));
 sg13g2_mux2_1 _27486_ (.A0(net3975),
    .A1(net6277),
    .S(_08397_),
    .X(_02805_));
 sg13g2_nand2_2 _27487_ (.Y(_08398_),
    .A(net5955),
    .B(_08278_));
 sg13g2_mux2_1 _27488_ (.A0(net6452),
    .A1(net6852),
    .S(_08398_),
    .X(_02806_));
 sg13g2_mux2_1 _27489_ (.A0(net6423),
    .A1(net6707),
    .S(_08398_),
    .X(_02807_));
 sg13g2_mux2_1 _27490_ (.A0(net6395),
    .A1(net6797),
    .S(_08398_),
    .X(_02808_));
 sg13g2_mux2_1 _27491_ (.A0(net6373),
    .A1(net7077),
    .S(_08398_),
    .X(_02809_));
 sg13g2_mux2_1 _27492_ (.A0(net6344),
    .A1(net6664),
    .S(_08398_),
    .X(_02810_));
 sg13g2_mux2_1 _27493_ (.A0(net6313),
    .A1(net6784),
    .S(_08398_),
    .X(_02811_));
 sg13g2_mux2_1 _27494_ (.A0(net6282),
    .A1(net4669),
    .S(_08398_),
    .X(_02812_));
 sg13g2_nor2_2 _27495_ (.A(net5965),
    .B(_08266_),
    .Y(_08399_));
 sg13g2_mux2_1 _27496_ (.A0(net4374),
    .A1(net6452),
    .S(_08399_),
    .X(_02813_));
 sg13g2_mux2_1 _27497_ (.A0(net4356),
    .A1(net6423),
    .S(_08399_),
    .X(_02814_));
 sg13g2_mux2_1 _27498_ (.A0(net4343),
    .A1(net6395),
    .S(_08399_),
    .X(_02815_));
 sg13g2_mux2_1 _27499_ (.A0(net3886),
    .A1(net6373),
    .S(_08399_),
    .X(_02816_));
 sg13g2_mux2_1 _27500_ (.A0(net3580),
    .A1(net6344),
    .S(_08399_),
    .X(_02817_));
 sg13g2_mux2_1 _27501_ (.A0(net3584),
    .A1(net6313),
    .S(_08399_),
    .X(_02818_));
 sg13g2_mux2_1 _27502_ (.A0(net4203),
    .A1(net6282),
    .S(_08399_),
    .X(_02819_));
 sg13g2_nor2_2 _27503_ (.A(_08266_),
    .B(net5952),
    .Y(_08400_));
 sg13g2_mux2_1 _27504_ (.A0(net3841),
    .A1(net6453),
    .S(_08400_),
    .X(_02820_));
 sg13g2_mux2_1 _27505_ (.A0(net3994),
    .A1(net6423),
    .S(_08400_),
    .X(_02821_));
 sg13g2_mux2_1 _27506_ (.A0(net3999),
    .A1(net6395),
    .S(_08400_),
    .X(_02822_));
 sg13g2_mux2_1 _27507_ (.A0(net3501),
    .A1(net6373),
    .S(_08400_),
    .X(_02823_));
 sg13g2_mux2_1 _27508_ (.A0(net3497),
    .A1(net6344),
    .S(_08400_),
    .X(_02824_));
 sg13g2_mux2_1 _27509_ (.A0(net3967),
    .A1(net6313),
    .S(_08400_),
    .X(_02825_));
 sg13g2_mux2_1 _27510_ (.A0(net4106),
    .A1(net6282),
    .S(_08400_),
    .X(_02826_));
 sg13g2_nor2_2 _27511_ (.A(net6029),
    .B(_08266_),
    .Y(_08401_));
 sg13g2_mux2_1 _27512_ (.A0(net4399),
    .A1(net6452),
    .S(_08401_),
    .X(_02827_));
 sg13g2_mux2_1 _27513_ (.A0(net4113),
    .A1(net6423),
    .S(_08401_),
    .X(_02828_));
 sg13g2_mux2_1 _27514_ (.A0(net4034),
    .A1(net6395),
    .S(_08401_),
    .X(_02829_));
 sg13g2_mux2_1 _27515_ (.A0(net4260),
    .A1(net6373),
    .S(_08401_),
    .X(_02830_));
 sg13g2_mux2_1 _27516_ (.A0(net4194),
    .A1(net6344),
    .S(_08401_),
    .X(_02831_));
 sg13g2_mux2_1 _27517_ (.A0(net4102),
    .A1(net6313),
    .S(_08401_),
    .X(_02832_));
 sg13g2_mux2_1 _27518_ (.A0(net3931),
    .A1(net6282),
    .S(_08401_),
    .X(_02833_));
 sg13g2_nand2_2 _27519_ (.Y(_08402_),
    .A(net5969),
    .B(_08269_));
 sg13g2_mux2_1 _27520_ (.A0(net6461),
    .A1(net6706),
    .S(_08402_),
    .X(_02834_));
 sg13g2_mux2_1 _27521_ (.A0(net6431),
    .A1(net4828),
    .S(_08402_),
    .X(_02835_));
 sg13g2_mux2_1 _27522_ (.A0(net6402),
    .A1(net4782),
    .S(_08402_),
    .X(_02836_));
 sg13g2_mux2_1 _27523_ (.A0(net6375),
    .A1(net6684),
    .S(_08402_),
    .X(_02837_));
 sg13g2_mux2_1 _27524_ (.A0(net6347),
    .A1(net6795),
    .S(_08402_),
    .X(_02838_));
 sg13g2_mux2_1 _27525_ (.A0(net6314),
    .A1(net4853),
    .S(_08402_),
    .X(_02839_));
 sg13g2_mux2_1 _27526_ (.A0(net6286),
    .A1(net6696),
    .S(_08402_),
    .X(_02840_));
 sg13g2_nand2_2 _27527_ (.Y(_08403_),
    .A(net5962),
    .B(_08269_));
 sg13g2_mux2_1 _27528_ (.A0(net6461),
    .A1(net7090),
    .S(_08403_),
    .X(_02841_));
 sg13g2_mux2_1 _27529_ (.A0(net6431),
    .A1(net6622),
    .S(_08403_),
    .X(_02842_));
 sg13g2_mux2_1 _27530_ (.A0(net6402),
    .A1(net4648),
    .S(_08403_),
    .X(_02843_));
 sg13g2_mux2_1 _27531_ (.A0(net6375),
    .A1(net4936),
    .S(_08403_),
    .X(_02844_));
 sg13g2_mux2_1 _27532_ (.A0(net6343),
    .A1(net4674),
    .S(_08403_),
    .X(_02845_));
 sg13g2_mux2_1 _27533_ (.A0(net6314),
    .A1(net7079),
    .S(_08403_),
    .X(_02846_));
 sg13g2_mux2_1 _27534_ (.A0(net6286),
    .A1(net6818),
    .S(_08403_),
    .X(_02847_));
 sg13g2_nand2_2 _27535_ (.Y(_08404_),
    .A(_08269_),
    .B(net5953));
 sg13g2_mux2_1 _27536_ (.A0(net6461),
    .A1(net6675),
    .S(_08404_),
    .X(_02848_));
 sg13g2_mux2_1 _27537_ (.A0(net6431),
    .A1(net6657),
    .S(_08404_),
    .X(_02849_));
 sg13g2_mux2_1 _27538_ (.A0(net6402),
    .A1(net6781),
    .S(_08404_),
    .X(_02850_));
 sg13g2_mux2_1 _27539_ (.A0(net6375),
    .A1(net7044),
    .S(_08404_),
    .X(_02851_));
 sg13g2_mux2_1 _27540_ (.A0(net6346),
    .A1(net6967),
    .S(_08404_),
    .X(_02852_));
 sg13g2_mux2_1 _27541_ (.A0(net6314),
    .A1(net4695),
    .S(_08404_),
    .X(_02853_));
 sg13g2_mux2_1 _27542_ (.A0(net6286),
    .A1(net6887),
    .S(_08404_),
    .X(_02854_));
 sg13g2_nand2_2 _27543_ (.Y(_08405_),
    .A(net5968),
    .B(_08269_));
 sg13g2_mux2_1 _27544_ (.A0(net6461),
    .A1(net6761),
    .S(_08405_),
    .X(_02855_));
 sg13g2_mux2_1 _27545_ (.A0(net6433),
    .A1(net4607),
    .S(_08405_),
    .X(_02856_));
 sg13g2_mux2_1 _27546_ (.A0(net6402),
    .A1(net6699),
    .S(_08405_),
    .X(_02857_));
 sg13g2_mux2_1 _27547_ (.A0(net6375),
    .A1(net6831),
    .S(_08405_),
    .X(_02858_));
 sg13g2_mux2_1 _27548_ (.A0(net6346),
    .A1(net4897),
    .S(_08405_),
    .X(_02859_));
 sg13g2_mux2_1 _27549_ (.A0(net6314),
    .A1(net4707),
    .S(_08405_),
    .X(_02860_));
 sg13g2_mux2_1 _27550_ (.A0(net6286),
    .A1(net4860),
    .S(_08405_),
    .X(_02861_));
 sg13g2_nand2_2 _27551_ (.Y(_08406_),
    .A(_08269_),
    .B(net5951));
 sg13g2_mux2_1 _27552_ (.A0(net6460),
    .A1(net4683),
    .S(_08406_),
    .X(_02862_));
 sg13g2_mux2_1 _27553_ (.A0(net6432),
    .A1(net6840),
    .S(_08406_),
    .X(_02863_));
 sg13g2_mux2_1 _27554_ (.A0(net6401),
    .A1(net6952),
    .S(_08406_),
    .X(_02864_));
 sg13g2_mux2_1 _27555_ (.A0(net6374),
    .A1(net4532),
    .S(_08406_),
    .X(_02865_));
 sg13g2_mux2_1 _27556_ (.A0(net6345),
    .A1(net4775),
    .S(_08406_),
    .X(_02866_));
 sg13g2_mux2_1 _27557_ (.A0(net6315),
    .A1(net4531),
    .S(_08406_),
    .X(_02867_));
 sg13g2_mux2_1 _27558_ (.A0(net6284),
    .A1(net4801),
    .S(_08406_),
    .X(_02868_));
 sg13g2_nor2_2 _27559_ (.A(_03128_),
    .B(net5952),
    .Y(_08407_));
 sg13g2_mux2_1 _27560_ (.A0(net3680),
    .A1(net6454),
    .S(_08407_),
    .X(_02869_));
 sg13g2_mux2_1 _27561_ (.A0(net4021),
    .A1(net6425),
    .S(_08407_),
    .X(_02870_));
 sg13g2_mux2_1 _27562_ (.A0(net3831),
    .A1(net6396),
    .S(_08407_),
    .X(_02871_));
 sg13g2_mux2_1 _27563_ (.A0(net3646),
    .A1(net6365),
    .S(_08407_),
    .X(_02872_));
 sg13g2_mux2_1 _27564_ (.A0(net3743),
    .A1(net6335),
    .S(_08407_),
    .X(_02873_));
 sg13g2_mux2_1 _27565_ (.A0(net4107),
    .A1(net6306),
    .S(_08407_),
    .X(_02874_));
 sg13g2_mux2_1 _27566_ (.A0(net3731),
    .A1(net6277),
    .S(_08407_),
    .X(_02875_));
 sg13g2_nor2_2 _27567_ (.A(_08270_),
    .B(_08294_),
    .Y(_08408_));
 sg13g2_mux2_1 _27568_ (.A0(net4412),
    .A1(net6460),
    .S(_08408_),
    .X(_02876_));
 sg13g2_mux2_1 _27569_ (.A0(net3426),
    .A1(net6432),
    .S(_08408_),
    .X(_02877_));
 sg13g2_mux2_1 _27570_ (.A0(net4128),
    .A1(net6401),
    .S(_08408_),
    .X(_02878_));
 sg13g2_mux2_1 _27571_ (.A0(net3840),
    .A1(net6374),
    .S(_08408_),
    .X(_02879_));
 sg13g2_mux2_1 _27572_ (.A0(net4213),
    .A1(net6345),
    .S(_08408_),
    .X(_02880_));
 sg13g2_mux2_1 _27573_ (.A0(net4401),
    .A1(net6315),
    .S(_08408_),
    .X(_02881_));
 sg13g2_mux2_1 _27574_ (.A0(net4085),
    .A1(net6285),
    .S(_08408_),
    .X(_02882_));
 sg13g2_nor2_2 _27575_ (.A(_08237_),
    .B(net5954),
    .Y(_08409_));
 sg13g2_mux2_1 _27576_ (.A0(net3948),
    .A1(net6460),
    .S(_08409_),
    .X(_02883_));
 sg13g2_mux2_1 _27577_ (.A0(net4136),
    .A1(net6432),
    .S(_08409_),
    .X(_02884_));
 sg13g2_mux2_1 _27578_ (.A0(net4066),
    .A1(net6401),
    .S(_08409_),
    .X(_02885_));
 sg13g2_mux2_1 _27579_ (.A0(net4172),
    .A1(net6374),
    .S(_08409_),
    .X(_02886_));
 sg13g2_mux2_1 _27580_ (.A0(net3768),
    .A1(net6345),
    .S(_08409_),
    .X(_02887_));
 sg13g2_mux2_1 _27581_ (.A0(net3866),
    .A1(net6315),
    .S(_08409_),
    .X(_02888_));
 sg13g2_mux2_1 _27582_ (.A0(net3503),
    .A1(net6285),
    .S(_08409_),
    .X(_02889_));
 sg13g2_nand2_2 _27583_ (.Y(_08410_),
    .A(_08269_),
    .B(net5950));
 sg13g2_mux2_1 _27584_ (.A0(net6459),
    .A1(net6770),
    .S(_08410_),
    .X(_02890_));
 sg13g2_mux2_1 _27585_ (.A0(net6433),
    .A1(net4826),
    .S(_08410_),
    .X(_02891_));
 sg13g2_mux2_1 _27586_ (.A0(net6402),
    .A1(net4746),
    .S(_08410_),
    .X(_02892_));
 sg13g2_mux2_1 _27587_ (.A0(net6376),
    .A1(net4571),
    .S(_08410_),
    .X(_02893_));
 sg13g2_mux2_1 _27588_ (.A0(net6343),
    .A1(net4734),
    .S(_08410_),
    .X(_02894_));
 sg13g2_mux2_1 _27589_ (.A0(net6314),
    .A1(net6890),
    .S(_08410_),
    .X(_02895_));
 sg13g2_mux2_1 _27590_ (.A0(net6284),
    .A1(net4821),
    .S(_08410_),
    .X(_02896_));
 sg13g2_nor2_2 _27591_ (.A(_03132_),
    .B(net5954),
    .Y(_08411_));
 sg13g2_mux2_1 _27592_ (.A0(net3805),
    .A1(net6459),
    .S(_08411_),
    .X(_02897_));
 sg13g2_mux2_1 _27593_ (.A0(net4359),
    .A1(net6433),
    .S(_08411_),
    .X(_02898_));
 sg13g2_mux2_1 _27594_ (.A0(net4039),
    .A1(net6403),
    .S(_08411_),
    .X(_02899_));
 sg13g2_mux2_1 _27595_ (.A0(net4207),
    .A1(net6376),
    .S(_08411_),
    .X(_02900_));
 sg13g2_mux2_1 _27596_ (.A0(net4117),
    .A1(net6343),
    .S(_08411_),
    .X(_02901_));
 sg13g2_mux2_1 _27597_ (.A0(net3481),
    .A1(net6314),
    .S(_08411_),
    .X(_02902_));
 sg13g2_mux2_1 _27598_ (.A0(net4024),
    .A1(net6284),
    .S(_08411_),
    .X(_02903_));
 sg13g2_nor2_2 _27599_ (.A(net5954),
    .B(_08275_),
    .Y(_08412_));
 sg13g2_mux2_1 _27600_ (.A0(net3934),
    .A1(net6459),
    .S(_08412_),
    .X(_02904_));
 sg13g2_mux2_1 _27601_ (.A0(net4308),
    .A1(net6433),
    .S(_08412_),
    .X(_02905_));
 sg13g2_mux2_1 _27602_ (.A0(net3627),
    .A1(net6402),
    .S(_08412_),
    .X(_02906_));
 sg13g2_mux2_1 _27603_ (.A0(net3942),
    .A1(net6375),
    .S(_08412_),
    .X(_02907_));
 sg13g2_mux2_1 _27604_ (.A0(net3857),
    .A1(net6343),
    .S(_08412_),
    .X(_02908_));
 sg13g2_mux2_1 _27605_ (.A0(net3855),
    .A1(net6314),
    .S(_08412_),
    .X(_02909_));
 sg13g2_mux2_1 _27606_ (.A0(net4111),
    .A1(net6284),
    .S(_08412_),
    .X(_02910_));
 sg13g2_nor2_2 _27607_ (.A(_08246_),
    .B(net5954),
    .Y(_08413_));
 sg13g2_mux2_1 _27608_ (.A0(net3859),
    .A1(net6459),
    .S(_08413_),
    .X(_02911_));
 sg13g2_mux2_1 _27609_ (.A0(net4446),
    .A1(net6433),
    .S(_08413_),
    .X(_02912_));
 sg13g2_mux2_1 _27610_ (.A0(net4417),
    .A1(net6403),
    .S(_08413_),
    .X(_02913_));
 sg13g2_mux2_1 _27611_ (.A0(net4170),
    .A1(net6375),
    .S(_08413_),
    .X(_02914_));
 sg13g2_mux2_1 _27612_ (.A0(net4171),
    .A1(net6343),
    .S(_08413_),
    .X(_02915_));
 sg13g2_mux2_1 _27613_ (.A0(net4280),
    .A1(net6315),
    .S(_08413_),
    .X(_02916_));
 sg13g2_mux2_1 _27614_ (.A0(net4004),
    .A1(net6284),
    .S(_08413_),
    .X(_02917_));
 sg13g2_nor2_2 _27615_ (.A(net5954),
    .B(_08279_),
    .Y(_08414_));
 sg13g2_mux2_1 _27616_ (.A0(net4272),
    .A1(net6459),
    .S(_08414_),
    .X(_02918_));
 sg13g2_mux2_1 _27617_ (.A0(net3616),
    .A1(net6431),
    .S(_08414_),
    .X(_02919_));
 sg13g2_mux2_1 _27618_ (.A0(net4229),
    .A1(net6401),
    .S(_08414_),
    .X(_02920_));
 sg13g2_mux2_1 _27619_ (.A0(net4281),
    .A1(net6373),
    .S(_08414_),
    .X(_02921_));
 sg13g2_mux2_1 _27620_ (.A0(net4139),
    .A1(net6343),
    .S(_08414_),
    .X(_02922_));
 sg13g2_mux2_1 _27621_ (.A0(net3508),
    .A1(net6316),
    .S(_08414_),
    .X(_02923_));
 sg13g2_mux2_1 _27622_ (.A0(net4749),
    .A1(net6282),
    .S(_08414_),
    .X(_02924_));
 sg13g2_nor2_2 _27623_ (.A(net5965),
    .B(net5954),
    .Y(_08415_));
 sg13g2_mux2_1 _27624_ (.A0(net4023),
    .A1(net6459),
    .S(_08415_),
    .X(_02925_));
 sg13g2_mux2_1 _27625_ (.A0(net4394),
    .A1(net6431),
    .S(_08415_),
    .X(_02926_));
 sg13g2_mux2_1 _27626_ (.A0(net3806),
    .A1(net6401),
    .S(_08415_),
    .X(_02927_));
 sg13g2_mux2_1 _27627_ (.A0(net4126),
    .A1(net6373),
    .S(_08415_),
    .X(_02928_));
 sg13g2_mux2_1 _27628_ (.A0(net3985),
    .A1(net6343),
    .S(_08415_),
    .X(_02929_));
 sg13g2_mux2_1 _27629_ (.A0(net4445),
    .A1(net6313),
    .S(_08415_),
    .X(_02930_));
 sg13g2_mux2_1 _27630_ (.A0(net3950),
    .A1(net6284),
    .S(_08415_),
    .X(_02931_));
 sg13g2_nor2_2 _27631_ (.A(net5954),
    .B(net5952),
    .Y(_08416_));
 sg13g2_mux2_1 _27632_ (.A0(net4137),
    .A1(net6459),
    .S(_08416_),
    .X(_02932_));
 sg13g2_mux2_1 _27633_ (.A0(net3378),
    .A1(net6431),
    .S(_08416_),
    .X(_02933_));
 sg13g2_mux2_1 _27634_ (.A0(net4123),
    .A1(net6401),
    .S(_08416_),
    .X(_02934_));
 sg13g2_mux2_1 _27635_ (.A0(net4264),
    .A1(net6373),
    .S(_08416_),
    .X(_02935_));
 sg13g2_mux2_1 _27636_ (.A0(net3441),
    .A1(net6343),
    .S(_08416_),
    .X(_02936_));
 sg13g2_mux2_1 _27637_ (.A0(net4160),
    .A1(net6313),
    .S(_08416_),
    .X(_02937_));
 sg13g2_mux2_1 _27638_ (.A0(net3682),
    .A1(net6284),
    .S(_08416_),
    .X(_02938_));
 sg13g2_nor2_2 _27639_ (.A(net6029),
    .B(_03128_),
    .Y(_08417_));
 sg13g2_mux2_1 _27640_ (.A0(net4037),
    .A1(net6454),
    .S(_08417_),
    .X(_02939_));
 sg13g2_mux2_1 _27641_ (.A0(net4396),
    .A1(net6425),
    .S(_08417_),
    .X(_02940_));
 sg13g2_mux2_1 _27642_ (.A0(net4177),
    .A1(net6396),
    .S(_08417_),
    .X(_02941_));
 sg13g2_mux2_1 _27643_ (.A0(net4129),
    .A1(net6365),
    .S(_08417_),
    .X(_02942_));
 sg13g2_mux2_1 _27644_ (.A0(net4271),
    .A1(net6335),
    .S(_08417_),
    .X(_02943_));
 sg13g2_mux2_1 _27645_ (.A0(net3986),
    .A1(net6307),
    .S(_08417_),
    .X(_02944_));
 sg13g2_mux2_1 _27646_ (.A0(net3513),
    .A1(net6277),
    .S(_08417_),
    .X(_02945_));
 sg13g2_nand2_2 _27647_ (.Y(_08418_),
    .A(net5969),
    .B(net5966));
 sg13g2_mux2_1 _27648_ (.A0(net6466),
    .A1(net4487),
    .S(_08418_),
    .X(_02946_));
 sg13g2_mux2_1 _27649_ (.A0(net6437),
    .A1(net6624),
    .S(_08418_),
    .X(_02947_));
 sg13g2_mux2_1 _27650_ (.A0(net6405),
    .A1(net4579),
    .S(_08418_),
    .X(_02948_));
 sg13g2_mux2_1 _27651_ (.A0(net6378),
    .A1(net4848),
    .S(_08418_),
    .X(_02949_));
 sg13g2_mux2_1 _27652_ (.A0(net6350),
    .A1(net4869),
    .S(_08418_),
    .X(_02950_));
 sg13g2_mux2_1 _27653_ (.A0(net6319),
    .A1(net6606),
    .S(_08418_),
    .X(_02951_));
 sg13g2_mux2_1 _27654_ (.A0(net6289),
    .A1(net4946),
    .S(_08418_),
    .X(_02952_));
 sg13g2_nand2_2 _27655_ (.Y(_08419_),
    .A(net5966),
    .B(net5962));
 sg13g2_mux2_1 _27656_ (.A0(net6466),
    .A1(net4795),
    .S(_08419_),
    .X(_02953_));
 sg13g2_mux2_1 _27657_ (.A0(net6434),
    .A1(net6721),
    .S(_08419_),
    .X(_02954_));
 sg13g2_mux2_1 _27658_ (.A0(net6405),
    .A1(net6861),
    .S(_08419_),
    .X(_02955_));
 sg13g2_mux2_1 _27659_ (.A0(net6378),
    .A1(net6701),
    .S(_08419_),
    .X(_02956_));
 sg13g2_mux2_1 _27660_ (.A0(net6350),
    .A1(net6867),
    .S(_08419_),
    .X(_02957_));
 sg13g2_mux2_1 _27661_ (.A0(net6319),
    .A1(net4745),
    .S(_08419_),
    .X(_02958_));
 sg13g2_mux2_1 _27662_ (.A0(net6289),
    .A1(net6897),
    .S(_08419_),
    .X(_02959_));
 sg13g2_nand2_2 _27663_ (.Y(_08420_),
    .A(net5966),
    .B(net5953));
 sg13g2_mux2_1 _27664_ (.A0(net6463),
    .A1(net7133),
    .S(_08420_),
    .X(_02960_));
 sg13g2_mux2_1 _27665_ (.A0(net6434),
    .A1(net6988),
    .S(_08420_),
    .X(_02961_));
 sg13g2_mux2_1 _27666_ (.A0(net6405),
    .A1(net7110),
    .S(_08420_),
    .X(_02962_));
 sg13g2_mux2_1 _27667_ (.A0(net6378),
    .A1(net6877),
    .S(_08420_),
    .X(_02963_));
 sg13g2_mux2_1 _27668_ (.A0(net6350),
    .A1(net4706),
    .S(_08420_),
    .X(_02964_));
 sg13g2_mux2_1 _27669_ (.A0(net6319),
    .A1(net6983),
    .S(_08420_),
    .X(_02965_));
 sg13g2_mux2_1 _27670_ (.A0(net6290),
    .A1(net6775),
    .S(_08420_),
    .X(_02966_));
 sg13g2_nand2_2 _27671_ (.Y(_08421_),
    .A(net6027),
    .B(net5962));
 sg13g2_mux2_1 _27672_ (.A0(net6455),
    .A1(net6853),
    .S(_08421_),
    .X(_02967_));
 sg13g2_mux2_1 _27673_ (.A0(net6426),
    .A1(net6649),
    .S(_08421_),
    .X(_02968_));
 sg13g2_mux2_1 _27674_ (.A0(net6397),
    .A1(net6971),
    .S(_08421_),
    .X(_02969_));
 sg13g2_mux2_1 _27675_ (.A0(net6368),
    .A1(net6841),
    .S(_08421_),
    .X(_02970_));
 sg13g2_mux2_1 _27676_ (.A0(net6341),
    .A1(net6938),
    .S(_08421_),
    .X(_02971_));
 sg13g2_mux2_1 _27677_ (.A0(net6309),
    .A1(net6663),
    .S(_08421_),
    .X(_02972_));
 sg13g2_mux2_1 _27678_ (.A0(net6279),
    .A1(net4925),
    .S(_08421_),
    .X(_02973_));
 sg13g2_nand2_2 _27679_ (.Y(_08422_),
    .A(net5967),
    .B(net5951));
 sg13g2_mux2_1 _27680_ (.A0(net6467),
    .A1(net4546),
    .S(_08422_),
    .X(_02974_));
 sg13g2_mux2_1 _27681_ (.A0(net6438),
    .A1(net4554),
    .S(_08422_),
    .X(_02975_));
 sg13g2_mux2_1 _27682_ (.A0(net6408),
    .A1(net4573),
    .S(_08422_),
    .X(_02976_));
 sg13g2_mux2_1 _27683_ (.A0(net6381),
    .A1(net6745),
    .S(_08422_),
    .X(_02977_));
 sg13g2_mux2_1 _27684_ (.A0(net6351),
    .A1(net6993),
    .S(_08422_),
    .X(_02978_));
 sg13g2_mux2_1 _27685_ (.A0(net6322),
    .A1(net7063),
    .S(_08422_),
    .X(_02979_));
 sg13g2_mux2_1 _27686_ (.A0(net6291),
    .A1(net7080),
    .S(_08422_),
    .X(_02980_));
 sg13g2_nand2_2 _27687_ (.Y(_08423_),
    .A(net5967),
    .B(_08251_));
 sg13g2_mux2_1 _27688_ (.A0(net6467),
    .A1(net6814),
    .S(_08423_),
    .X(_02981_));
 sg13g2_mux2_1 _27689_ (.A0(net6438),
    .A1(net6780),
    .S(_08423_),
    .X(_02982_));
 sg13g2_mux2_1 _27690_ (.A0(net6408),
    .A1(net4810),
    .S(_08423_),
    .X(_02983_));
 sg13g2_mux2_1 _27691_ (.A0(net6381),
    .A1(net4728),
    .S(_08423_),
    .X(_02984_));
 sg13g2_mux2_1 _27692_ (.A0(net6351),
    .A1(net4565),
    .S(_08423_),
    .X(_02985_));
 sg13g2_mux2_1 _27693_ (.A0(net6322),
    .A1(net4924),
    .S(_08423_),
    .X(_02986_));
 sg13g2_mux2_1 _27694_ (.A0(net6291),
    .A1(net4634),
    .S(_08423_),
    .X(_02987_));
 sg13g2_nand2_2 _27695_ (.Y(_08424_),
    .A(net5967),
    .B(_08293_));
 sg13g2_mux2_1 _27696_ (.A0(net6467),
    .A1(net4783),
    .S(_08424_),
    .X(_02988_));
 sg13g2_mux2_1 _27697_ (.A0(net6438),
    .A1(net6791),
    .S(_08424_),
    .X(_02989_));
 sg13g2_mux2_1 _27698_ (.A0(net6408),
    .A1(net6973),
    .S(_08424_),
    .X(_02990_));
 sg13g2_mux2_1 _27699_ (.A0(net6381),
    .A1(net6949),
    .S(_08424_),
    .X(_02991_));
 sg13g2_mux2_1 _27700_ (.A0(net6351),
    .A1(net6998),
    .S(_08424_),
    .X(_02992_));
 sg13g2_mux2_1 _27701_ (.A0(net6322),
    .A1(net4572),
    .S(_08424_),
    .X(_02993_));
 sg13g2_mux2_1 _27702_ (.A0(net6291),
    .A1(net7022),
    .S(_08424_),
    .X(_02994_));
 sg13g2_nand2_2 _27703_ (.Y(_08425_),
    .A(net5967),
    .B(_08236_));
 sg13g2_mux2_1 _27704_ (.A0(net6467),
    .A1(net6729),
    .S(_08425_),
    .X(_02995_));
 sg13g2_mux2_1 _27705_ (.A0(net6438),
    .A1(net6718),
    .S(_08425_),
    .X(_02996_));
 sg13g2_mux2_1 _27706_ (.A0(net6408),
    .A1(net7021),
    .S(_08425_),
    .X(_02997_));
 sg13g2_mux2_1 _27707_ (.A0(net6381),
    .A1(net4933),
    .S(_08425_),
    .X(_02998_));
 sg13g2_mux2_1 _27708_ (.A0(net6351),
    .A1(net6820),
    .S(_08425_),
    .X(_02999_));
 sg13g2_mux2_1 _27709_ (.A0(net6322),
    .A1(net6635),
    .S(_08425_),
    .X(_03000_));
 sg13g2_mux2_1 _27710_ (.A0(net6291),
    .A1(net6839),
    .S(_08425_),
    .X(_03001_));
 sg13g2_nand2_2 _27711_ (.Y(_08426_),
    .A(net5966),
    .B(net5950));
 sg13g2_mux2_1 _27712_ (.A0(net6467),
    .A1(net4823),
    .S(_08426_),
    .X(_03002_));
 sg13g2_mux2_1 _27713_ (.A0(net6440),
    .A1(net6834),
    .S(_08426_),
    .X(_03003_));
 sg13g2_mux2_1 _27714_ (.A0(net6408),
    .A1(net6786),
    .S(_08426_),
    .X(_03004_));
 sg13g2_mux2_1 _27715_ (.A0(net6381),
    .A1(net4679),
    .S(_08426_),
    .X(_03005_));
 sg13g2_mux2_1 _27716_ (.A0(net6353),
    .A1(net7053),
    .S(_08426_),
    .X(_03006_));
 sg13g2_mux2_1 _27717_ (.A0(net6322),
    .A1(net6902),
    .S(_08426_),
    .X(_03007_));
 sg13g2_mux2_1 _27718_ (.A0(net6291),
    .A1(net4829),
    .S(_08426_),
    .X(_03008_));
 sg13g2_a21oi_1 _27719_ (.A1(_08727_),
    .A2(net5735),
    .Y(_08427_),
    .B1(_08740_));
 sg13g2_nand2_1 _27720_ (.Y(_08428_),
    .A(_07429_),
    .B(_08427_));
 sg13g2_o21ai_1 _27721_ (.B1(_08428_),
    .Y(_08429_),
    .A1(_09018_),
    .A2(_07453_));
 sg13g2_nor3_1 _27722_ (.A(_08740_),
    .B(net5731),
    .C(_07437_),
    .Y(_08430_));
 sg13g2_nor2b_1 _27723_ (.A(net5730),
    .B_N(_08430_),
    .Y(_08431_));
 sg13g2_nor3_1 _27724_ (.A(_07465_),
    .B(_08429_),
    .C(_08431_),
    .Y(_08432_));
 sg13g2_a22oi_1 _27725_ (.Y(_03009_),
    .B1(_07466_),
    .B2(_08432_),
    .A2(net5820),
    .A1(_08577_));
 sg13g2_nor2_1 _27726_ (.A(net7407),
    .B(net5822),
    .Y(_08433_));
 sg13g2_nor3_1 _27727_ (.A(net5733),
    .B(_08991_),
    .C(_07454_),
    .Y(_08434_));
 sg13g2_nor3_1 _27728_ (.A(net5820),
    .B(_08429_),
    .C(_08434_),
    .Y(_08435_));
 sg13g2_o21ai_1 _27729_ (.B1(_08954_),
    .Y(_03010_),
    .A1(_08433_),
    .A2(_08435_));
 sg13g2_nor2_1 _27730_ (.A(net5736),
    .B(net5730),
    .Y(_08436_));
 sg13g2_o21ai_1 _27731_ (.B1(_08436_),
    .Y(_08437_),
    .A1(net5733),
    .A2(_08757_));
 sg13g2_nand3_1 _27732_ (.B(_07460_),
    .C(_08437_),
    .A(_07437_),
    .Y(_08438_));
 sg13g2_nand3_1 _27733_ (.B(net5731),
    .C(_08438_),
    .A(_08739_),
    .Y(_08439_));
 sg13g2_nor3_1 _27734_ (.A(_08835_),
    .B(_08990_),
    .C(_07454_),
    .Y(_08440_));
 sg13g2_nor3_1 _27735_ (.A(_07465_),
    .B(_08430_),
    .C(_08440_),
    .Y(_08441_));
 sg13g2_a22oi_1 _27736_ (.Y(_03011_),
    .B1(_08439_),
    .B2(_08441_),
    .A2(net5820),
    .A1(_08576_));
 sg13g2_a22oi_1 _27737_ (.Y(_03012_),
    .B1(_07472_),
    .B2(_08439_),
    .A2(net5819),
    .A1(_08574_));
 sg13g2_nor3_2 _27738_ (.A(_08746_),
    .B(_08763_),
    .C(_08831_),
    .Y(_08442_));
 sg13g2_a21oi_2 _27739_ (.B1(_08442_),
    .Y(_08443_),
    .A2(_08896_),
    .A1(_08741_));
 sg13g2_a22oi_1 _27740_ (.Y(_03013_),
    .B1(_07434_),
    .B2(_08443_),
    .A2(net5819),
    .A1(_08589_));
 sg13g2_nand4_1 _27741_ (.B(net5731),
    .C(_08989_),
    .A(net5755),
    .Y(_08444_),
    .D(_07420_));
 sg13g2_nand3_1 _27742_ (.B(_07440_),
    .C(_08444_),
    .A(_07439_),
    .Y(_08445_));
 sg13g2_o21ai_1 _27743_ (.B1(_07436_),
    .Y(_08446_),
    .A1(_09018_),
    .A2(_07454_));
 sg13g2_nor3_1 _27744_ (.A(_07464_),
    .B(_08445_),
    .C(_08446_),
    .Y(_08447_));
 sg13g2_a22oi_1 _27745_ (.Y(_03014_),
    .B1(_08443_),
    .B2(_08447_),
    .A2(net5819),
    .A1(_08588_));
 sg13g2_nand2_1 _27746_ (.Y(_08448_),
    .A(_08756_),
    .B(_08442_));
 sg13g2_nor2_1 _27747_ (.A(_07435_),
    .B(_08443_),
    .Y(_08449_));
 sg13g2_a22oi_1 _27748_ (.Y(_03015_),
    .B1(_08448_),
    .B2(_08449_),
    .A2(net5819),
    .A1(_08586_));
 sg13g2_nand3_1 _27749_ (.B(_07434_),
    .C(_08442_),
    .A(net5731),
    .Y(_08450_));
 sg13g2_o21ai_1 _27750_ (.B1(_08450_),
    .Y(_08451_),
    .A1(net7376),
    .A2(net5824));
 sg13g2_inv_1 _27751_ (.Y(_03016_),
    .A(_08451_));
 sg13g2_nand3b_1 _27752_ (.B(_09121_),
    .C(_09125_),
    .Y(_08452_),
    .A_N(_09113_));
 sg13g2_o21ai_1 _27753_ (.B1(\atari2600.tia.vid_ypos[3] ),
    .Y(_08453_),
    .A1(\atari2600.tia.vid_ypos[2] ),
    .A2(_08702_));
 sg13g2_a21o_1 _27754_ (.A2(_08453_),
    .A1(_09643_),
    .B1(_10114_),
    .X(_08454_));
 sg13g2_a21oi_2 _27755_ (.B1(_09343_),
    .Y(_08455_),
    .A2(_08454_),
    .A1(_00130_));
 sg13g2_nand2_1 _27756_ (.Y(_08456_),
    .A(\atari2600.tia.cx[14] ),
    .B(_10063_));
 sg13g2_nand3_1 _27757_ (.B(_04675_),
    .C(_04681_),
    .A(\gamepad_pmod.decoder.data_reg[3] ),
    .Y(_08457_));
 sg13g2_o21ai_1 _27758_ (.B1(_08457_),
    .Y(_08458_),
    .A1(net5),
    .A2(_04675_));
 sg13g2_nor3_2 _27759_ (.A(net5564),
    .B(net5492),
    .C(_08458_),
    .Y(_08459_));
 sg13g2_a221oi_1 _27760_ (.B2(\atari2600.tia.cx[12] ),
    .C1(_08459_),
    .B1(_05374_),
    .A1(\atari2600.tia.cx[2] ),
    .Y(_08460_),
    .A2(_09306_));
 sg13g2_a22oi_1 _27761_ (.Y(_08461_),
    .B1(_09444_),
    .B2(\atari2600.tia.cx[10] ),
    .A2(_09172_),
    .A1(\atari2600.tia.cx[4] ));
 sg13g2_a221oi_1 _27762_ (.B2(\atari2600.tia.cx[1] ),
    .C1(_08455_),
    .B1(_06572_),
    .A1(\atari2600.tia.cx[6] ),
    .Y(_08462_),
    .A2(_09211_));
 sg13g2_nand4_1 _27763_ (.B(_08460_),
    .C(_08461_),
    .A(_08456_),
    .Y(_08463_),
    .D(_08462_));
 sg13g2_a21oi_2 _27764_ (.B1(_08463_),
    .Y(_08464_),
    .A2(_09401_),
    .A1(\atari2600.tia.cx[8] ));
 sg13g2_nor3_1 _27765_ (.A(_09147_),
    .B(net5550),
    .C(net5404),
    .Y(_08465_));
 sg13g2_nor3_1 _27766_ (.A(_08452_),
    .B(_08464_),
    .C(_08465_),
    .Y(_08466_));
 sg13g2_a21o_1 _27767_ (.A2(_08452_),
    .A1(net4341),
    .B1(_08466_),
    .X(_03017_));
 sg13g2_a22oi_1 _27768_ (.Y(_08467_),
    .B1(_10063_),
    .B2(\atari2600.tia.cx[13] ),
    .A2(_09211_),
    .A1(\atari2600.tia.cx[5] ));
 sg13g2_a22oi_1 _27769_ (.Y(_08468_),
    .B1(_06572_),
    .B2(\atari2600.tia.cx[0] ),
    .A2(_09401_),
    .A1(\atari2600.tia.cx[7] ));
 sg13g2_a22oi_1 _27770_ (.Y(_08469_),
    .B1(_09444_),
    .B2(\atari2600.tia.cx[9] ),
    .A2(_09172_),
    .A1(\atari2600.tia.cx[3] ));
 sg13g2_nand3_1 _27771_ (.B(_08468_),
    .C(_08469_),
    .A(_08467_),
    .Y(_08470_));
 sg13g2_a21oi_2 _27772_ (.B1(_08470_),
    .Y(_08471_),
    .A2(_05374_),
    .A1(\atari2600.tia.cx[11] ));
 sg13g2_nor3_1 _27773_ (.A(_08452_),
    .B(_08465_),
    .C(_08471_),
    .Y(_08472_));
 sg13g2_a21o_1 _27774_ (.A2(_08452_),
    .A1(net4423),
    .B1(_08472_),
    .X(_03018_));
 sg13g2_dfrbp_1 _27775_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net98),
    .D(_00177_),
    .Q_N(_13827_),
    .Q(\flash_rom.addr_in[16] ));
 sg13g2_dfrbp_1 _27776_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2699),
    .D(_00178_),
    .Q_N(_13826_),
    .Q(\flash_rom.addr_in[17] ));
 sg13g2_dfrbp_1 _27777_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2698),
    .D(_00179_),
    .Q_N(_13825_),
    .Q(\flash_rom.addr_in[18] ));
 sg13g2_dfrbp_1 _27778_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2697),
    .D(_00180_),
    .Q_N(_13824_),
    .Q(\flash_rom.addr_in[19] ));
 sg13g2_dfrbp_1 _27779_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2696),
    .D(_00181_),
    .Q_N(_13823_),
    .Q(\atari2600.ram[90][0] ));
 sg13g2_dfrbp_1 _27780_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2695),
    .D(_00182_),
    .Q_N(_13822_),
    .Q(\atari2600.ram[90][1] ));
 sg13g2_dfrbp_1 _27781_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2694),
    .D(_00183_),
    .Q_N(_13821_),
    .Q(\atari2600.ram[90][2] ));
 sg13g2_dfrbp_1 _27782_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2693),
    .D(_00184_),
    .Q_N(_13820_),
    .Q(\atari2600.ram[90][3] ));
 sg13g2_dfrbp_1 _27783_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2692),
    .D(_00185_),
    .Q_N(_13819_),
    .Q(\atari2600.ram[90][4] ));
 sg13g2_dfrbp_1 _27784_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2691),
    .D(_00186_),
    .Q_N(_13818_),
    .Q(\atari2600.ram[90][5] ));
 sg13g2_dfrbp_1 _27785_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2690),
    .D(_00187_),
    .Q_N(_13817_),
    .Q(\atari2600.ram[90][6] ));
 sg13g2_dfrbp_1 _27786_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2689),
    .D(_00188_),
    .Q_N(_13816_),
    .Q(\atari2600.ram[90][7] ));
 sg13g2_dfrbp_1 _27787_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2688),
    .D(_00189_),
    .Q_N(_13815_),
    .Q(\atari2600.ram[2][0] ));
 sg13g2_dfrbp_1 _27788_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2687),
    .D(_00190_),
    .Q_N(_13814_),
    .Q(\atari2600.ram[2][1] ));
 sg13g2_dfrbp_1 _27789_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2686),
    .D(_00191_),
    .Q_N(_13813_),
    .Q(\atari2600.ram[2][2] ));
 sg13g2_dfrbp_1 _27790_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2685),
    .D(_00192_),
    .Q_N(_13812_),
    .Q(\atari2600.ram[2][3] ));
 sg13g2_dfrbp_1 _27791_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2684),
    .D(_00193_),
    .Q_N(_13811_),
    .Q(\atari2600.ram[2][4] ));
 sg13g2_dfrbp_1 _27792_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2683),
    .D(_00194_),
    .Q_N(_13810_),
    .Q(\atari2600.ram[2][5] ));
 sg13g2_dfrbp_1 _27793_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2682),
    .D(_00195_),
    .Q_N(_13809_),
    .Q(\atari2600.ram[2][6] ));
 sg13g2_dfrbp_1 _27794_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2681),
    .D(_00196_),
    .Q_N(_13808_),
    .Q(\atari2600.ram[2][7] ));
 sg13g2_dfrbp_1 _27795_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2680),
    .D(_00197_),
    .Q_N(_13807_),
    .Q(\atari2600.ram[94][0] ));
 sg13g2_dfrbp_1 _27796_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2679),
    .D(_00198_),
    .Q_N(_13806_),
    .Q(\atari2600.ram[94][1] ));
 sg13g2_dfrbp_1 _27797_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2678),
    .D(_00199_),
    .Q_N(_13805_),
    .Q(\atari2600.ram[94][2] ));
 sg13g2_dfrbp_1 _27798_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2677),
    .D(_00200_),
    .Q_N(_13804_),
    .Q(\atari2600.ram[94][3] ));
 sg13g2_dfrbp_1 _27799_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2676),
    .D(_00201_),
    .Q_N(_13803_),
    .Q(\atari2600.ram[94][4] ));
 sg13g2_dfrbp_1 _27800_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2675),
    .D(_00202_),
    .Q_N(_13802_),
    .Q(\atari2600.ram[94][5] ));
 sg13g2_dfrbp_1 _27801_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2674),
    .D(_00203_),
    .Q_N(_13801_),
    .Q(\atari2600.ram[94][6] ));
 sg13g2_dfrbp_1 _27802_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2673),
    .D(_00204_),
    .Q_N(_13800_),
    .Q(\atari2600.ram[94][7] ));
 sg13g2_dfrbp_1 _27803_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2672),
    .D(_00205_),
    .Q_N(_13799_),
    .Q(\atari2600.ram[76][0] ));
 sg13g2_dfrbp_1 _27804_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2671),
    .D(_00206_),
    .Q_N(_13798_),
    .Q(\atari2600.ram[76][1] ));
 sg13g2_dfrbp_1 _27805_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2670),
    .D(_00207_),
    .Q_N(_13797_),
    .Q(\atari2600.ram[76][2] ));
 sg13g2_dfrbp_1 _27806_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2669),
    .D(_00208_),
    .Q_N(_13796_),
    .Q(\atari2600.ram[76][3] ));
 sg13g2_dfrbp_1 _27807_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2668),
    .D(_00209_),
    .Q_N(_13795_),
    .Q(\atari2600.ram[76][4] ));
 sg13g2_dfrbp_1 _27808_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2667),
    .D(_00210_),
    .Q_N(_13794_),
    .Q(\atari2600.ram[76][5] ));
 sg13g2_dfrbp_1 _27809_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2666),
    .D(_00211_),
    .Q_N(_13793_),
    .Q(\atari2600.ram[76][6] ));
 sg13g2_dfrbp_1 _27810_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2665),
    .D(_00212_),
    .Q_N(_13792_),
    .Q(\atari2600.ram[76][7] ));
 sg13g2_dfrbp_1 _27811_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2664),
    .D(_00213_),
    .Q_N(_13791_),
    .Q(\atari2600.ram[93][0] ));
 sg13g2_dfrbp_1 _27812_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2663),
    .D(_00214_),
    .Q_N(_13790_),
    .Q(\atari2600.ram[93][1] ));
 sg13g2_dfrbp_1 _27813_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2662),
    .D(_00215_),
    .Q_N(_13789_),
    .Q(\atari2600.ram[93][2] ));
 sg13g2_dfrbp_1 _27814_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2661),
    .D(_00216_),
    .Q_N(_13788_),
    .Q(\atari2600.ram[93][3] ));
 sg13g2_dfrbp_1 _27815_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2660),
    .D(_00217_),
    .Q_N(_13787_),
    .Q(\atari2600.ram[93][4] ));
 sg13g2_dfrbp_1 _27816_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2659),
    .D(_00218_),
    .Q_N(_13786_),
    .Q(\atari2600.ram[93][5] ));
 sg13g2_dfrbp_1 _27817_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2658),
    .D(_00219_),
    .Q_N(_13785_),
    .Q(\atari2600.ram[93][6] ));
 sg13g2_dfrbp_1 _27818_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2657),
    .D(_00220_),
    .Q_N(_13784_),
    .Q(\atari2600.ram[93][7] ));
 sg13g2_dfrbp_1 _27819_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net2656),
    .D(_00221_),
    .Q_N(_13783_),
    .Q(\atari2600.ram[78][0] ));
 sg13g2_dfrbp_1 _27820_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2655),
    .D(_00222_),
    .Q_N(_13782_),
    .Q(\atari2600.ram[78][1] ));
 sg13g2_dfrbp_1 _27821_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2654),
    .D(_00223_),
    .Q_N(_13781_),
    .Q(\atari2600.ram[78][2] ));
 sg13g2_dfrbp_1 _27822_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2653),
    .D(_00224_),
    .Q_N(_13780_),
    .Q(\atari2600.ram[78][3] ));
 sg13g2_dfrbp_1 _27823_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2652),
    .D(_00225_),
    .Q_N(_13779_),
    .Q(\atari2600.ram[78][4] ));
 sg13g2_dfrbp_1 _27824_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net2651),
    .D(_00226_),
    .Q_N(_13778_),
    .Q(\atari2600.ram[78][5] ));
 sg13g2_dfrbp_1 _27825_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net2650),
    .D(_00227_),
    .Q_N(_13777_),
    .Q(\atari2600.ram[78][6] ));
 sg13g2_dfrbp_1 _27826_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net2649),
    .D(_00228_),
    .Q_N(_13776_),
    .Q(\atari2600.ram[78][7] ));
 sg13g2_dfrbp_1 _27827_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2648),
    .D(_00229_),
    .Q_N(_13775_),
    .Q(\atari2600.ram[71][0] ));
 sg13g2_dfrbp_1 _27828_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2647),
    .D(_00230_),
    .Q_N(_13774_),
    .Q(\atari2600.ram[71][1] ));
 sg13g2_dfrbp_1 _27829_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2646),
    .D(_00231_),
    .Q_N(_13773_),
    .Q(\atari2600.ram[71][2] ));
 sg13g2_dfrbp_1 _27830_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2645),
    .D(_00232_),
    .Q_N(_13772_),
    .Q(\atari2600.ram[71][3] ));
 sg13g2_dfrbp_1 _27831_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2644),
    .D(_00233_),
    .Q_N(_13771_),
    .Q(\atari2600.ram[71][4] ));
 sg13g2_dfrbp_1 _27832_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2643),
    .D(_00234_),
    .Q_N(_13770_),
    .Q(\atari2600.ram[71][5] ));
 sg13g2_dfrbp_1 _27833_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2642),
    .D(_00235_),
    .Q_N(_13769_),
    .Q(\atari2600.ram[71][6] ));
 sg13g2_dfrbp_1 _27834_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2641),
    .D(_00236_),
    .Q_N(_13768_),
    .Q(\atari2600.ram[71][7] ));
 sg13g2_dfrbp_1 _27835_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2640),
    .D(_00237_),
    .Q_N(_13767_),
    .Q(\scanline[9][0] ));
 sg13g2_dfrbp_1 _27836_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2639),
    .D(_00238_),
    .Q_N(_13766_),
    .Q(\scanline[9][1] ));
 sg13g2_dfrbp_1 _27837_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2638),
    .D(_00239_),
    .Q_N(_13765_),
    .Q(\scanline[9][2] ));
 sg13g2_dfrbp_1 _27838_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2637),
    .D(_00240_),
    .Q_N(_13764_),
    .Q(\scanline[9][3] ));
 sg13g2_dfrbp_1 _27839_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2636),
    .D(_00241_),
    .Q_N(_13763_),
    .Q(\scanline[9][4] ));
 sg13g2_dfrbp_1 _27840_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2635),
    .D(_00242_),
    .Q_N(_13762_),
    .Q(\scanline[9][5] ));
 sg13g2_dfrbp_1 _27841_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2634),
    .D(_00243_),
    .Q_N(_13761_),
    .Q(\scanline[9][6] ));
 sg13g2_dfrbp_1 _27842_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2633),
    .D(_00244_),
    .Q_N(_13760_),
    .Q(\atari2600.ram[22][0] ));
 sg13g2_dfrbp_1 _27843_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2632),
    .D(_00245_),
    .Q_N(_13759_),
    .Q(\atari2600.ram[22][1] ));
 sg13g2_dfrbp_1 _27844_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2631),
    .D(_00246_),
    .Q_N(_13758_),
    .Q(\atari2600.ram[22][2] ));
 sg13g2_dfrbp_1 _27845_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2630),
    .D(_00247_),
    .Q_N(_13757_),
    .Q(\atari2600.ram[22][3] ));
 sg13g2_dfrbp_1 _27846_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2629),
    .D(_00248_),
    .Q_N(_13756_),
    .Q(\atari2600.ram[22][4] ));
 sg13g2_dfrbp_1 _27847_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2628),
    .D(_00249_),
    .Q_N(_13755_),
    .Q(\atari2600.ram[22][5] ));
 sg13g2_dfrbp_1 _27848_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2627),
    .D(_00250_),
    .Q_N(_13754_),
    .Q(\atari2600.ram[22][6] ));
 sg13g2_dfrbp_1 _27849_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2626),
    .D(_00251_),
    .Q_N(_13753_),
    .Q(\atari2600.ram[22][7] ));
 sg13g2_dfrbp_1 _27850_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2625),
    .D(_00252_),
    .Q_N(_13752_),
    .Q(\atari2600.ram[26][0] ));
 sg13g2_dfrbp_1 _27851_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net2624),
    .D(_00253_),
    .Q_N(_13751_),
    .Q(\atari2600.ram[26][1] ));
 sg13g2_dfrbp_1 _27852_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2623),
    .D(_00254_),
    .Q_N(_13750_),
    .Q(\atari2600.ram[26][2] ));
 sg13g2_dfrbp_1 _27853_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2622),
    .D(_00255_),
    .Q_N(_13749_),
    .Q(\atari2600.ram[26][3] ));
 sg13g2_dfrbp_1 _27854_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2621),
    .D(_00256_),
    .Q_N(_13748_),
    .Q(\atari2600.ram[26][4] ));
 sg13g2_dfrbp_1 _27855_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2620),
    .D(_00257_),
    .Q_N(_13747_),
    .Q(\atari2600.ram[26][5] ));
 sg13g2_dfrbp_1 _27856_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2619),
    .D(_00258_),
    .Q_N(_13746_),
    .Q(\atari2600.ram[26][6] ));
 sg13g2_dfrbp_1 _27857_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2618),
    .D(_00259_),
    .Q_N(_13745_),
    .Q(\atari2600.ram[26][7] ));
 sg13g2_dfrbp_1 _27858_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2617),
    .D(_00260_),
    .Q_N(_13744_),
    .Q(spi_restart));
 sg13g2_dfrbp_1 _27859_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net99),
    .D(_00261_),
    .Q_N(_13828_),
    .Q(\flash_rom.stall_read ));
 sg13g2_dfrbp_1 _27860_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net188),
    .D(net2932),
    .Q_N(_13829_),
    .Q(spi_data_ready_last));
 sg13g2_dfrbp_1 _27861_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2616),
    .D(_00000_),
    .Q_N(_13743_),
    .Q(rom_data_pending));
 sg13g2_dfrbp_1 _27862_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2615),
    .D(_00262_),
    .Q_N(_00169_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _27863_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2614),
    .D(net7470),
    .Q_N(_13742_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _27864_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2613),
    .D(_00264_),
    .Q_N(_13741_),
    .Q(\rom_last_read_addr[0] ));
 sg13g2_dfrbp_1 _27865_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2612),
    .D(net7076),
    .Q_N(_13740_),
    .Q(\rom_last_read_addr[1] ));
 sg13g2_dfrbp_1 _27866_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2611),
    .D(net4510),
    .Q_N(_13739_),
    .Q(\rom_last_read_addr[2] ));
 sg13g2_dfrbp_1 _27867_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2610),
    .D(net4671),
    .Q_N(_13738_),
    .Q(\rom_last_read_addr[3] ));
 sg13g2_dfrbp_1 _27868_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2609),
    .D(net6627),
    .Q_N(_13737_),
    .Q(\rom_last_read_addr[4] ));
 sg13g2_dfrbp_1 _27869_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2608),
    .D(net4337),
    .Q_N(_13736_),
    .Q(\rom_last_read_addr[5] ));
 sg13g2_dfrbp_1 _27870_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2607),
    .D(net7247),
    .Q_N(_13735_),
    .Q(\rom_last_read_addr[6] ));
 sg13g2_dfrbp_1 _27871_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2606),
    .D(net7114),
    .Q_N(_13734_),
    .Q(\rom_last_read_addr[7] ));
 sg13g2_dfrbp_1 _27872_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2605),
    .D(net4920),
    .Q_N(_13733_),
    .Q(\rom_last_read_addr[8] ));
 sg13g2_dfrbp_1 _27873_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2604),
    .D(net7330),
    .Q_N(_13732_),
    .Q(\rom_last_read_addr[9] ));
 sg13g2_dfrbp_1 _27874_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2603),
    .D(net4371),
    .Q_N(_13731_),
    .Q(\rom_last_read_addr[10] ));
 sg13g2_dfrbp_1 _27875_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2602),
    .D(net6965),
    .Q_N(_13730_),
    .Q(\rom_last_read_addr[11] ));
 sg13g2_dfrbp_1 _27876_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2601),
    .D(_00276_),
    .Q_N(_13729_),
    .Q(\atari2600.ram[7][0] ));
 sg13g2_dfrbp_1 _27877_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2600),
    .D(_00277_),
    .Q_N(_13728_),
    .Q(\atari2600.ram[7][1] ));
 sg13g2_dfrbp_1 _27878_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2599),
    .D(_00278_),
    .Q_N(_13727_),
    .Q(\atari2600.ram[7][2] ));
 sg13g2_dfrbp_1 _27879_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2598),
    .D(_00279_),
    .Q_N(_13726_),
    .Q(\atari2600.ram[7][3] ));
 sg13g2_dfrbp_1 _27880_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2597),
    .D(_00280_),
    .Q_N(_13725_),
    .Q(\atari2600.ram[7][4] ));
 sg13g2_dfrbp_1 _27881_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2596),
    .D(_00281_),
    .Q_N(_13724_),
    .Q(\atari2600.ram[7][5] ));
 sg13g2_dfrbp_1 _27882_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2595),
    .D(_00282_),
    .Q_N(_13723_),
    .Q(\atari2600.ram[7][6] ));
 sg13g2_dfrbp_1 _27883_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2594),
    .D(_00283_),
    .Q_N(_13722_),
    .Q(\atari2600.ram[7][7] ));
 sg13g2_dfrbp_1 _27884_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2593),
    .D(net7166),
    .Q_N(_00093_),
    .Q(\rom_next_addr_in_queue[0] ));
 sg13g2_dfrbp_1 _27885_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2592),
    .D(net7224),
    .Q_N(_13721_),
    .Q(\rom_next_addr_in_queue[1] ));
 sg13g2_dfrbp_1 _27886_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2591),
    .D(_00286_),
    .Q_N(_13720_),
    .Q(\rom_next_addr_in_queue[2] ));
 sg13g2_dfrbp_1 _27887_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2590),
    .D(_00287_),
    .Q_N(_13719_),
    .Q(\rom_next_addr_in_queue[3] ));
 sg13g2_dfrbp_1 _27888_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2589),
    .D(_00288_),
    .Q_N(_13718_),
    .Q(\rom_next_addr_in_queue[4] ));
 sg13g2_dfrbp_1 _27889_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2588),
    .D(_00289_),
    .Q_N(_13717_),
    .Q(\rom_next_addr_in_queue[5] ));
 sg13g2_dfrbp_1 _27890_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2587),
    .D(_00290_),
    .Q_N(_13716_),
    .Q(\rom_next_addr_in_queue[6] ));
 sg13g2_dfrbp_1 _27891_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2586),
    .D(net7423),
    .Q_N(_13715_),
    .Q(\rom_next_addr_in_queue[7] ));
 sg13g2_dfrbp_1 _27892_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2585),
    .D(_00292_),
    .Q_N(_13714_),
    .Q(\rom_next_addr_in_queue[8] ));
 sg13g2_dfrbp_1 _27893_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2584),
    .D(_00293_),
    .Q_N(_13713_),
    .Q(\rom_next_addr_in_queue[9] ));
 sg13g2_dfrbp_1 _27894_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2583),
    .D(net7324),
    .Q_N(_13712_),
    .Q(\rom_next_addr_in_queue[10] ));
 sg13g2_dfrbp_1 _27895_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2582),
    .D(_00295_),
    .Q_N(_13711_),
    .Q(\rom_next_addr_in_queue[11] ));
 sg13g2_dfrbp_1 _27896_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2581),
    .D(net7375),
    .Q_N(_13710_),
    .Q(\audio_pwm_accumulator[0] ));
 sg13g2_dfrbp_1 _27897_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2580),
    .D(_00297_),
    .Q_N(_13709_),
    .Q(\audio_pwm_accumulator[1] ));
 sg13g2_dfrbp_1 _27898_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2579),
    .D(_00298_),
    .Q_N(_13708_),
    .Q(\audio_pwm_accumulator[2] ));
 sg13g2_dfrbp_1 _27899_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2578),
    .D(_00299_),
    .Q_N(_13707_),
    .Q(\audio_pwm_accumulator[3] ));
 sg13g2_dfrbp_1 _27900_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2577),
    .D(_00300_),
    .Q_N(_13706_),
    .Q(\audio_pwm_accumulator[4] ));
 sg13g2_dfrbp_1 _27901_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net2576),
    .D(_00301_),
    .Q_N(_13705_),
    .Q(audio_pwm));
 sg13g2_dfrbp_1 _27902_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2575),
    .D(_00302_),
    .Q_N(_13704_),
    .Q(\r_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27903_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2574),
    .D(_00303_),
    .Q_N(_13703_),
    .Q(\r_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27904_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2573),
    .D(_00304_),
    .Q_N(_13702_),
    .Q(\r_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27905_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2572),
    .D(_00305_),
    .Q_N(_13701_),
    .Q(\r_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27906_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2571),
    .D(_00306_),
    .Q_N(_13700_),
    .Q(\r_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27907_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2570),
    .D(_00307_),
    .Q_N(_13699_),
    .Q(\r_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27908_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2569),
    .D(_00308_),
    .Q_N(_13698_),
    .Q(\r_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27909_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2568),
    .D(_00309_),
    .Q_N(_13697_),
    .Q(\r_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27910_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2567),
    .D(_00310_),
    .Q_N(_13696_),
    .Q(\r_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27911_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2566),
    .D(_00311_),
    .Q_N(_13695_),
    .Q(\g_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27912_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2565),
    .D(_00312_),
    .Q_N(_13694_),
    .Q(\g_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27913_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2564),
    .D(_00313_),
    .Q_N(_00069_),
    .Q(\g_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27914_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2563),
    .D(_00314_),
    .Q_N(_13693_),
    .Q(\g_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27915_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2562),
    .D(_00315_),
    .Q_N(_13692_),
    .Q(\g_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27916_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2561),
    .D(_00316_),
    .Q_N(_13691_),
    .Q(\g_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27917_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2560),
    .D(_00317_),
    .Q_N(_13690_),
    .Q(\g_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27918_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2559),
    .D(_00318_),
    .Q_N(_13689_),
    .Q(\g_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27919_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2558),
    .D(_00319_),
    .Q_N(_13688_),
    .Q(\g_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27920_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2557),
    .D(_00320_),
    .Q_N(_13687_),
    .Q(\b_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27921_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2556),
    .D(_00321_),
    .Q_N(_13686_),
    .Q(\b_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27922_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2555),
    .D(_00322_),
    .Q_N(_13685_),
    .Q(\b_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27923_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2554),
    .D(_00323_),
    .Q_N(_13684_),
    .Q(\b_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27924_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2553),
    .D(_00324_),
    .Q_N(_13683_),
    .Q(\b_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27925_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2552),
    .D(_00325_),
    .Q_N(_13682_),
    .Q(\b_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27926_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2551),
    .D(_00326_),
    .Q_N(_13681_),
    .Q(\b_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27927_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2550),
    .D(_00327_),
    .Q_N(_13680_),
    .Q(\b_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27928_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2549),
    .D(_00328_),
    .Q_N(_13679_),
    .Q(\b_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27929_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2548),
    .D(_00329_),
    .Q_N(_13678_),
    .Q(\r_pwm_even[1] ));
 sg13g2_dfrbp_1 _27930_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2547),
    .D(net7359),
    .Q_N(_13677_),
    .Q(\r_pwm_even[2] ));
 sg13g2_dfrbp_1 _27931_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2546),
    .D(_00331_),
    .Q_N(_13676_),
    .Q(\r_pwm_even[3] ));
 sg13g2_dfrbp_1 _27932_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2545),
    .D(_00332_),
    .Q_N(_13675_),
    .Q(\r_pwm_even[4] ));
 sg13g2_dfrbp_1 _27933_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2544),
    .D(_00333_),
    .Q_N(_13674_),
    .Q(\r_pwm_even[5] ));
 sg13g2_dfrbp_1 _27934_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2543),
    .D(_00334_),
    .Q_N(_13673_),
    .Q(\r_pwm_even[6] ));
 sg13g2_dfrbp_1 _27935_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2542),
    .D(_00335_),
    .Q_N(_13672_),
    .Q(\r_pwm_even[7] ));
 sg13g2_dfrbp_1 _27936_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2541),
    .D(_00336_),
    .Q_N(_13671_),
    .Q(\r_pwm_even[8] ));
 sg13g2_dfrbp_1 _27937_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2540),
    .D(_00337_),
    .Q_N(_13670_),
    .Q(\r_pwm_even[9] ));
 sg13g2_dfrbp_1 _27938_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2539),
    .D(net4277),
    .Q_N(_13669_),
    .Q(\g_pwm_even[1] ));
 sg13g2_dfrbp_1 _27939_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2538),
    .D(_00339_),
    .Q_N(_13668_),
    .Q(\g_pwm_even[2] ));
 sg13g2_dfrbp_1 _27940_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2537),
    .D(_00340_),
    .Q_N(_13667_),
    .Q(\g_pwm_even[3] ));
 sg13g2_dfrbp_1 _27941_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2536),
    .D(_00341_),
    .Q_N(_13666_),
    .Q(\g_pwm_even[4] ));
 sg13g2_dfrbp_1 _27942_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2535),
    .D(_00342_),
    .Q_N(_13665_),
    .Q(\g_pwm_even[5] ));
 sg13g2_dfrbp_1 _27943_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2534),
    .D(_00343_),
    .Q_N(_13664_),
    .Q(\g_pwm_even[6] ));
 sg13g2_dfrbp_1 _27944_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2533),
    .D(_00344_),
    .Q_N(_13663_),
    .Q(\g_pwm_even[7] ));
 sg13g2_dfrbp_1 _27945_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2532),
    .D(_00345_),
    .Q_N(_13662_),
    .Q(\g_pwm_even[8] ));
 sg13g2_dfrbp_1 _27946_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2531),
    .D(_00346_),
    .Q_N(_13661_),
    .Q(\g_pwm_even[9] ));
 sg13g2_dfrbp_1 _27947_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2530),
    .D(net2934),
    .Q_N(_00167_),
    .Q(\frame_counter[0] ));
 sg13g2_dfrbp_1 _27948_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2529),
    .D(net4245),
    .Q_N(_13660_),
    .Q(\frame_counter[1] ));
 sg13g2_dfrbp_1 _27949_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net218),
    .D(_00349_),
    .Q_N(_13830_),
    .Q(\frame_counter[2] ));
 sg13g2_dfrbp_1 _27950_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2528),
    .D(net2931),
    .Q_N(_13659_),
    .Q(tia_vsync_last));
 sg13g2_dfrbp_1 _27951_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2527),
    .D(_00350_),
    .Q_N(_13658_),
    .Q(\atari2600.input_switches[0] ));
 sg13g2_dfrbp_1 _27952_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2526),
    .D(_00351_),
    .Q_N(_13657_),
    .Q(\atari2600.input_switches[1] ));
 sg13g2_dfrbp_1 _27953_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2525),
    .D(_00352_),
    .Q_N(_13656_),
    .Q(\atari2600.input_switches[2] ));
 sg13g2_dfrbp_1 _27954_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2524),
    .D(_00353_),
    .Q_N(_13655_),
    .Q(\atari2600.input_switches[3] ));
 sg13g2_dfrbp_1 _27955_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2523),
    .D(_00354_),
    .Q_N(_13654_),
    .Q(\b_pwm_even[1] ));
 sg13g2_dfrbp_1 _27956_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2522),
    .D(_00355_),
    .Q_N(_13653_),
    .Q(\b_pwm_even[2] ));
 sg13g2_dfrbp_1 _27957_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2521),
    .D(_00356_),
    .Q_N(_13652_),
    .Q(\b_pwm_even[3] ));
 sg13g2_dfrbp_1 _27958_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2520),
    .D(_00357_),
    .Q_N(_13651_),
    .Q(\b_pwm_even[4] ));
 sg13g2_dfrbp_1 _27959_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2519),
    .D(_00358_),
    .Q_N(_13650_),
    .Q(\b_pwm_even[5] ));
 sg13g2_dfrbp_1 _27960_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2518),
    .D(_00359_),
    .Q_N(_13649_),
    .Q(\b_pwm_even[6] ));
 sg13g2_dfrbp_1 _27961_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2517),
    .D(_00360_),
    .Q_N(_13648_),
    .Q(\b_pwm_even[7] ));
 sg13g2_dfrbp_1 _27962_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2516),
    .D(_00361_),
    .Q_N(_13647_),
    .Q(\b_pwm_even[8] ));
 sg13g2_dfrbp_1 _27963_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2515),
    .D(_00362_),
    .Q_N(_13646_),
    .Q(\b_pwm_even[9] ));
 sg13g2_dfrbp_1 _27964_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2514),
    .D(_00363_),
    .Q_N(_13645_),
    .Q(\atari2600.ram[73][0] ));
 sg13g2_dfrbp_1 _27965_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2513),
    .D(_00364_),
    .Q_N(_13644_),
    .Q(\atari2600.ram[73][1] ));
 sg13g2_dfrbp_1 _27966_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2512),
    .D(_00365_),
    .Q_N(_13643_),
    .Q(\atari2600.ram[73][2] ));
 sg13g2_dfrbp_1 _27967_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2511),
    .D(_00366_),
    .Q_N(_13642_),
    .Q(\atari2600.ram[73][3] ));
 sg13g2_dfrbp_1 _27968_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2510),
    .D(_00367_),
    .Q_N(_13641_),
    .Q(\atari2600.ram[73][4] ));
 sg13g2_dfrbp_1 _27969_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2509),
    .D(_00368_),
    .Q_N(_13640_),
    .Q(\atari2600.ram[73][5] ));
 sg13g2_dfrbp_1 _27970_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2508),
    .D(_00369_),
    .Q_N(_13639_),
    .Q(\atari2600.ram[73][6] ));
 sg13g2_dfrbp_1 _27971_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net2507),
    .D(_00370_),
    .Q_N(_13638_),
    .Q(\atari2600.ram[73][7] ));
 sg13g2_dfrbp_1 _27972_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2506),
    .D(_00371_),
    .Q_N(_13637_),
    .Q(\atari2600.ram[127][0] ));
 sg13g2_dfrbp_1 _27973_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net2505),
    .D(_00372_),
    .Q_N(_13636_),
    .Q(\atari2600.ram[127][1] ));
 sg13g2_dfrbp_1 _27974_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2504),
    .D(_00373_),
    .Q_N(_13635_),
    .Q(\atari2600.ram[127][2] ));
 sg13g2_dfrbp_1 _27975_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2503),
    .D(_00374_),
    .Q_N(_13634_),
    .Q(\atari2600.ram[127][3] ));
 sg13g2_dfrbp_1 _27976_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2502),
    .D(_00375_),
    .Q_N(_13633_),
    .Q(\atari2600.ram[127][4] ));
 sg13g2_dfrbp_1 _27977_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2501),
    .D(_00376_),
    .Q_N(_13632_),
    .Q(\atari2600.ram[127][5] ));
 sg13g2_dfrbp_1 _27978_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net2500),
    .D(_00377_),
    .Q_N(_13631_),
    .Q(\atari2600.ram[127][6] ));
 sg13g2_dfrbp_1 _27979_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net219),
    .D(_00378_),
    .Q_N(_13831_),
    .Q(\atari2600.ram[127][7] ));
 sg13g2_dfrbp_1 _27980_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net6543),
    .D(_00171_),
    .Q_N(_13832_),
    .Q(\atari2600.cpu.state[0] ));
 sg13g2_dfrbp_1 _27981_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net6543),
    .D(_00172_),
    .Q_N(_13833_),
    .Q(\atari2600.cpu.state[1] ));
 sg13g2_dfrbp_1 _27982_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net6543),
    .D(_00173_),
    .Q_N(_13630_),
    .Q(\atari2600.cpu.state[2] ));
 sg13g2_dfrbp_1 _27983_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net6543),
    .D(_00176_),
    .Q_N(\atari2600.cpu.state[3] ),
    .Q(_00170_));
 sg13g2_dfrbp_1 _27984_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net6543),
    .D(_00174_),
    .Q_N(_13834_),
    .Q(\atari2600.cpu.state[4] ));
 sg13g2_dfrbp_1 _27985_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net6545),
    .D(_00175_),
    .Q_N(_13629_),
    .Q(\atari2600.cpu.state[5] ));
 sg13g2_dfrbp_1 _27986_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2499),
    .D(_00379_),
    .Q_N(_13628_),
    .Q(\atari2600.ram[87][0] ));
 sg13g2_dfrbp_1 _27987_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2498),
    .D(_00380_),
    .Q_N(_13627_),
    .Q(\atari2600.ram[87][1] ));
 sg13g2_dfrbp_1 _27988_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2497),
    .D(_00381_),
    .Q_N(_13626_),
    .Q(\atari2600.ram[87][2] ));
 sg13g2_dfrbp_1 _27989_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2496),
    .D(_00382_),
    .Q_N(_13625_),
    .Q(\atari2600.ram[87][3] ));
 sg13g2_dfrbp_1 _27990_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2495),
    .D(_00383_),
    .Q_N(_13624_),
    .Q(\atari2600.ram[87][4] ));
 sg13g2_dfrbp_1 _27991_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2494),
    .D(_00384_),
    .Q_N(_13623_),
    .Q(\atari2600.ram[87][5] ));
 sg13g2_dfrbp_1 _27992_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2493),
    .D(_00385_),
    .Q_N(_13622_),
    .Q(\atari2600.ram[87][6] ));
 sg13g2_dfrbp_1 _27993_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2492),
    .D(_00386_),
    .Q_N(_13621_),
    .Q(\atari2600.ram[87][7] ));
 sg13g2_dfrbp_1 _27994_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2491),
    .D(_00387_),
    .Q_N(_13620_),
    .Q(\atari2600.ram[83][0] ));
 sg13g2_dfrbp_1 _27995_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2490),
    .D(_00388_),
    .Q_N(_13619_),
    .Q(\atari2600.ram[83][1] ));
 sg13g2_dfrbp_1 _27996_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2489),
    .D(_00389_),
    .Q_N(_13618_),
    .Q(\atari2600.ram[83][2] ));
 sg13g2_dfrbp_1 _27997_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2488),
    .D(_00390_),
    .Q_N(_13617_),
    .Q(\atari2600.ram[83][3] ));
 sg13g2_dfrbp_1 _27998_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2487),
    .D(_00391_),
    .Q_N(_13616_),
    .Q(\atari2600.ram[83][4] ));
 sg13g2_dfrbp_1 _27999_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2486),
    .D(_00392_),
    .Q_N(_13615_),
    .Q(\atari2600.ram[83][5] ));
 sg13g2_dfrbp_1 _28000_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2485),
    .D(_00393_),
    .Q_N(_13614_),
    .Q(\atari2600.ram[83][6] ));
 sg13g2_dfrbp_1 _28001_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2484),
    .D(_00394_),
    .Q_N(_13613_),
    .Q(\atari2600.ram[83][7] ));
 sg13g2_dfrbp_1 _28002_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2483),
    .D(_00395_),
    .Q_N(_13612_),
    .Q(\atari2600.ram[84][0] ));
 sg13g2_dfrbp_1 _28003_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2482),
    .D(_00396_),
    .Q_N(_13611_),
    .Q(\atari2600.ram[84][1] ));
 sg13g2_dfrbp_1 _28004_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2481),
    .D(_00397_),
    .Q_N(_13610_),
    .Q(\atari2600.ram[84][2] ));
 sg13g2_dfrbp_1 _28005_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2480),
    .D(_00398_),
    .Q_N(_13609_),
    .Q(\atari2600.ram[84][3] ));
 sg13g2_dfrbp_1 _28006_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2479),
    .D(_00399_),
    .Q_N(_13608_),
    .Q(\atari2600.ram[84][4] ));
 sg13g2_dfrbp_1 _28007_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2478),
    .D(_00400_),
    .Q_N(_13607_),
    .Q(\atari2600.ram[84][5] ));
 sg13g2_dfrbp_1 _28008_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2477),
    .D(_00401_),
    .Q_N(_13606_),
    .Q(\atari2600.ram[84][6] ));
 sg13g2_dfrbp_1 _28009_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2476),
    .D(_00402_),
    .Q_N(_13605_),
    .Q(\atari2600.ram[84][7] ));
 sg13g2_dfrbp_1 _28010_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2475),
    .D(_00403_),
    .Q_N(_13604_),
    .Q(\atari2600.ram[80][0] ));
 sg13g2_dfrbp_1 _28011_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2474),
    .D(_00404_),
    .Q_N(_13603_),
    .Q(\atari2600.ram[80][1] ));
 sg13g2_dfrbp_1 _28012_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2473),
    .D(_00405_),
    .Q_N(_13602_),
    .Q(\atari2600.ram[80][2] ));
 sg13g2_dfrbp_1 _28013_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2472),
    .D(_00406_),
    .Q_N(_13601_),
    .Q(\atari2600.ram[80][3] ));
 sg13g2_dfrbp_1 _28014_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2471),
    .D(_00407_),
    .Q_N(_13600_),
    .Q(\atari2600.ram[80][4] ));
 sg13g2_dfrbp_1 _28015_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2470),
    .D(_00408_),
    .Q_N(_13599_),
    .Q(\atari2600.ram[80][5] ));
 sg13g2_dfrbp_1 _28016_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2469),
    .D(_00409_),
    .Q_N(_13598_),
    .Q(\atari2600.ram[80][6] ));
 sg13g2_dfrbp_1 _28017_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2468),
    .D(_00410_),
    .Q_N(_13597_),
    .Q(\atari2600.ram[80][7] ));
 sg13g2_dfrbp_1 _28018_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2467),
    .D(_00411_),
    .Q_N(_13596_),
    .Q(\atari2600.ram[85][0] ));
 sg13g2_dfrbp_1 _28019_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2466),
    .D(_00412_),
    .Q_N(_13595_),
    .Q(\atari2600.ram[85][1] ));
 sg13g2_dfrbp_1 _28020_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2465),
    .D(_00413_),
    .Q_N(_13594_),
    .Q(\atari2600.ram[85][2] ));
 sg13g2_dfrbp_1 _28021_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2464),
    .D(_00414_),
    .Q_N(_13593_),
    .Q(\atari2600.ram[85][3] ));
 sg13g2_dfrbp_1 _28022_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2463),
    .D(_00415_),
    .Q_N(_13592_),
    .Q(\atari2600.ram[85][4] ));
 sg13g2_dfrbp_1 _28023_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2462),
    .D(_00416_),
    .Q_N(_13591_),
    .Q(\atari2600.ram[85][5] ));
 sg13g2_dfrbp_1 _28024_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2461),
    .D(_00417_),
    .Q_N(_13590_),
    .Q(\atari2600.ram[85][6] ));
 sg13g2_dfrbp_1 _28025_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2460),
    .D(_00418_),
    .Q_N(_13589_),
    .Q(\atari2600.ram[85][7] ));
 sg13g2_dfrbp_1 _28026_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2459),
    .D(_00419_),
    .Q_N(_13588_),
    .Q(\atari2600.ram[81][0] ));
 sg13g2_dfrbp_1 _28027_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2458),
    .D(_00420_),
    .Q_N(_13587_),
    .Q(\atari2600.ram[81][1] ));
 sg13g2_dfrbp_1 _28028_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2457),
    .D(_00421_),
    .Q_N(_13586_),
    .Q(\atari2600.ram[81][2] ));
 sg13g2_dfrbp_1 _28029_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2456),
    .D(_00422_),
    .Q_N(_13585_),
    .Q(\atari2600.ram[81][3] ));
 sg13g2_dfrbp_1 _28030_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2455),
    .D(_00423_),
    .Q_N(_13584_),
    .Q(\atari2600.ram[81][4] ));
 sg13g2_dfrbp_1 _28031_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2454),
    .D(_00424_),
    .Q_N(_13583_),
    .Q(\atari2600.ram[81][5] ));
 sg13g2_dfrbp_1 _28032_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2453),
    .D(_00425_),
    .Q_N(_13582_),
    .Q(\atari2600.ram[81][6] ));
 sg13g2_dfrbp_1 _28033_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2452),
    .D(_00426_),
    .Q_N(_13581_),
    .Q(\atari2600.ram[81][7] ));
 sg13g2_dfrbp_1 _28034_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2451),
    .D(_00427_),
    .Q_N(_13580_),
    .Q(\atari2600.ram[86][0] ));
 sg13g2_dfrbp_1 _28035_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2450),
    .D(_00428_),
    .Q_N(_13579_),
    .Q(\atari2600.ram[86][1] ));
 sg13g2_dfrbp_1 _28036_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2449),
    .D(_00429_),
    .Q_N(_13578_),
    .Q(\atari2600.ram[86][2] ));
 sg13g2_dfrbp_1 _28037_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2448),
    .D(_00430_),
    .Q_N(_13577_),
    .Q(\atari2600.ram[86][3] ));
 sg13g2_dfrbp_1 _28038_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2447),
    .D(_00431_),
    .Q_N(_13576_),
    .Q(\atari2600.ram[86][4] ));
 sg13g2_dfrbp_1 _28039_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2446),
    .D(_00432_),
    .Q_N(_13575_),
    .Q(\atari2600.ram[86][5] ));
 sg13g2_dfrbp_1 _28040_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2445),
    .D(_00433_),
    .Q_N(_13574_),
    .Q(\atari2600.ram[86][6] ));
 sg13g2_dfrbp_1 _28041_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2444),
    .D(_00434_),
    .Q_N(_13573_),
    .Q(\atari2600.ram[86][7] ));
 sg13g2_dfrbp_1 _28042_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2443),
    .D(_00435_),
    .Q_N(_13572_),
    .Q(\atari2600.ram[82][0] ));
 sg13g2_dfrbp_1 _28043_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2442),
    .D(_00436_),
    .Q_N(_13571_),
    .Q(\atari2600.ram[82][1] ));
 sg13g2_dfrbp_1 _28044_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2441),
    .D(_00437_),
    .Q_N(_13570_),
    .Q(\atari2600.ram[82][2] ));
 sg13g2_dfrbp_1 _28045_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2440),
    .D(_00438_),
    .Q_N(_13569_),
    .Q(\atari2600.ram[82][3] ));
 sg13g2_dfrbp_1 _28046_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2439),
    .D(_00439_),
    .Q_N(_13568_),
    .Q(\atari2600.ram[82][4] ));
 sg13g2_dfrbp_1 _28047_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2438),
    .D(_00440_),
    .Q_N(_13567_),
    .Q(\atari2600.ram[82][5] ));
 sg13g2_dfrbp_1 _28048_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2437),
    .D(_00441_),
    .Q_N(_13566_),
    .Q(\atari2600.ram[82][6] ));
 sg13g2_dfrbp_1 _28049_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2436),
    .D(_00442_),
    .Q_N(_13565_),
    .Q(\atari2600.ram[82][7] ));
 sg13g2_dfrbp_1 _28050_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2435),
    .D(_00443_),
    .Q_N(_13564_),
    .Q(\atari2600.ram[12][0] ));
 sg13g2_dfrbp_1 _28051_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2434),
    .D(_00444_),
    .Q_N(_13563_),
    .Q(\atari2600.ram[12][1] ));
 sg13g2_dfrbp_1 _28052_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2433),
    .D(_00445_),
    .Q_N(_13562_),
    .Q(\atari2600.ram[12][2] ));
 sg13g2_dfrbp_1 _28053_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2432),
    .D(_00446_),
    .Q_N(_13561_),
    .Q(\atari2600.ram[12][3] ));
 sg13g2_dfrbp_1 _28054_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2431),
    .D(_00447_),
    .Q_N(_13560_),
    .Q(\atari2600.ram[12][4] ));
 sg13g2_dfrbp_1 _28055_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2430),
    .D(_00448_),
    .Q_N(_13559_),
    .Q(\atari2600.ram[12][5] ));
 sg13g2_dfrbp_1 _28056_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2429),
    .D(_00449_),
    .Q_N(_13558_),
    .Q(\atari2600.ram[12][6] ));
 sg13g2_dfrbp_1 _28057_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2428),
    .D(_00450_),
    .Q_N(_13557_),
    .Q(\atari2600.ram[12][7] ));
 sg13g2_dfrbp_1 _28058_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net2427),
    .D(_00451_),
    .Q_N(_13556_),
    .Q(\atari2600.ram[77][0] ));
 sg13g2_dfrbp_1 _28059_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net2426),
    .D(_00452_),
    .Q_N(_13555_),
    .Q(\atari2600.ram[77][1] ));
 sg13g2_dfrbp_1 _28060_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2425),
    .D(_00453_),
    .Q_N(_13554_),
    .Q(\atari2600.ram[77][2] ));
 sg13g2_dfrbp_1 _28061_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2424),
    .D(_00454_),
    .Q_N(_13553_),
    .Q(\atari2600.ram[77][3] ));
 sg13g2_dfrbp_1 _28062_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2423),
    .D(_00455_),
    .Q_N(_13552_),
    .Q(\atari2600.ram[77][4] ));
 sg13g2_dfrbp_1 _28063_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2422),
    .D(_00456_),
    .Q_N(_13551_),
    .Q(\atari2600.ram[77][5] ));
 sg13g2_dfrbp_1 _28064_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2421),
    .D(_00457_),
    .Q_N(_13550_),
    .Q(\atari2600.ram[77][6] ));
 sg13g2_dfrbp_1 _28065_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net301),
    .D(_00458_),
    .Q_N(_13835_),
    .Q(\atari2600.ram[77][7] ));
 sg13g2_dfrbp_1 _28066_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net302),
    .D(_00009_),
    .Q_N(_13836_),
    .Q(\internal_rom_data[0] ));
 sg13g2_dfrbp_1 _28067_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net303),
    .D(_00010_),
    .Q_N(_13837_),
    .Q(\internal_rom_data[1] ));
 sg13g2_dfrbp_1 _28068_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net304),
    .D(_00011_),
    .Q_N(_13838_),
    .Q(\internal_rom_data[2] ));
 sg13g2_dfrbp_1 _28069_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net305),
    .D(_00012_),
    .Q_N(_13839_),
    .Q(\internal_rom_data[3] ));
 sg13g2_dfrbp_1 _28070_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net306),
    .D(_00013_),
    .Q_N(_13840_),
    .Q(\internal_rom_data[4] ));
 sg13g2_dfrbp_1 _28071_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net307),
    .D(_00014_),
    .Q_N(_13841_),
    .Q(\internal_rom_data[5] ));
 sg13g2_dfrbp_1 _28072_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net805),
    .D(_00015_),
    .Q_N(_13842_),
    .Q(\internal_rom_data[6] ));
 sg13g2_dfrbp_1 _28073_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2420),
    .D(_00016_),
    .Q_N(_13549_),
    .Q(\internal_rom_data[7] ));
 sg13g2_dfrbp_1 _28074_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2419),
    .D(_00459_),
    .Q_N(_13548_),
    .Q(\atari2600.cpu.ABH[0] ));
 sg13g2_dfrbp_1 _28075_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2418),
    .D(_00460_),
    .Q_N(_13547_),
    .Q(\atari2600.cpu.ABH[1] ));
 sg13g2_dfrbp_1 _28076_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2417),
    .D(_00461_),
    .Q_N(_13546_),
    .Q(\atari2600.cpu.ABH[2] ));
 sg13g2_dfrbp_1 _28077_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net2416),
    .D(_00462_),
    .Q_N(_13545_),
    .Q(\atari2600.cpu.ABH[3] ));
 sg13g2_dfrbp_1 _28078_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2415),
    .D(_00463_),
    .Q_N(_13544_),
    .Q(\atari2600.cpu.ABH[4] ));
 sg13g2_dfrbp_1 _28079_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2414),
    .D(_00464_),
    .Q_N(_13543_),
    .Q(\atari2600.ram[95][0] ));
 sg13g2_dfrbp_1 _28080_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2413),
    .D(_00465_),
    .Q_N(_13542_),
    .Q(\atari2600.ram[95][1] ));
 sg13g2_dfrbp_1 _28081_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2412),
    .D(_00466_),
    .Q_N(_13541_),
    .Q(\atari2600.ram[95][2] ));
 sg13g2_dfrbp_1 _28082_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2411),
    .D(_00467_),
    .Q_N(_13540_),
    .Q(\atari2600.ram[95][3] ));
 sg13g2_dfrbp_1 _28083_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2410),
    .D(_00468_),
    .Q_N(_13539_),
    .Q(\atari2600.ram[95][4] ));
 sg13g2_dfrbp_1 _28084_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2409),
    .D(_00469_),
    .Q_N(_13538_),
    .Q(\atari2600.ram[95][5] ));
 sg13g2_dfrbp_1 _28085_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2408),
    .D(_00470_),
    .Q_N(_13537_),
    .Q(\atari2600.ram[95][6] ));
 sg13g2_dfrbp_1 _28086_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2407),
    .D(_00471_),
    .Q_N(_13536_),
    .Q(\atari2600.ram[95][7] ));
 sg13g2_dfrbp_1 _28087_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2406),
    .D(_00472_),
    .Q_N(_13535_),
    .Q(\atari2600.ram[13][0] ));
 sg13g2_dfrbp_1 _28088_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2405),
    .D(_00473_),
    .Q_N(_13534_),
    .Q(\atari2600.ram[13][1] ));
 sg13g2_dfrbp_1 _28089_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2404),
    .D(_00474_),
    .Q_N(_13533_),
    .Q(\atari2600.ram[13][2] ));
 sg13g2_dfrbp_1 _28090_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2403),
    .D(_00475_),
    .Q_N(_13532_),
    .Q(\atari2600.ram[13][3] ));
 sg13g2_dfrbp_1 _28091_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2402),
    .D(_00476_),
    .Q_N(_13531_),
    .Q(\atari2600.ram[13][4] ));
 sg13g2_dfrbp_1 _28092_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2401),
    .D(_00477_),
    .Q_N(_13530_),
    .Q(\atari2600.ram[13][5] ));
 sg13g2_dfrbp_1 _28093_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2400),
    .D(_00478_),
    .Q_N(_13529_),
    .Q(\atari2600.ram[13][6] ));
 sg13g2_dfrbp_1 _28094_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2399),
    .D(_00479_),
    .Q_N(_13528_),
    .Q(\atari2600.ram[13][7] ));
 sg13g2_dfrbp_1 _28095_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2398),
    .D(_00480_),
    .Q_N(_13527_),
    .Q(\atari2600.ram[96][0] ));
 sg13g2_dfrbp_1 _28096_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2397),
    .D(_00481_),
    .Q_N(_13526_),
    .Q(\atari2600.ram[96][1] ));
 sg13g2_dfrbp_1 _28097_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2396),
    .D(_00482_),
    .Q_N(_13525_),
    .Q(\atari2600.ram[96][2] ));
 sg13g2_dfrbp_1 _28098_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2395),
    .D(_00483_),
    .Q_N(_13524_),
    .Q(\atari2600.ram[96][3] ));
 sg13g2_dfrbp_1 _28099_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2394),
    .D(_00484_),
    .Q_N(_13523_),
    .Q(\atari2600.ram[96][4] ));
 sg13g2_dfrbp_1 _28100_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2393),
    .D(_00485_),
    .Q_N(_13522_),
    .Q(\atari2600.ram[96][5] ));
 sg13g2_dfrbp_1 _28101_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2392),
    .D(_00486_),
    .Q_N(_13521_),
    .Q(\atari2600.ram[96][6] ));
 sg13g2_dfrbp_1 _28102_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2391),
    .D(_00487_),
    .Q_N(_13520_),
    .Q(\atari2600.ram[96][7] ));
 sg13g2_dfrbp_1 _28103_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2390),
    .D(_00488_),
    .Q_N(_13519_),
    .Q(\atari2600.ram[97][0] ));
 sg13g2_dfrbp_1 _28104_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2389),
    .D(_00489_),
    .Q_N(_13518_),
    .Q(\atari2600.ram[97][1] ));
 sg13g2_dfrbp_1 _28105_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2388),
    .D(_00490_),
    .Q_N(_13517_),
    .Q(\atari2600.ram[97][2] ));
 sg13g2_dfrbp_1 _28106_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2387),
    .D(_00491_),
    .Q_N(_13516_),
    .Q(\atari2600.ram[97][3] ));
 sg13g2_dfrbp_1 _28107_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2386),
    .D(_00492_),
    .Q_N(_13515_),
    .Q(\atari2600.ram[97][4] ));
 sg13g2_dfrbp_1 _28108_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2385),
    .D(_00493_),
    .Q_N(_13514_),
    .Q(\atari2600.ram[97][5] ));
 sg13g2_dfrbp_1 _28109_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2384),
    .D(_00494_),
    .Q_N(_13513_),
    .Q(\atari2600.ram[97][6] ));
 sg13g2_dfrbp_1 _28110_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2383),
    .D(_00495_),
    .Q_N(_13512_),
    .Q(\atari2600.ram[97][7] ));
 sg13g2_dfrbp_1 _28111_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2382),
    .D(_00496_),
    .Q_N(_13511_),
    .Q(\atari2600.ram[98][0] ));
 sg13g2_dfrbp_1 _28112_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2381),
    .D(_00497_),
    .Q_N(_13510_),
    .Q(\atari2600.ram[98][1] ));
 sg13g2_dfrbp_1 _28113_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2380),
    .D(_00498_),
    .Q_N(_13509_),
    .Q(\atari2600.ram[98][2] ));
 sg13g2_dfrbp_1 _28114_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2379),
    .D(_00499_),
    .Q_N(_13508_),
    .Q(\atari2600.ram[98][3] ));
 sg13g2_dfrbp_1 _28115_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2378),
    .D(_00500_),
    .Q_N(_13507_),
    .Q(\atari2600.ram[98][4] ));
 sg13g2_dfrbp_1 _28116_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2377),
    .D(_00501_),
    .Q_N(_13506_),
    .Q(\atari2600.ram[98][5] ));
 sg13g2_dfrbp_1 _28117_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2376),
    .D(_00502_),
    .Q_N(_13505_),
    .Q(\atari2600.ram[98][6] ));
 sg13g2_dfrbp_1 _28118_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2375),
    .D(_00503_),
    .Q_N(_13504_),
    .Q(\atari2600.ram[98][7] ));
 sg13g2_dfrbp_1 _28119_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2374),
    .D(_00504_),
    .Q_N(_13503_),
    .Q(\atari2600.ram[0][0] ));
 sg13g2_dfrbp_1 _28120_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2373),
    .D(_00505_),
    .Q_N(_13502_),
    .Q(\atari2600.ram[0][1] ));
 sg13g2_dfrbp_1 _28121_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2372),
    .D(_00506_),
    .Q_N(_13501_),
    .Q(\atari2600.ram[0][2] ));
 sg13g2_dfrbp_1 _28122_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2371),
    .D(_00507_),
    .Q_N(_13500_),
    .Q(\atari2600.ram[0][3] ));
 sg13g2_dfrbp_1 _28123_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2370),
    .D(_00508_),
    .Q_N(_13499_),
    .Q(\atari2600.ram[0][4] ));
 sg13g2_dfrbp_1 _28124_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2369),
    .D(_00509_),
    .Q_N(_13498_),
    .Q(\atari2600.ram[0][5] ));
 sg13g2_dfrbp_1 _28125_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net2368),
    .D(_00510_),
    .Q_N(_13497_),
    .Q(\atari2600.ram[0][6] ));
 sg13g2_dfrbp_1 _28126_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net2367),
    .D(_00511_),
    .Q_N(_13496_),
    .Q(\atari2600.ram[0][7] ));
 sg13g2_dfrbp_1 _28127_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2366),
    .D(_00512_),
    .Q_N(_13495_),
    .Q(\atari2600.ram[100][0] ));
 sg13g2_dfrbp_1 _28128_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2365),
    .D(_00513_),
    .Q_N(_13494_),
    .Q(\atari2600.ram[100][1] ));
 sg13g2_dfrbp_1 _28129_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2364),
    .D(_00514_),
    .Q_N(_13493_),
    .Q(\atari2600.ram[100][2] ));
 sg13g2_dfrbp_1 _28130_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2363),
    .D(_00515_),
    .Q_N(_13492_),
    .Q(\atari2600.ram[100][3] ));
 sg13g2_dfrbp_1 _28131_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2362),
    .D(_00516_),
    .Q_N(_13491_),
    .Q(\atari2600.ram[100][4] ));
 sg13g2_dfrbp_1 _28132_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2361),
    .D(_00517_),
    .Q_N(_13490_),
    .Q(\atari2600.ram[100][5] ));
 sg13g2_dfrbp_1 _28133_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2360),
    .D(_00518_),
    .Q_N(_13489_),
    .Q(\atari2600.ram[100][6] ));
 sg13g2_dfrbp_1 _28134_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2359),
    .D(_00519_),
    .Q_N(_13488_),
    .Q(\atari2600.ram[100][7] ));
 sg13g2_dfrbp_1 _28135_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2358),
    .D(_00520_),
    .Q_N(_13487_),
    .Q(\atari2600.ram[101][0] ));
 sg13g2_dfrbp_1 _28136_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2357),
    .D(_00521_),
    .Q_N(_13486_),
    .Q(\atari2600.ram[101][1] ));
 sg13g2_dfrbp_1 _28137_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2356),
    .D(_00522_),
    .Q_N(_13485_),
    .Q(\atari2600.ram[101][2] ));
 sg13g2_dfrbp_1 _28138_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2355),
    .D(_00523_),
    .Q_N(_13484_),
    .Q(\atari2600.ram[101][3] ));
 sg13g2_dfrbp_1 _28139_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2354),
    .D(_00524_),
    .Q_N(_13483_),
    .Q(\atari2600.ram[101][4] ));
 sg13g2_dfrbp_1 _28140_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2353),
    .D(_00525_),
    .Q_N(_13482_),
    .Q(\atari2600.ram[101][5] ));
 sg13g2_dfrbp_1 _28141_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2352),
    .D(_00526_),
    .Q_N(_13481_),
    .Q(\atari2600.ram[101][6] ));
 sg13g2_dfrbp_1 _28142_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2351),
    .D(_00527_),
    .Q_N(_13480_),
    .Q(\atari2600.ram[101][7] ));
 sg13g2_dfrbp_1 _28143_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2350),
    .D(_00528_),
    .Q_N(_13479_),
    .Q(\atari2600.ram[102][0] ));
 sg13g2_dfrbp_1 _28144_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2349),
    .D(_00529_),
    .Q_N(_13478_),
    .Q(\atari2600.ram[102][1] ));
 sg13g2_dfrbp_1 _28145_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2348),
    .D(_00530_),
    .Q_N(_13477_),
    .Q(\atari2600.ram[102][2] ));
 sg13g2_dfrbp_1 _28146_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2347),
    .D(_00531_),
    .Q_N(_13476_),
    .Q(\atari2600.ram[102][3] ));
 sg13g2_dfrbp_1 _28147_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2346),
    .D(_00532_),
    .Q_N(_13475_),
    .Q(\atari2600.ram[102][4] ));
 sg13g2_dfrbp_1 _28148_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2345),
    .D(_00533_),
    .Q_N(_13474_),
    .Q(\atari2600.ram[102][5] ));
 sg13g2_dfrbp_1 _28149_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net2344),
    .D(_00534_),
    .Q_N(_13473_),
    .Q(\atari2600.ram[102][6] ));
 sg13g2_dfrbp_1 _28150_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2343),
    .D(_00535_),
    .Q_N(_13472_),
    .Q(\atari2600.ram[102][7] ));
 sg13g2_dfrbp_1 _28151_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2342),
    .D(_00536_),
    .Q_N(_13471_),
    .Q(\atari2600.ram[103][0] ));
 sg13g2_dfrbp_1 _28152_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2341),
    .D(_00537_),
    .Q_N(_13470_),
    .Q(\atari2600.ram[103][1] ));
 sg13g2_dfrbp_1 _28153_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2340),
    .D(_00538_),
    .Q_N(_13469_),
    .Q(\atari2600.ram[103][2] ));
 sg13g2_dfrbp_1 _28154_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2339),
    .D(_00539_),
    .Q_N(_13468_),
    .Q(\atari2600.ram[103][3] ));
 sg13g2_dfrbp_1 _28155_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2338),
    .D(_00540_),
    .Q_N(_13467_),
    .Q(\atari2600.ram[103][4] ));
 sg13g2_dfrbp_1 _28156_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2337),
    .D(_00541_),
    .Q_N(_13466_),
    .Q(\atari2600.ram[103][5] ));
 sg13g2_dfrbp_1 _28157_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2336),
    .D(_00542_),
    .Q_N(_13465_),
    .Q(\atari2600.ram[103][6] ));
 sg13g2_dfrbp_1 _28158_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2335),
    .D(_00543_),
    .Q_N(_13464_),
    .Q(\atari2600.ram[103][7] ));
 sg13g2_dfrbp_1 _28159_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2334),
    .D(_00544_),
    .Q_N(_13463_),
    .Q(\atari2600.ram[104][0] ));
 sg13g2_dfrbp_1 _28160_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2333),
    .D(_00545_),
    .Q_N(_13462_),
    .Q(\atari2600.ram[104][1] ));
 sg13g2_dfrbp_1 _28161_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2332),
    .D(_00546_),
    .Q_N(_13461_),
    .Q(\atari2600.ram[104][2] ));
 sg13g2_dfrbp_1 _28162_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2331),
    .D(_00547_),
    .Q_N(_13460_),
    .Q(\atari2600.ram[104][3] ));
 sg13g2_dfrbp_1 _28163_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2330),
    .D(_00548_),
    .Q_N(_13459_),
    .Q(\atari2600.ram[104][4] ));
 sg13g2_dfrbp_1 _28164_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2329),
    .D(_00549_),
    .Q_N(_13458_),
    .Q(\atari2600.ram[104][5] ));
 sg13g2_dfrbp_1 _28165_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2328),
    .D(_00550_),
    .Q_N(_13457_),
    .Q(\atari2600.ram[104][6] ));
 sg13g2_dfrbp_1 _28166_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2327),
    .D(_00551_),
    .Q_N(_13456_),
    .Q(\atari2600.ram[104][7] ));
 sg13g2_dfrbp_1 _28167_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2326),
    .D(_00552_),
    .Q_N(_13455_),
    .Q(\atari2600.ram[105][0] ));
 sg13g2_dfrbp_1 _28168_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2325),
    .D(_00553_),
    .Q_N(_13454_),
    .Q(\atari2600.ram[105][1] ));
 sg13g2_dfrbp_1 _28169_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2324),
    .D(_00554_),
    .Q_N(_13453_),
    .Q(\atari2600.ram[105][2] ));
 sg13g2_dfrbp_1 _28170_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2323),
    .D(_00555_),
    .Q_N(_13452_),
    .Q(\atari2600.ram[105][3] ));
 sg13g2_dfrbp_1 _28171_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net2322),
    .D(_00556_),
    .Q_N(_13451_),
    .Q(\atari2600.ram[105][4] ));
 sg13g2_dfrbp_1 _28172_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2321),
    .D(_00557_),
    .Q_N(_13450_),
    .Q(\atari2600.ram[105][5] ));
 sg13g2_dfrbp_1 _28173_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2320),
    .D(_00558_),
    .Q_N(_13449_),
    .Q(\atari2600.ram[105][6] ));
 sg13g2_dfrbp_1 _28174_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2319),
    .D(_00559_),
    .Q_N(_13448_),
    .Q(\atari2600.ram[105][7] ));
 sg13g2_dfrbp_1 _28175_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2318),
    .D(_00560_),
    .Q_N(_13447_),
    .Q(\atari2600.ram[106][0] ));
 sg13g2_dfrbp_1 _28176_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2317),
    .D(_00561_),
    .Q_N(_13446_),
    .Q(\atari2600.ram[106][1] ));
 sg13g2_dfrbp_1 _28177_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2316),
    .D(_00562_),
    .Q_N(_13445_),
    .Q(\atari2600.ram[106][2] ));
 sg13g2_dfrbp_1 _28178_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2315),
    .D(_00563_),
    .Q_N(_13444_),
    .Q(\atari2600.ram[106][3] ));
 sg13g2_dfrbp_1 _28179_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2314),
    .D(_00564_),
    .Q_N(_13443_),
    .Q(\atari2600.ram[106][4] ));
 sg13g2_dfrbp_1 _28180_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2313),
    .D(_00565_),
    .Q_N(_13442_),
    .Q(\atari2600.ram[106][5] ));
 sg13g2_dfrbp_1 _28181_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2312),
    .D(_00566_),
    .Q_N(_13441_),
    .Q(\atari2600.ram[106][6] ));
 sg13g2_dfrbp_1 _28182_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2311),
    .D(_00567_),
    .Q_N(_13440_),
    .Q(\atari2600.ram[106][7] ));
 sg13g2_dfrbp_1 _28183_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2310),
    .D(_00568_),
    .Q_N(_13439_),
    .Q(\atari2600.ram[107][0] ));
 sg13g2_dfrbp_1 _28184_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2309),
    .D(_00569_),
    .Q_N(_13438_),
    .Q(\atari2600.ram[107][1] ));
 sg13g2_dfrbp_1 _28185_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2308),
    .D(_00570_),
    .Q_N(_13437_),
    .Q(\atari2600.ram[107][2] ));
 sg13g2_dfrbp_1 _28186_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2307),
    .D(_00571_),
    .Q_N(_13436_),
    .Q(\atari2600.ram[107][3] ));
 sg13g2_dfrbp_1 _28187_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2306),
    .D(_00572_),
    .Q_N(_13435_),
    .Q(\atari2600.ram[107][4] ));
 sg13g2_dfrbp_1 _28188_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net2305),
    .D(_00573_),
    .Q_N(_13434_),
    .Q(\atari2600.ram[107][5] ));
 sg13g2_dfrbp_1 _28189_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2304),
    .D(_00574_),
    .Q_N(_13433_),
    .Q(\atari2600.ram[107][6] ));
 sg13g2_dfrbp_1 _28190_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2303),
    .D(_00575_),
    .Q_N(_13432_),
    .Q(\atari2600.ram[107][7] ));
 sg13g2_dfrbp_1 _28191_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2302),
    .D(_00576_),
    .Q_N(_13431_),
    .Q(\atari2600.ram[108][0] ));
 sg13g2_dfrbp_1 _28192_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2301),
    .D(_00577_),
    .Q_N(_13430_),
    .Q(\atari2600.ram[108][1] ));
 sg13g2_dfrbp_1 _28193_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2300),
    .D(_00578_),
    .Q_N(_13429_),
    .Q(\atari2600.ram[108][2] ));
 sg13g2_dfrbp_1 _28194_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2299),
    .D(_00579_),
    .Q_N(_13428_),
    .Q(\atari2600.ram[108][3] ));
 sg13g2_dfrbp_1 _28195_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2298),
    .D(_00580_),
    .Q_N(_13427_),
    .Q(\atari2600.ram[108][4] ));
 sg13g2_dfrbp_1 _28196_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2297),
    .D(_00581_),
    .Q_N(_13426_),
    .Q(\atari2600.ram[108][5] ));
 sg13g2_dfrbp_1 _28197_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2296),
    .D(_00582_),
    .Q_N(_13425_),
    .Q(\atari2600.ram[108][6] ));
 sg13g2_dfrbp_1 _28198_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2295),
    .D(_00583_),
    .Q_N(_13424_),
    .Q(\atari2600.ram[108][7] ));
 sg13g2_dfrbp_1 _28199_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2294),
    .D(_00584_),
    .Q_N(_13423_),
    .Q(\atari2600.ram[10][0] ));
 sg13g2_dfrbp_1 _28200_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2293),
    .D(_00585_),
    .Q_N(_13422_),
    .Q(\atari2600.ram[10][1] ));
 sg13g2_dfrbp_1 _28201_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2292),
    .D(_00586_),
    .Q_N(_13421_),
    .Q(\atari2600.ram[10][2] ));
 sg13g2_dfrbp_1 _28202_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2291),
    .D(_00587_),
    .Q_N(_13420_),
    .Q(\atari2600.ram[10][3] ));
 sg13g2_dfrbp_1 _28203_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2290),
    .D(_00588_),
    .Q_N(_13419_),
    .Q(\atari2600.ram[10][4] ));
 sg13g2_dfrbp_1 _28204_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net2289),
    .D(_00589_),
    .Q_N(_13418_),
    .Q(\atari2600.ram[10][5] ));
 sg13g2_dfrbp_1 _28205_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2288),
    .D(_00590_),
    .Q_N(_13417_),
    .Q(\atari2600.ram[10][6] ));
 sg13g2_dfrbp_1 _28206_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2287),
    .D(_00591_),
    .Q_N(_13416_),
    .Q(\atari2600.ram[10][7] ));
 sg13g2_dfrbp_1 _28207_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2286),
    .D(_00592_),
    .Q_N(_13415_),
    .Q(\atari2600.ram[110][0] ));
 sg13g2_dfrbp_1 _28208_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2285),
    .D(_00593_),
    .Q_N(_13414_),
    .Q(\atari2600.ram[110][1] ));
 sg13g2_dfrbp_1 _28209_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2284),
    .D(_00594_),
    .Q_N(_13413_),
    .Q(\atari2600.ram[110][2] ));
 sg13g2_dfrbp_1 _28210_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2283),
    .D(_00595_),
    .Q_N(_13412_),
    .Q(\atari2600.ram[110][3] ));
 sg13g2_dfrbp_1 _28211_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2282),
    .D(_00596_),
    .Q_N(_13411_),
    .Q(\atari2600.ram[110][4] ));
 sg13g2_dfrbp_1 _28212_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2281),
    .D(_00597_),
    .Q_N(_13410_),
    .Q(\atari2600.ram[110][5] ));
 sg13g2_dfrbp_1 _28213_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2280),
    .D(_00598_),
    .Q_N(_13409_),
    .Q(\atari2600.ram[110][6] ));
 sg13g2_dfrbp_1 _28214_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2279),
    .D(_00599_),
    .Q_N(_13408_),
    .Q(\atari2600.ram[110][7] ));
 sg13g2_dfrbp_1 _28215_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2278),
    .D(_00600_),
    .Q_N(_13407_),
    .Q(\atari2600.ram[111][0] ));
 sg13g2_dfrbp_1 _28216_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net2277),
    .D(_00601_),
    .Q_N(_13406_),
    .Q(\atari2600.ram[111][1] ));
 sg13g2_dfrbp_1 _28217_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2276),
    .D(_00602_),
    .Q_N(_13405_),
    .Q(\atari2600.ram[111][2] ));
 sg13g2_dfrbp_1 _28218_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2275),
    .D(_00603_),
    .Q_N(_13404_),
    .Q(\atari2600.ram[111][3] ));
 sg13g2_dfrbp_1 _28219_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net2274),
    .D(_00604_),
    .Q_N(_13403_),
    .Q(\atari2600.ram[111][4] ));
 sg13g2_dfrbp_1 _28220_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2273),
    .D(_00605_),
    .Q_N(_13402_),
    .Q(\atari2600.ram[111][5] ));
 sg13g2_dfrbp_1 _28221_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2272),
    .D(_00606_),
    .Q_N(_13401_),
    .Q(\atari2600.ram[111][6] ));
 sg13g2_dfrbp_1 _28222_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2271),
    .D(_00607_),
    .Q_N(_13400_),
    .Q(\atari2600.ram[111][7] ));
 sg13g2_dfrbp_1 _28223_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2270),
    .D(_00608_),
    .Q_N(_13399_),
    .Q(\atari2600.ram[112][0] ));
 sg13g2_dfrbp_1 _28224_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2269),
    .D(_00609_),
    .Q_N(_13398_),
    .Q(\atari2600.ram[112][1] ));
 sg13g2_dfrbp_1 _28225_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2268),
    .D(_00610_),
    .Q_N(_13397_),
    .Q(\atari2600.ram[112][2] ));
 sg13g2_dfrbp_1 _28226_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2267),
    .D(_00611_),
    .Q_N(_13396_),
    .Q(\atari2600.ram[112][3] ));
 sg13g2_dfrbp_1 _28227_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2266),
    .D(_00612_),
    .Q_N(_13395_),
    .Q(\atari2600.ram[112][4] ));
 sg13g2_dfrbp_1 _28228_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2265),
    .D(_00613_),
    .Q_N(_13394_),
    .Q(\atari2600.ram[112][5] ));
 sg13g2_dfrbp_1 _28229_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2264),
    .D(_00614_),
    .Q_N(_13393_),
    .Q(\atari2600.ram[112][6] ));
 sg13g2_dfrbp_1 _28230_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2263),
    .D(_00615_),
    .Q_N(_13392_),
    .Q(\atari2600.ram[112][7] ));
 sg13g2_dfrbp_1 _28231_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2262),
    .D(_00616_),
    .Q_N(_13391_),
    .Q(\atari2600.ram[113][0] ));
 sg13g2_dfrbp_1 _28232_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net2261),
    .D(_00617_),
    .Q_N(_13390_),
    .Q(\atari2600.ram[113][1] ));
 sg13g2_dfrbp_1 _28233_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2260),
    .D(_00618_),
    .Q_N(_13389_),
    .Q(\atari2600.ram[113][2] ));
 sg13g2_dfrbp_1 _28234_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2259),
    .D(_00619_),
    .Q_N(_13388_),
    .Q(\atari2600.ram[113][3] ));
 sg13g2_dfrbp_1 _28235_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2258),
    .D(_00620_),
    .Q_N(_13387_),
    .Q(\atari2600.ram[113][4] ));
 sg13g2_dfrbp_1 _28236_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2257),
    .D(_00621_),
    .Q_N(_13386_),
    .Q(\atari2600.ram[113][5] ));
 sg13g2_dfrbp_1 _28237_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2256),
    .D(_00622_),
    .Q_N(_13385_),
    .Q(\atari2600.ram[113][6] ));
 sg13g2_dfrbp_1 _28238_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2255),
    .D(_00623_),
    .Q_N(_13384_),
    .Q(\atari2600.ram[113][7] ));
 sg13g2_dfrbp_1 _28239_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2254),
    .D(_00624_),
    .Q_N(_13383_),
    .Q(\atari2600.ram[114][0] ));
 sg13g2_dfrbp_1 _28240_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2253),
    .D(_00625_),
    .Q_N(_13382_),
    .Q(\atari2600.ram[114][1] ));
 sg13g2_dfrbp_1 _28241_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2252),
    .D(_00626_),
    .Q_N(_13381_),
    .Q(\atari2600.ram[114][2] ));
 sg13g2_dfrbp_1 _28242_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2251),
    .D(_00627_),
    .Q_N(_13380_),
    .Q(\atari2600.ram[114][3] ));
 sg13g2_dfrbp_1 _28243_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2250),
    .D(_00628_),
    .Q_N(_13379_),
    .Q(\atari2600.ram[114][4] ));
 sg13g2_dfrbp_1 _28244_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2249),
    .D(_00629_),
    .Q_N(_13378_),
    .Q(\atari2600.ram[114][5] ));
 sg13g2_dfrbp_1 _28245_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2248),
    .D(_00630_),
    .Q_N(_13377_),
    .Q(\atari2600.ram[114][6] ));
 sg13g2_dfrbp_1 _28246_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2247),
    .D(_00631_),
    .Q_N(_13376_),
    .Q(\atari2600.ram[114][7] ));
 sg13g2_dfrbp_1 _28247_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2246),
    .D(_00632_),
    .Q_N(_13375_),
    .Q(\atari2600.ram[115][0] ));
 sg13g2_dfrbp_1 _28248_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2245),
    .D(_00633_),
    .Q_N(_13374_),
    .Q(\atari2600.ram[115][1] ));
 sg13g2_dfrbp_1 _28249_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2244),
    .D(_00634_),
    .Q_N(_13373_),
    .Q(\atari2600.ram[115][2] ));
 sg13g2_dfrbp_1 _28250_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2243),
    .D(_00635_),
    .Q_N(_13372_),
    .Q(\atari2600.ram[115][3] ));
 sg13g2_dfrbp_1 _28251_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2242),
    .D(_00636_),
    .Q_N(_13371_),
    .Q(\atari2600.ram[115][4] ));
 sg13g2_dfrbp_1 _28252_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2241),
    .D(_00637_),
    .Q_N(_13370_),
    .Q(\atari2600.ram[115][5] ));
 sg13g2_dfrbp_1 _28253_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2240),
    .D(_00638_),
    .Q_N(_13369_),
    .Q(\atari2600.ram[115][6] ));
 sg13g2_dfrbp_1 _28254_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2239),
    .D(_00639_),
    .Q_N(_13368_),
    .Q(\atari2600.ram[115][7] ));
 sg13g2_dfrbp_1 _28255_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2238),
    .D(_00640_),
    .Q_N(_13367_),
    .Q(\atari2600.ram[116][0] ));
 sg13g2_dfrbp_1 _28256_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2237),
    .D(_00641_),
    .Q_N(_13366_),
    .Q(\atari2600.ram[116][1] ));
 sg13g2_dfrbp_1 _28257_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2236),
    .D(_00642_),
    .Q_N(_13365_),
    .Q(\atari2600.ram[116][2] ));
 sg13g2_dfrbp_1 _28258_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net2235),
    .D(_00643_),
    .Q_N(_13364_),
    .Q(\atari2600.ram[116][3] ));
 sg13g2_dfrbp_1 _28259_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2234),
    .D(_00644_),
    .Q_N(_13363_),
    .Q(\atari2600.ram[116][4] ));
 sg13g2_dfrbp_1 _28260_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2233),
    .D(_00645_),
    .Q_N(_13362_),
    .Q(\atari2600.ram[116][5] ));
 sg13g2_dfrbp_1 _28261_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net2232),
    .D(_00646_),
    .Q_N(_13361_),
    .Q(\atari2600.ram[116][6] ));
 sg13g2_dfrbp_1 _28262_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net2231),
    .D(_00647_),
    .Q_N(_13360_),
    .Q(\atari2600.ram[116][7] ));
 sg13g2_dfrbp_1 _28263_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2230),
    .D(_00648_),
    .Q_N(_13359_),
    .Q(\atari2600.ram[117][0] ));
 sg13g2_dfrbp_1 _28264_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2229),
    .D(_00649_),
    .Q_N(_13358_),
    .Q(\atari2600.ram[117][1] ));
 sg13g2_dfrbp_1 _28265_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2228),
    .D(_00650_),
    .Q_N(_13357_),
    .Q(\atari2600.ram[117][2] ));
 sg13g2_dfrbp_1 _28266_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2227),
    .D(_00651_),
    .Q_N(_13356_),
    .Q(\atari2600.ram[117][3] ));
 sg13g2_dfrbp_1 _28267_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net2226),
    .D(_00652_),
    .Q_N(_13355_),
    .Q(\atari2600.ram[117][4] ));
 sg13g2_dfrbp_1 _28268_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2225),
    .D(_00653_),
    .Q_N(_13354_),
    .Q(\atari2600.ram[117][5] ));
 sg13g2_dfrbp_1 _28269_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net2224),
    .D(_00654_),
    .Q_N(_13353_),
    .Q(\atari2600.ram[117][6] ));
 sg13g2_dfrbp_1 _28270_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2223),
    .D(_00655_),
    .Q_N(_13352_),
    .Q(\atari2600.ram[117][7] ));
 sg13g2_dfrbp_1 _28271_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2222),
    .D(_00656_),
    .Q_N(_13351_),
    .Q(\atari2600.ram[118][0] ));
 sg13g2_dfrbp_1 _28272_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2221),
    .D(_00657_),
    .Q_N(_13350_),
    .Q(\atari2600.ram[118][1] ));
 sg13g2_dfrbp_1 _28273_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2220),
    .D(_00658_),
    .Q_N(_13349_),
    .Q(\atari2600.ram[118][2] ));
 sg13g2_dfrbp_1 _28274_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net2219),
    .D(_00659_),
    .Q_N(_13348_),
    .Q(\atari2600.ram[118][3] ));
 sg13g2_dfrbp_1 _28275_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net2218),
    .D(_00660_),
    .Q_N(_13347_),
    .Q(\atari2600.ram[118][4] ));
 sg13g2_dfrbp_1 _28276_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net2217),
    .D(_00661_),
    .Q_N(_13346_),
    .Q(\atari2600.ram[118][5] ));
 sg13g2_dfrbp_1 _28277_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2216),
    .D(_00662_),
    .Q_N(_13345_),
    .Q(\atari2600.ram[118][6] ));
 sg13g2_dfrbp_1 _28278_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2215),
    .D(_00663_),
    .Q_N(_13344_),
    .Q(\atari2600.ram[118][7] ));
 sg13g2_dfrbp_1 _28279_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2214),
    .D(_00664_),
    .Q_N(_13343_),
    .Q(\atari2600.ram[11][0] ));
 sg13g2_dfrbp_1 _28280_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2213),
    .D(_00665_),
    .Q_N(_13342_),
    .Q(\atari2600.ram[11][1] ));
 sg13g2_dfrbp_1 _28281_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2212),
    .D(_00666_),
    .Q_N(_13341_),
    .Q(\atari2600.ram[11][2] ));
 sg13g2_dfrbp_1 _28282_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2211),
    .D(_00667_),
    .Q_N(_13340_),
    .Q(\atari2600.ram[11][3] ));
 sg13g2_dfrbp_1 _28283_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2210),
    .D(_00668_),
    .Q_N(_13339_),
    .Q(\atari2600.ram[11][4] ));
 sg13g2_dfrbp_1 _28284_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2209),
    .D(_00669_),
    .Q_N(_13338_),
    .Q(\atari2600.ram[11][5] ));
 sg13g2_dfrbp_1 _28285_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2208),
    .D(_00670_),
    .Q_N(_13337_),
    .Q(\atari2600.ram[11][6] ));
 sg13g2_dfrbp_1 _28286_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2207),
    .D(_00671_),
    .Q_N(_13336_),
    .Q(\atari2600.ram[11][7] ));
 sg13g2_dfrbp_1 _28287_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2206),
    .D(_00672_),
    .Q_N(_13335_),
    .Q(\atari2600.ram[120][0] ));
 sg13g2_dfrbp_1 _28288_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2205),
    .D(_00673_),
    .Q_N(_13334_),
    .Q(\atari2600.ram[120][1] ));
 sg13g2_dfrbp_1 _28289_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2204),
    .D(_00674_),
    .Q_N(_13333_),
    .Q(\atari2600.ram[120][2] ));
 sg13g2_dfrbp_1 _28290_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2203),
    .D(_00675_),
    .Q_N(_13332_),
    .Q(\atari2600.ram[120][3] ));
 sg13g2_dfrbp_1 _28291_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2202),
    .D(_00676_),
    .Q_N(_13331_),
    .Q(\atari2600.ram[120][4] ));
 sg13g2_dfrbp_1 _28292_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2201),
    .D(_00677_),
    .Q_N(_13330_),
    .Q(\atari2600.ram[120][5] ));
 sg13g2_dfrbp_1 _28293_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2200),
    .D(_00678_),
    .Q_N(_13329_),
    .Q(\atari2600.ram[120][6] ));
 sg13g2_dfrbp_1 _28294_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2199),
    .D(_00679_),
    .Q_N(_13328_),
    .Q(\atari2600.ram[120][7] ));
 sg13g2_dfrbp_1 _28295_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2198),
    .D(_00680_),
    .Q_N(_13327_),
    .Q(\atari2600.ram[121][0] ));
 sg13g2_dfrbp_1 _28296_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2197),
    .D(_00681_),
    .Q_N(_13326_),
    .Q(\atari2600.ram[121][1] ));
 sg13g2_dfrbp_1 _28297_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2196),
    .D(_00682_),
    .Q_N(_13325_),
    .Q(\atari2600.ram[121][2] ));
 sg13g2_dfrbp_1 _28298_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2195),
    .D(_00683_),
    .Q_N(_13324_),
    .Q(\atari2600.ram[121][3] ));
 sg13g2_dfrbp_1 _28299_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2194),
    .D(_00684_),
    .Q_N(_13323_),
    .Q(\atari2600.ram[121][4] ));
 sg13g2_dfrbp_1 _28300_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2193),
    .D(_00685_),
    .Q_N(_13322_),
    .Q(\atari2600.ram[121][5] ));
 sg13g2_dfrbp_1 _28301_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2192),
    .D(_00686_),
    .Q_N(_13321_),
    .Q(\atari2600.ram[121][6] ));
 sg13g2_dfrbp_1 _28302_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2191),
    .D(_00687_),
    .Q_N(_13320_),
    .Q(\atari2600.ram[121][7] ));
 sg13g2_dfrbp_1 _28303_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2190),
    .D(_00688_),
    .Q_N(_13319_),
    .Q(\atari2600.ram[122][0] ));
 sg13g2_dfrbp_1 _28304_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2189),
    .D(_00689_),
    .Q_N(_13318_),
    .Q(\atari2600.ram[122][1] ));
 sg13g2_dfrbp_1 _28305_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2188),
    .D(_00690_),
    .Q_N(_13317_),
    .Q(\atari2600.ram[122][2] ));
 sg13g2_dfrbp_1 _28306_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2187),
    .D(_00691_),
    .Q_N(_13316_),
    .Q(\atari2600.ram[122][3] ));
 sg13g2_dfrbp_1 _28307_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2186),
    .D(_00692_),
    .Q_N(_13315_),
    .Q(\atari2600.ram[122][4] ));
 sg13g2_dfrbp_1 _28308_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2185),
    .D(_00693_),
    .Q_N(_13314_),
    .Q(\atari2600.ram[122][5] ));
 sg13g2_dfrbp_1 _28309_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2184),
    .D(_00694_),
    .Q_N(_13313_),
    .Q(\atari2600.ram[122][6] ));
 sg13g2_dfrbp_1 _28310_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2183),
    .D(_00695_),
    .Q_N(_13312_),
    .Q(\atari2600.ram[122][7] ));
 sg13g2_dfrbp_1 _28311_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2182),
    .D(_00696_),
    .Q_N(_13311_),
    .Q(\atari2600.ram[123][0] ));
 sg13g2_dfrbp_1 _28312_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2181),
    .D(_00697_),
    .Q_N(_13310_),
    .Q(\atari2600.ram[123][1] ));
 sg13g2_dfrbp_1 _28313_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2180),
    .D(_00698_),
    .Q_N(_13309_),
    .Q(\atari2600.ram[123][2] ));
 sg13g2_dfrbp_1 _28314_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2179),
    .D(_00699_),
    .Q_N(_13308_),
    .Q(\atari2600.ram[123][3] ));
 sg13g2_dfrbp_1 _28315_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2178),
    .D(_00700_),
    .Q_N(_13307_),
    .Q(\atari2600.ram[123][4] ));
 sg13g2_dfrbp_1 _28316_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2177),
    .D(_00701_),
    .Q_N(_13306_),
    .Q(\atari2600.ram[123][5] ));
 sg13g2_dfrbp_1 _28317_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2176),
    .D(_00702_),
    .Q_N(_13305_),
    .Q(\atari2600.ram[123][6] ));
 sg13g2_dfrbp_1 _28318_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2175),
    .D(_00703_),
    .Q_N(_13304_),
    .Q(\atari2600.ram[123][7] ));
 sg13g2_dfrbp_1 _28319_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2174),
    .D(_00704_),
    .Q_N(_13303_),
    .Q(\atari2600.ram[124][0] ));
 sg13g2_dfrbp_1 _28320_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net2173),
    .D(_00705_),
    .Q_N(_13302_),
    .Q(\atari2600.ram[124][1] ));
 sg13g2_dfrbp_1 _28321_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2172),
    .D(_00706_),
    .Q_N(_13301_),
    .Q(\atari2600.ram[124][2] ));
 sg13g2_dfrbp_1 _28322_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2171),
    .D(_00707_),
    .Q_N(_13300_),
    .Q(\atari2600.ram[124][3] ));
 sg13g2_dfrbp_1 _28323_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2170),
    .D(_00708_),
    .Q_N(_13299_),
    .Q(\atari2600.ram[124][4] ));
 sg13g2_dfrbp_1 _28324_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net2169),
    .D(_00709_),
    .Q_N(_13298_),
    .Q(\atari2600.ram[124][5] ));
 sg13g2_dfrbp_1 _28325_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net2168),
    .D(_00710_),
    .Q_N(_13297_),
    .Q(\atari2600.ram[124][6] ));
 sg13g2_dfrbp_1 _28326_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net2167),
    .D(_00711_),
    .Q_N(_13296_),
    .Q(\atari2600.ram[124][7] ));
 sg13g2_dfrbp_1 _28327_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2166),
    .D(_00712_),
    .Q_N(_13295_),
    .Q(\atari2600.ram[125][0] ));
 sg13g2_dfrbp_1 _28328_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net2165),
    .D(_00713_),
    .Q_N(_13294_),
    .Q(\atari2600.ram[125][1] ));
 sg13g2_dfrbp_1 _28329_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2164),
    .D(_00714_),
    .Q_N(_13293_),
    .Q(\atari2600.ram[125][2] ));
 sg13g2_dfrbp_1 _28330_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2163),
    .D(_00715_),
    .Q_N(_13292_),
    .Q(\atari2600.ram[125][3] ));
 sg13g2_dfrbp_1 _28331_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2162),
    .D(_00716_),
    .Q_N(_13291_),
    .Q(\atari2600.ram[125][4] ));
 sg13g2_dfrbp_1 _28332_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2161),
    .D(_00717_),
    .Q_N(_13290_),
    .Q(\atari2600.ram[125][5] ));
 sg13g2_dfrbp_1 _28333_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net2160),
    .D(_00718_),
    .Q_N(_13289_),
    .Q(\atari2600.ram[125][6] ));
 sg13g2_dfrbp_1 _28334_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2159),
    .D(_00719_),
    .Q_N(_13288_),
    .Q(\atari2600.ram[125][7] ));
 sg13g2_dfrbp_1 _28335_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2158),
    .D(_00720_),
    .Q_N(_13287_),
    .Q(\atari2600.ram[126][0] ));
 sg13g2_dfrbp_1 _28336_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net2157),
    .D(_00721_),
    .Q_N(_13286_),
    .Q(\atari2600.ram[126][1] ));
 sg13g2_dfrbp_1 _28337_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2156),
    .D(_00722_),
    .Q_N(_13285_),
    .Q(\atari2600.ram[126][2] ));
 sg13g2_dfrbp_1 _28338_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2155),
    .D(_00723_),
    .Q_N(_13284_),
    .Q(\atari2600.ram[126][3] ));
 sg13g2_dfrbp_1 _28339_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2154),
    .D(_00724_),
    .Q_N(_13283_),
    .Q(\atari2600.ram[126][4] ));
 sg13g2_dfrbp_1 _28340_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2153),
    .D(_00725_),
    .Q_N(_13282_),
    .Q(\atari2600.ram[126][5] ));
 sg13g2_dfrbp_1 _28341_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net2152),
    .D(_00726_),
    .Q_N(_13281_),
    .Q(\atari2600.ram[126][6] ));
 sg13g2_dfrbp_1 _28342_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net2151),
    .D(_00727_),
    .Q_N(_13280_),
    .Q(\atari2600.ram[126][7] ));
 sg13g2_dfrbp_1 _28343_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2150),
    .D(_00728_),
    .Q_N(_13279_),
    .Q(\atari2600.ram[92][0] ));
 sg13g2_dfrbp_1 _28344_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2149),
    .D(_00729_),
    .Q_N(_13278_),
    .Q(\atari2600.ram[92][1] ));
 sg13g2_dfrbp_1 _28345_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2148),
    .D(_00730_),
    .Q_N(_13277_),
    .Q(\atari2600.ram[92][2] ));
 sg13g2_dfrbp_1 _28346_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2147),
    .D(_00731_),
    .Q_N(_13276_),
    .Q(\atari2600.ram[92][3] ));
 sg13g2_dfrbp_1 _28347_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2146),
    .D(_00732_),
    .Q_N(_13275_),
    .Q(\atari2600.ram[92][4] ));
 sg13g2_dfrbp_1 _28348_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2145),
    .D(_00733_),
    .Q_N(_13274_),
    .Q(\atari2600.ram[92][5] ));
 sg13g2_dfrbp_1 _28349_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2144),
    .D(_00734_),
    .Q_N(_13273_),
    .Q(\atari2600.ram[92][6] ));
 sg13g2_dfrbp_1 _28350_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2143),
    .D(_00735_),
    .Q_N(_13272_),
    .Q(\atari2600.ram[92][7] ));
 sg13g2_dfrbp_1 _28351_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2142),
    .D(_00736_),
    .Q_N(_13271_),
    .Q(\atari2600.cpu.AXYS[3][0] ));
 sg13g2_dfrbp_1 _28352_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2141),
    .D(_00737_),
    .Q_N(_13270_),
    .Q(\atari2600.cpu.AXYS[3][1] ));
 sg13g2_dfrbp_1 _28353_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2140),
    .D(_00738_),
    .Q_N(_13269_),
    .Q(\atari2600.cpu.AXYS[3][2] ));
 sg13g2_dfrbp_1 _28354_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2139),
    .D(_00739_),
    .Q_N(_13268_),
    .Q(\atari2600.cpu.AXYS[3][3] ));
 sg13g2_dfrbp_1 _28355_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2138),
    .D(net3335),
    .Q_N(_13267_),
    .Q(\atari2600.cpu.AXYS[3][4] ));
 sg13g2_dfrbp_1 _28356_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2137),
    .D(_00741_),
    .Q_N(_13266_),
    .Q(\atari2600.cpu.AXYS[3][5] ));
 sg13g2_dfrbp_1 _28357_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2136),
    .D(_00742_),
    .Q_N(_13265_),
    .Q(\atari2600.cpu.AXYS[3][6] ));
 sg13g2_dfrbp_1 _28358_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2135),
    .D(_00743_),
    .Q_N(_13264_),
    .Q(\atari2600.cpu.AXYS[3][7] ));
 sg13g2_dfrbp_1 _28359_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2134),
    .D(_00744_),
    .Q_N(_13263_),
    .Q(\atari2600.ram[19][0] ));
 sg13g2_dfrbp_1 _28360_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net2133),
    .D(_00745_),
    .Q_N(_13262_),
    .Q(\atari2600.ram[19][1] ));
 sg13g2_dfrbp_1 _28361_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net2132),
    .D(_00746_),
    .Q_N(_13261_),
    .Q(\atari2600.ram[19][2] ));
 sg13g2_dfrbp_1 _28362_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2131),
    .D(_00747_),
    .Q_N(_13260_),
    .Q(\atari2600.ram[19][3] ));
 sg13g2_dfrbp_1 _28363_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2130),
    .D(_00748_),
    .Q_N(_13259_),
    .Q(\atari2600.ram[19][4] ));
 sg13g2_dfrbp_1 _28364_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2129),
    .D(_00749_),
    .Q_N(_13258_),
    .Q(\atari2600.ram[19][5] ));
 sg13g2_dfrbp_1 _28365_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2128),
    .D(_00750_),
    .Q_N(_13257_),
    .Q(\atari2600.ram[19][6] ));
 sg13g2_dfrbp_1 _28366_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net2127),
    .D(_00751_),
    .Q_N(_13256_),
    .Q(\atari2600.ram[19][7] ));
 sg13g2_dfrbp_1 _28367_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2126),
    .D(_00752_),
    .Q_N(_13255_),
    .Q(\atari2600.ram[29][0] ));
 sg13g2_dfrbp_1 _28368_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2125),
    .D(_00753_),
    .Q_N(_13254_),
    .Q(\atari2600.ram[29][1] ));
 sg13g2_dfrbp_1 _28369_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2124),
    .D(_00754_),
    .Q_N(_13253_),
    .Q(\atari2600.ram[29][2] ));
 sg13g2_dfrbp_1 _28370_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2123),
    .D(_00755_),
    .Q_N(_13252_),
    .Q(\atari2600.ram[29][3] ));
 sg13g2_dfrbp_1 _28371_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2122),
    .D(_00756_),
    .Q_N(_13251_),
    .Q(\atari2600.ram[29][4] ));
 sg13g2_dfrbp_1 _28372_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2121),
    .D(_00757_),
    .Q_N(_13250_),
    .Q(\atari2600.ram[29][5] ));
 sg13g2_dfrbp_1 _28373_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2120),
    .D(_00758_),
    .Q_N(_13249_),
    .Q(\atari2600.ram[29][6] ));
 sg13g2_dfrbp_1 _28374_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2119),
    .D(_00759_),
    .Q_N(_13248_),
    .Q(\atari2600.ram[29][7] ));
 sg13g2_dfrbp_1 _28375_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2118),
    .D(_00760_),
    .Q_N(_13247_),
    .Q(\atari2600.ram[39][0] ));
 sg13g2_dfrbp_1 _28376_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2117),
    .D(_00761_),
    .Q_N(_13246_),
    .Q(\atari2600.ram[39][1] ));
 sg13g2_dfrbp_1 _28377_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2116),
    .D(_00762_),
    .Q_N(_13245_),
    .Q(\atari2600.ram[39][2] ));
 sg13g2_dfrbp_1 _28378_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2115),
    .D(_00763_),
    .Q_N(_13244_),
    .Q(\atari2600.ram[39][3] ));
 sg13g2_dfrbp_1 _28379_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2114),
    .D(_00764_),
    .Q_N(_13243_),
    .Q(\atari2600.ram[39][4] ));
 sg13g2_dfrbp_1 _28380_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net2113),
    .D(_00765_),
    .Q_N(_13242_),
    .Q(\atari2600.ram[39][5] ));
 sg13g2_dfrbp_1 _28381_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2112),
    .D(_00766_),
    .Q_N(_13241_),
    .Q(\atari2600.ram[39][6] ));
 sg13g2_dfrbp_1 _28382_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2111),
    .D(_00767_),
    .Q_N(_13240_),
    .Q(\atari2600.ram[39][7] ));
 sg13g2_dfrbp_1 _28383_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2110),
    .D(_00768_),
    .Q_N(_13239_),
    .Q(\atari2600.ram[49][0] ));
 sg13g2_dfrbp_1 _28384_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2109),
    .D(_00769_),
    .Q_N(_13238_),
    .Q(\atari2600.ram[49][1] ));
 sg13g2_dfrbp_1 _28385_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net2108),
    .D(_00770_),
    .Q_N(_13237_),
    .Q(\atari2600.ram[49][2] ));
 sg13g2_dfrbp_1 _28386_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net2107),
    .D(_00771_),
    .Q_N(_13236_),
    .Q(\atari2600.ram[49][3] ));
 sg13g2_dfrbp_1 _28387_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2106),
    .D(_00772_),
    .Q_N(_13235_),
    .Q(\atari2600.ram[49][4] ));
 sg13g2_dfrbp_1 _28388_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2105),
    .D(_00773_),
    .Q_N(_13234_),
    .Q(\atari2600.ram[49][5] ));
 sg13g2_dfrbp_1 _28389_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net2104),
    .D(_00774_),
    .Q_N(_13233_),
    .Q(\atari2600.ram[49][6] ));
 sg13g2_dfrbp_1 _28390_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2103),
    .D(_00775_),
    .Q_N(_13232_),
    .Q(\atari2600.ram[49][7] ));
 sg13g2_dfrbp_1 _28391_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2102),
    .D(_00776_),
    .Q_N(_13231_),
    .Q(\atari2600.ram[59][0] ));
 sg13g2_dfrbp_1 _28392_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2101),
    .D(_00777_),
    .Q_N(_13230_),
    .Q(\atari2600.ram[59][1] ));
 sg13g2_dfrbp_1 _28393_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net2100),
    .D(_00778_),
    .Q_N(_13229_),
    .Q(\atari2600.ram[59][2] ));
 sg13g2_dfrbp_1 _28394_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2099),
    .D(_00779_),
    .Q_N(_13228_),
    .Q(\atari2600.ram[59][3] ));
 sg13g2_dfrbp_1 _28395_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2098),
    .D(_00780_),
    .Q_N(_13227_),
    .Q(\atari2600.ram[59][4] ));
 sg13g2_dfrbp_1 _28396_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2097),
    .D(_00781_),
    .Q_N(_13226_),
    .Q(\atari2600.ram[59][5] ));
 sg13g2_dfrbp_1 _28397_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2096),
    .D(_00782_),
    .Q_N(_13225_),
    .Q(\atari2600.ram[59][6] ));
 sg13g2_dfrbp_1 _28398_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2095),
    .D(_00783_),
    .Q_N(_13224_),
    .Q(\atari2600.ram[59][7] ));
 sg13g2_dfrbp_1 _28399_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2094),
    .D(_00784_),
    .Q_N(_13223_),
    .Q(\atari2600.ram[69][0] ));
 sg13g2_dfrbp_1 _28400_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2093),
    .D(_00785_),
    .Q_N(_13222_),
    .Q(\atari2600.ram[69][1] ));
 sg13g2_dfrbp_1 _28401_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2092),
    .D(_00786_),
    .Q_N(_13221_),
    .Q(\atari2600.ram[69][2] ));
 sg13g2_dfrbp_1 _28402_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2091),
    .D(_00787_),
    .Q_N(_13220_),
    .Q(\atari2600.ram[69][3] ));
 sg13g2_dfrbp_1 _28403_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2090),
    .D(_00788_),
    .Q_N(_13219_),
    .Q(\atari2600.ram[69][4] ));
 sg13g2_dfrbp_1 _28404_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2089),
    .D(_00789_),
    .Q_N(_13218_),
    .Q(\atari2600.ram[69][5] ));
 sg13g2_dfrbp_1 _28405_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2088),
    .D(_00790_),
    .Q_N(_13217_),
    .Q(\atari2600.ram[69][6] ));
 sg13g2_dfrbp_1 _28406_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2087),
    .D(_00791_),
    .Q_N(_13216_),
    .Q(\atari2600.ram[69][7] ));
 sg13g2_dfrbp_1 _28407_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net2086),
    .D(_00792_),
    .Q_N(_13215_),
    .Q(\atari2600.ram[79][0] ));
 sg13g2_dfrbp_1 _28408_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2085),
    .D(_00793_),
    .Q_N(_13214_),
    .Q(\atari2600.ram[79][1] ));
 sg13g2_dfrbp_1 _28409_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2084),
    .D(_00794_),
    .Q_N(_13213_),
    .Q(\atari2600.ram[79][2] ));
 sg13g2_dfrbp_1 _28410_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net2083),
    .D(_00795_),
    .Q_N(_13212_),
    .Q(\atari2600.ram[79][3] ));
 sg13g2_dfrbp_1 _28411_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net2082),
    .D(_00796_),
    .Q_N(_13211_),
    .Q(\atari2600.ram[79][4] ));
 sg13g2_dfrbp_1 _28412_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net2081),
    .D(_00797_),
    .Q_N(_13210_),
    .Q(\atari2600.ram[79][5] ));
 sg13g2_dfrbp_1 _28413_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net2080),
    .D(_00798_),
    .Q_N(_13209_),
    .Q(\atari2600.ram[79][6] ));
 sg13g2_dfrbp_1 _28414_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net2079),
    .D(_00799_),
    .Q_N(_13208_),
    .Q(\atari2600.ram[79][7] ));
 sg13g2_dfrbp_1 _28415_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2078),
    .D(_00800_),
    .Q_N(_13207_),
    .Q(\atari2600.ram[89][0] ));
 sg13g2_dfrbp_1 _28416_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2077),
    .D(_00801_),
    .Q_N(_13206_),
    .Q(\atari2600.ram[89][1] ));
 sg13g2_dfrbp_1 _28417_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2076),
    .D(_00802_),
    .Q_N(_13205_),
    .Q(\atari2600.ram[89][2] ));
 sg13g2_dfrbp_1 _28418_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2075),
    .D(_00803_),
    .Q_N(_13204_),
    .Q(\atari2600.ram[89][3] ));
 sg13g2_dfrbp_1 _28419_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2074),
    .D(_00804_),
    .Q_N(_13203_),
    .Q(\atari2600.ram[89][4] ));
 sg13g2_dfrbp_1 _28420_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2073),
    .D(_00805_),
    .Q_N(_13202_),
    .Q(\atari2600.ram[89][5] ));
 sg13g2_dfrbp_1 _28421_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2072),
    .D(_00806_),
    .Q_N(_13201_),
    .Q(\atari2600.ram[89][6] ));
 sg13g2_dfrbp_1 _28422_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2071),
    .D(_00807_),
    .Q_N(_13200_),
    .Q(\atari2600.ram[89][7] ));
 sg13g2_dfrbp_1 _28423_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2070),
    .D(_00808_),
    .Q_N(_13199_),
    .Q(\atari2600.ram[99][0] ));
 sg13g2_dfrbp_1 _28424_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2069),
    .D(_00809_),
    .Q_N(_13198_),
    .Q(\atari2600.ram[99][1] ));
 sg13g2_dfrbp_1 _28425_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2068),
    .D(_00810_),
    .Q_N(_13197_),
    .Q(\atari2600.ram[99][2] ));
 sg13g2_dfrbp_1 _28426_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2067),
    .D(_00811_),
    .Q_N(_13196_),
    .Q(\atari2600.ram[99][3] ));
 sg13g2_dfrbp_1 _28427_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2066),
    .D(_00812_),
    .Q_N(_13195_),
    .Q(\atari2600.ram[99][4] ));
 sg13g2_dfrbp_1 _28428_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2065),
    .D(_00813_),
    .Q_N(_13194_),
    .Q(\atari2600.ram[99][5] ));
 sg13g2_dfrbp_1 _28429_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2064),
    .D(_00814_),
    .Q_N(_13193_),
    .Q(\atari2600.ram[99][6] ));
 sg13g2_dfrbp_1 _28430_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2063),
    .D(_00815_),
    .Q_N(_13192_),
    .Q(\atari2600.ram[99][7] ));
 sg13g2_dfrbp_1 _28431_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net2062),
    .D(_00816_),
    .Q_N(_13191_),
    .Q(\atari2600.ram[109][0] ));
 sg13g2_dfrbp_1 _28432_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net2061),
    .D(_00817_),
    .Q_N(_13190_),
    .Q(\atari2600.ram[109][1] ));
 sg13g2_dfrbp_1 _28433_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2060),
    .D(_00818_),
    .Q_N(_13189_),
    .Q(\atari2600.ram[109][2] ));
 sg13g2_dfrbp_1 _28434_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2059),
    .D(_00819_),
    .Q_N(_13188_),
    .Q(\atari2600.ram[109][3] ));
 sg13g2_dfrbp_1 _28435_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2058),
    .D(_00820_),
    .Q_N(_13187_),
    .Q(\atari2600.ram[109][4] ));
 sg13g2_dfrbp_1 _28436_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net2057),
    .D(_00821_),
    .Q_N(_13186_),
    .Q(\atari2600.ram[109][5] ));
 sg13g2_dfrbp_1 _28437_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2056),
    .D(_00822_),
    .Q_N(_13185_),
    .Q(\atari2600.ram[109][6] ));
 sg13g2_dfrbp_1 _28438_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net2055),
    .D(_00823_),
    .Q_N(_13184_),
    .Q(\atari2600.ram[109][7] ));
 sg13g2_dfrbp_1 _28439_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net2054),
    .D(_00824_),
    .Q_N(_13183_),
    .Q(\atari2600.ram[119][0] ));
 sg13g2_dfrbp_1 _28440_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2053),
    .D(_00825_),
    .Q_N(_13182_),
    .Q(\atari2600.ram[119][1] ));
 sg13g2_dfrbp_1 _28441_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net2052),
    .D(_00826_),
    .Q_N(_13181_),
    .Q(\atari2600.ram[119][2] ));
 sg13g2_dfrbp_1 _28442_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2051),
    .D(_00827_),
    .Q_N(_13180_),
    .Q(\atari2600.ram[119][3] ));
 sg13g2_dfrbp_1 _28443_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net2050),
    .D(_00828_),
    .Q_N(_13179_),
    .Q(\atari2600.ram[119][4] ));
 sg13g2_dfrbp_1 _28444_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net2049),
    .D(_00829_),
    .Q_N(_13178_),
    .Q(\atari2600.ram[119][5] ));
 sg13g2_dfrbp_1 _28445_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net2048),
    .D(_00830_),
    .Q_N(_13177_),
    .Q(\atari2600.ram[119][6] ));
 sg13g2_dfrbp_1 _28446_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net2047),
    .D(_00831_),
    .Q_N(_13176_),
    .Q(\atari2600.ram[119][7] ));
 sg13g2_dfrbp_1 _28447_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net2046),
    .D(_00832_),
    .Q_N(_13175_),
    .Q(\atari2600.ram[74][0] ));
 sg13g2_dfrbp_1 _28448_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2045),
    .D(_00833_),
    .Q_N(_13174_),
    .Q(\atari2600.ram[74][1] ));
 sg13g2_dfrbp_1 _28449_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2044),
    .D(_00834_),
    .Q_N(_13173_),
    .Q(\atari2600.ram[74][2] ));
 sg13g2_dfrbp_1 _28450_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2043),
    .D(_00835_),
    .Q_N(_13172_),
    .Q(\atari2600.ram[74][3] ));
 sg13g2_dfrbp_1 _28451_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net2042),
    .D(_00836_),
    .Q_N(_13171_),
    .Q(\atari2600.ram[74][4] ));
 sg13g2_dfrbp_1 _28452_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net2041),
    .D(_00837_),
    .Q_N(_13170_),
    .Q(\atari2600.ram[74][5] ));
 sg13g2_dfrbp_1 _28453_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net2040),
    .D(_00838_),
    .Q_N(_13169_),
    .Q(\atari2600.ram[74][6] ));
 sg13g2_dfrbp_1 _28454_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net2039),
    .D(_00839_),
    .Q_N(_13168_),
    .Q(\atari2600.ram[74][7] ));
 sg13g2_dfrbp_1 _28455_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net2038),
    .D(_00840_),
    .Q_N(_13167_),
    .Q(\atari2600.ram[75][0] ));
 sg13g2_dfrbp_1 _28456_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2037),
    .D(_00841_),
    .Q_N(_13166_),
    .Q(\atari2600.ram[75][1] ));
 sg13g2_dfrbp_1 _28457_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net2036),
    .D(_00842_),
    .Q_N(_13165_),
    .Q(\atari2600.ram[75][2] ));
 sg13g2_dfrbp_1 _28458_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net2035),
    .D(_00843_),
    .Q_N(_13164_),
    .Q(\atari2600.ram[75][3] ));
 sg13g2_dfrbp_1 _28459_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2034),
    .D(_00844_),
    .Q_N(_13163_),
    .Q(\atari2600.ram[75][4] ));
 sg13g2_dfrbp_1 _28460_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2033),
    .D(_00845_),
    .Q_N(_13162_),
    .Q(\atari2600.ram[75][5] ));
 sg13g2_dfrbp_1 _28461_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net2032),
    .D(_00846_),
    .Q_N(_13161_),
    .Q(\atari2600.ram[75][6] ));
 sg13g2_dfrbp_1 _28462_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net2031),
    .D(_00847_),
    .Q_N(_13160_),
    .Q(\atari2600.ram[75][7] ));
 sg13g2_dfrbp_1 _28463_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net2030),
    .D(_00848_),
    .Q_N(_13159_),
    .Q(\atari2600.ram[35][0] ));
 sg13g2_dfrbp_1 _28464_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2029),
    .D(_00849_),
    .Q_N(_13158_),
    .Q(\atari2600.ram[35][1] ));
 sg13g2_dfrbp_1 _28465_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2028),
    .D(_00850_),
    .Q_N(_13157_),
    .Q(\atari2600.ram[35][2] ));
 sg13g2_dfrbp_1 _28466_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2027),
    .D(_00851_),
    .Q_N(_13156_),
    .Q(\atari2600.ram[35][3] ));
 sg13g2_dfrbp_1 _28467_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2026),
    .D(_00852_),
    .Q_N(_13155_),
    .Q(\atari2600.ram[35][4] ));
 sg13g2_dfrbp_1 _28468_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2025),
    .D(_00853_),
    .Q_N(_13154_),
    .Q(\atari2600.ram[35][5] ));
 sg13g2_dfrbp_1 _28469_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net2024),
    .D(_00854_),
    .Q_N(_13153_),
    .Q(\atari2600.ram[35][6] ));
 sg13g2_dfrbp_1 _28470_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2023),
    .D(_00855_),
    .Q_N(_13152_),
    .Q(\atari2600.ram[35][7] ));
 sg13g2_dfrbp_1 _28471_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2022),
    .D(_00856_),
    .Q_N(_13151_),
    .Q(\atari2600.cpu.ALU.BI7 ));
 sg13g2_dfrbp_1 _28472_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net2021),
    .D(net7271),
    .Q_N(_13150_),
    .Q(\atari2600.pia.diag[0] ));
 sg13g2_dfrbp_1 _28473_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2020),
    .D(_00858_),
    .Q_N(_13149_),
    .Q(\atari2600.pia.diag[1] ));
 sg13g2_dfrbp_1 _28474_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2019),
    .D(net7314),
    .Q_N(_13148_),
    .Q(\atari2600.pia.diag[2] ));
 sg13g2_dfrbp_1 _28475_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2018),
    .D(net7109),
    .Q_N(_13147_),
    .Q(\atari2600.pia.diag[3] ));
 sg13g2_dfrbp_1 _28476_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2017),
    .D(net7275),
    .Q_N(_13146_),
    .Q(\atari2600.pia.diag[4] ));
 sg13g2_dfrbp_1 _28477_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net2016),
    .D(_00862_),
    .Q_N(_13145_),
    .Q(\atari2600.pia.diag[5] ));
 sg13g2_dfrbp_1 _28478_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2015),
    .D(net7278),
    .Q_N(_13144_),
    .Q(\atari2600.pia.diag[6] ));
 sg13g2_dfrbp_1 _28479_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2014),
    .D(_00864_),
    .Q_N(_13143_),
    .Q(\atari2600.pia.diag[7] ));
 sg13g2_dfrbp_1 _28480_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2013),
    .D(net3727),
    .Q_N(_13142_),
    .Q(\atari2600.pia.instat[1] ));
 sg13g2_dfrbp_1 _28481_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2012),
    .D(_00866_),
    .Q_N(_13141_),
    .Q(\atari2600.pia.dat_o[0] ));
 sg13g2_dfrbp_1 _28482_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2011),
    .D(net4493),
    .Q_N(_13140_),
    .Q(\atari2600.pia.dat_o[1] ));
 sg13g2_dfrbp_1 _28483_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2010),
    .D(net4644),
    .Q_N(_13139_),
    .Q(\atari2600.pia.dat_o[2] ));
 sg13g2_dfrbp_1 _28484_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2009),
    .D(net7129),
    .Q_N(_13138_),
    .Q(\atari2600.pia.dat_o[3] ));
 sg13g2_dfrbp_1 _28485_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2008),
    .D(net7168),
    .Q_N(_13137_),
    .Q(\atari2600.pia.dat_o[4] ));
 sg13g2_dfrbp_1 _28486_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2007),
    .D(net7158),
    .Q_N(_13136_),
    .Q(\atari2600.pia.dat_o[5] ));
 sg13g2_dfrbp_1 _28487_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2006),
    .D(net4460),
    .Q_N(_13135_),
    .Q(\atari2600.pia.dat_o[6] ));
 sg13g2_dfrbp_1 _28488_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2005),
    .D(net4780),
    .Q_N(_13134_),
    .Q(\atari2600.pia.dat_o[7] ));
 sg13g2_dfrbp_1 _28489_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2004),
    .D(_00874_),
    .Q_N(_13133_),
    .Q(\atari2600.pia.time_counter[0] ));
 sg13g2_dfrbp_1 _28490_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net2003),
    .D(_00875_),
    .Q_N(_13132_),
    .Q(\atari2600.pia.time_counter[1] ));
 sg13g2_dfrbp_1 _28491_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2002),
    .D(_00876_),
    .Q_N(_13131_),
    .Q(\atari2600.pia.time_counter[2] ));
 sg13g2_dfrbp_1 _28492_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2001),
    .D(_00877_),
    .Q_N(_13130_),
    .Q(\atari2600.pia.time_counter[3] ));
 sg13g2_dfrbp_1 _28493_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2000),
    .D(_00878_),
    .Q_N(_13129_),
    .Q(\atari2600.pia.time_counter[4] ));
 sg13g2_dfrbp_1 _28494_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1999),
    .D(_00879_),
    .Q_N(_13128_),
    .Q(\atari2600.pia.time_counter[5] ));
 sg13g2_dfrbp_1 _28495_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1998),
    .D(_00880_),
    .Q_N(_00083_),
    .Q(\atari2600.pia.time_counter[6] ));
 sg13g2_dfrbp_1 _28496_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1997),
    .D(net7339),
    .Q_N(_13127_),
    .Q(\atari2600.pia.time_counter[7] ));
 sg13g2_dfrbp_1 _28497_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1996),
    .D(net7019),
    .Q_N(_13126_),
    .Q(\atari2600.pia.time_counter[8] ));
 sg13g2_dfrbp_1 _28498_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1995),
    .D(_00883_),
    .Q_N(_13125_),
    .Q(\atari2600.pia.time_counter[9] ));
 sg13g2_dfrbp_1 _28499_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1994),
    .D(_00884_),
    .Q_N(_00084_),
    .Q(\atari2600.pia.time_counter[10] ));
 sg13g2_dfrbp_1 _28500_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1993),
    .D(_00885_),
    .Q_N(_13124_),
    .Q(\atari2600.pia.time_counter[11] ));
 sg13g2_dfrbp_1 _28501_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1992),
    .D(_00886_),
    .Q_N(_13123_),
    .Q(\atari2600.pia.time_counter[12] ));
 sg13g2_dfrbp_1 _28502_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1991),
    .D(_00887_),
    .Q_N(_13122_),
    .Q(\atari2600.pia.time_counter[13] ));
 sg13g2_dfrbp_1 _28503_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1990),
    .D(_00888_),
    .Q_N(_13121_),
    .Q(\atari2600.pia.time_counter[14] ));
 sg13g2_dfrbp_1 _28504_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1989),
    .D(net6598),
    .Q_N(_13120_),
    .Q(\atari2600.pia.time_counter[15] ));
 sg13g2_dfrbp_1 _28505_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1988),
    .D(net7025),
    .Q_N(_13119_),
    .Q(\atari2600.pia.time_counter[16] ));
 sg13g2_dfrbp_1 _28506_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1987),
    .D(_00891_),
    .Q_N(_13118_),
    .Q(\atari2600.pia.time_counter[17] ));
 sg13g2_dfrbp_1 _28507_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1986),
    .D(_00892_),
    .Q_N(_13117_),
    .Q(\atari2600.pia.time_counter[18] ));
 sg13g2_dfrbp_1 _28508_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1985),
    .D(_00893_),
    .Q_N(_13116_),
    .Q(\atari2600.pia.time_counter[19] ));
 sg13g2_dfrbp_1 _28509_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1984),
    .D(_00894_),
    .Q_N(_13115_),
    .Q(\atari2600.pia.time_counter[20] ));
 sg13g2_dfrbp_1 _28510_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1983),
    .D(_00895_),
    .Q_N(_13114_),
    .Q(\atari2600.pia.time_counter[21] ));
 sg13g2_dfrbp_1 _28511_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1981),
    .D(net3619),
    .Q_N(_13113_),
    .Q(\atari2600.pia.time_counter[22] ));
 sg13g2_dfrbp_1 _28512_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1979),
    .D(_00897_),
    .Q_N(_13112_),
    .Q(\atari2600.pia.time_counter[23] ));
 sg13g2_dfrbp_1 _28513_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1977),
    .D(_00898_),
    .Q_N(_13111_),
    .Q(\atari2600.pia.underflow ));
 sg13g2_dfrbp_1 _28514_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1976),
    .D(_00899_),
    .Q_N(_13110_),
    .Q(\atari2600.pia.reset_timer[0] ));
 sg13g2_dfrbp_1 _28515_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1975),
    .D(_00900_),
    .Q_N(_13109_),
    .Q(\atari2600.pia.reset_timer[1] ));
 sg13g2_dfrbp_1 _28516_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1974),
    .D(_00901_),
    .Q_N(_13108_),
    .Q(\atari2600.pia.reset_timer[2] ));
 sg13g2_dfrbp_1 _28517_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1973),
    .D(_00902_),
    .Q_N(_13107_),
    .Q(\atari2600.pia.reset_timer[3] ));
 sg13g2_dfrbp_1 _28518_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1972),
    .D(_00903_),
    .Q_N(_13106_),
    .Q(\atari2600.pia.reset_timer[4] ));
 sg13g2_dfrbp_1 _28519_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1971),
    .D(_00904_),
    .Q_N(_13105_),
    .Q(\atari2600.pia.reset_timer[5] ));
 sg13g2_dfrbp_1 _28520_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1970),
    .D(_00905_),
    .Q_N(_13104_),
    .Q(\atari2600.pia.reset_timer[6] ));
 sg13g2_dfrbp_1 _28521_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1969),
    .D(_00906_),
    .Q_N(_13103_),
    .Q(\atari2600.pia.reset_timer[7] ));
 sg13g2_dfrbp_1 _28522_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1968),
    .D(_00907_),
    .Q_N(_13102_),
    .Q(\atari2600.pia.swa_dir[0] ));
 sg13g2_dfrbp_1 _28523_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1967),
    .D(_00908_),
    .Q_N(_13101_),
    .Q(\atari2600.pia.swa_dir[1] ));
 sg13g2_dfrbp_1 _28524_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1966),
    .D(_00909_),
    .Q_N(_13100_),
    .Q(\atari2600.pia.swa_dir[2] ));
 sg13g2_dfrbp_1 _28525_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1965),
    .D(_00910_),
    .Q_N(_13099_),
    .Q(\atari2600.pia.swa_dir[3] ));
 sg13g2_dfrbp_1 _28526_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1964),
    .D(_00911_),
    .Q_N(_13098_),
    .Q(\atari2600.pia.swa_dir[4] ));
 sg13g2_dfrbp_1 _28527_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1963),
    .D(_00912_),
    .Q_N(_13097_),
    .Q(\atari2600.pia.swa_dir[5] ));
 sg13g2_dfrbp_1 _28528_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1962),
    .D(_00913_),
    .Q_N(_13096_),
    .Q(\atari2600.pia.swa_dir[6] ));
 sg13g2_dfrbp_1 _28529_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1961),
    .D(_00914_),
    .Q_N(_13095_),
    .Q(\atari2600.pia.swa_dir[7] ));
 sg13g2_dfrbp_1 _28530_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1960),
    .D(net7041),
    .Q_N(_13094_),
    .Q(\atari2600.tia.old_grp1[0] ));
 sg13g2_dfrbp_1 _28531_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1959),
    .D(net6765),
    .Q_N(_13093_),
    .Q(\atari2600.tia.old_grp1[1] ));
 sg13g2_dfrbp_1 _28532_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1958),
    .D(net7140),
    .Q_N(_13092_),
    .Q(\atari2600.tia.old_grp1[2] ));
 sg13g2_dfrbp_1 _28533_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1957),
    .D(net4942),
    .Q_N(_13091_),
    .Q(\atari2600.tia.old_grp1[3] ));
 sg13g2_dfrbp_1 _28534_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1956),
    .D(net4526),
    .Q_N(_13090_),
    .Q(\atari2600.tia.old_grp1[4] ));
 sg13g2_dfrbp_1 _28535_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1955),
    .D(net4347),
    .Q_N(_13089_),
    .Q(\atari2600.tia.old_grp1[5] ));
 sg13g2_dfrbp_1 _28536_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1954),
    .D(net4705),
    .Q_N(_13088_),
    .Q(\atari2600.tia.old_grp1[6] ));
 sg13g2_dfrbp_1 _28537_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1953),
    .D(net4575),
    .Q_N(_13087_),
    .Q(\atari2600.tia.old_grp1[7] ));
 sg13g2_dfrbp_1 _28538_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1952),
    .D(_00923_),
    .Q_N(_13086_),
    .Q(\atari2600.tia.p0_spacing[4] ));
 sg13g2_dfrbp_1 _28539_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1950),
    .D(_00924_),
    .Q_N(_13085_),
    .Q(\atari2600.tia.p0_spacing[5] ));
 sg13g2_dfrbp_1 _28540_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1948),
    .D(_00925_),
    .Q_N(_13084_),
    .Q(\atari2600.tia.p0_spacing[6] ));
 sg13g2_dfrbp_1 _28541_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1946),
    .D(_00926_),
    .Q_N(_13083_),
    .Q(\atari2600.tia.p1_w[3] ));
 sg13g2_dfrbp_1 _28542_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1944),
    .D(_00927_),
    .Q_N(_13082_),
    .Q(\atari2600.tia.p1_w[4] ));
 sg13g2_dfrbp_1 _28543_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1943),
    .D(_00928_),
    .Q_N(_13081_),
    .Q(\atari2600.tia.p1_w[5] ));
 sg13g2_dfrbp_1 _28544_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1942),
    .D(_00929_),
    .Q_N(_13080_),
    .Q(\atari2600.tia.p1_scale[0] ));
 sg13g2_dfrbp_1 _28545_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1941),
    .D(_00930_),
    .Q_N(_13079_),
    .Q(\atari2600.tia.p1_scale[1] ));
 sg13g2_dfrbp_1 _28546_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1940),
    .D(_00931_),
    .Q_N(_13078_),
    .Q(\atari2600.tia.p0_scale[0] ));
 sg13g2_dfrbp_1 _28547_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1939),
    .D(_00932_),
    .Q_N(_13077_),
    .Q(\atari2600.tia.p0_scale[1] ));
 sg13g2_dfrbp_1 _28548_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1938),
    .D(_00933_),
    .Q_N(_13076_),
    .Q(\atari2600.tia.p0_w[3] ));
 sg13g2_dfrbp_1 _28549_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1937),
    .D(_00934_),
    .Q_N(_13075_),
    .Q(\atari2600.tia.p0_w[4] ));
 sg13g2_dfrbp_1 _28550_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1936),
    .D(_00935_),
    .Q_N(_13074_),
    .Q(\atari2600.tia.p0_w[5] ));
 sg13g2_dfrbp_1 _28551_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1935),
    .D(_00936_),
    .Q_N(_13073_),
    .Q(\atari2600.pia.interval[3] ));
 sg13g2_dfrbp_1 _28552_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1934),
    .D(_00937_),
    .Q_N(_13072_),
    .Q(\atari2600.pia.interval[6] ));
 sg13g2_dfrbp_1 _28553_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1933),
    .D(_00938_),
    .Q_N(_13071_),
    .Q(\atari2600.pia.interval[10] ));
 sg13g2_dfrbp_1 _28554_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1932),
    .D(_00939_),
    .Q_N(_13070_),
    .Q(\atari2600.tia.m1_w[0] ));
 sg13g2_dfrbp_1 _28555_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1931),
    .D(_00940_),
    .Q_N(_13069_),
    .Q(\atari2600.tia.m1_w[1] ));
 sg13g2_dfrbp_1 _28556_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1930),
    .D(_00941_),
    .Q_N(_13068_),
    .Q(\atari2600.tia.m1_w[2] ));
 sg13g2_dfrbp_1 _28557_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1929),
    .D(_00942_),
    .Q_N(_13067_),
    .Q(\atari2600.tia.m1_w[3] ));
 sg13g2_dfrbp_1 _28558_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1928),
    .D(_00943_),
    .Q_N(_13066_),
    .Q(\atari2600.tia.m0_w[0] ));
 sg13g2_dfrbp_1 _28559_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1927),
    .D(_00944_),
    .Q_N(_13065_),
    .Q(\atari2600.tia.m0_w[1] ));
 sg13g2_dfrbp_1 _28560_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1926),
    .D(_00945_),
    .Q_N(_13064_),
    .Q(\atari2600.tia.m0_w[2] ));
 sg13g2_dfrbp_1 _28561_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1925),
    .D(_00946_),
    .Q_N(_13063_),
    .Q(\atari2600.tia.m0_w[3] ));
 sg13g2_dfrbp_1 _28562_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1924),
    .D(_00947_),
    .Q_N(_13062_),
    .Q(\atari2600.tia.ball_w[0] ));
 sg13g2_dfrbp_1 _28563_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1923),
    .D(_00948_),
    .Q_N(_13061_),
    .Q(\atari2600.tia.ball_w[1] ));
 sg13g2_dfrbp_1 _28564_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1922),
    .D(_00949_),
    .Q_N(_13060_),
    .Q(\atari2600.tia.ball_w[2] ));
 sg13g2_dfrbp_1 _28565_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1921),
    .D(_00950_),
    .Q_N(_13059_),
    .Q(\atari2600.tia.ball_w[3] ));
 sg13g2_dfrbp_1 _28566_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1920),
    .D(_00951_),
    .Q_N(_13058_),
    .Q(\flash_rom.addr[0] ));
 sg13g2_dfrbp_1 _28567_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1919),
    .D(_00952_),
    .Q_N(_13057_),
    .Q(\flash_rom.addr[1] ));
 sg13g2_dfrbp_1 _28568_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1918),
    .D(_00953_),
    .Q_N(_13056_),
    .Q(\flash_rom.addr[2] ));
 sg13g2_dfrbp_1 _28569_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1917),
    .D(_00954_),
    .Q_N(_13055_),
    .Q(\flash_rom.addr[3] ));
 sg13g2_dfrbp_1 _28570_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1916),
    .D(_00955_),
    .Q_N(_13054_),
    .Q(\flash_rom.addr[4] ));
 sg13g2_dfrbp_1 _28571_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1915),
    .D(_00956_),
    .Q_N(_13053_),
    .Q(\flash_rom.addr[5] ));
 sg13g2_dfrbp_1 _28572_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1914),
    .D(_00957_),
    .Q_N(_13052_),
    .Q(\flash_rom.addr[6] ));
 sg13g2_dfrbp_1 _28573_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1913),
    .D(_00958_),
    .Q_N(_13051_),
    .Q(\flash_rom.addr[7] ));
 sg13g2_dfrbp_1 _28574_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1912),
    .D(_00959_),
    .Q_N(_13050_),
    .Q(\flash_rom.addr[8] ));
 sg13g2_dfrbp_1 _28575_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1911),
    .D(_00960_),
    .Q_N(_13049_),
    .Q(\flash_rom.addr[9] ));
 sg13g2_dfrbp_1 _28576_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1910),
    .D(_00961_),
    .Q_N(_13048_),
    .Q(\flash_rom.addr[10] ));
 sg13g2_dfrbp_1 _28577_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1909),
    .D(_00962_),
    .Q_N(_13047_),
    .Q(\flash_rom.addr[11] ));
 sg13g2_dfrbp_1 _28578_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1908),
    .D(net2995),
    .Q_N(_13046_),
    .Q(\flash_rom.addr[16] ));
 sg13g2_dfrbp_1 _28579_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1907),
    .D(net4518),
    .Q_N(_13045_),
    .Q(\flash_rom.addr[17] ));
 sg13g2_dfrbp_1 _28580_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1906),
    .D(net7195),
    .Q_N(_13044_),
    .Q(\flash_rom.addr[18] ));
 sg13g2_dfrbp_1 _28581_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1905),
    .D(net4426),
    .Q_N(_13043_),
    .Q(\flash_rom.addr[19] ));
 sg13g2_dfrbp_1 _28582_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1904),
    .D(_00967_),
    .Q_N(_13042_),
    .Q(\atari2600.ram[53][0] ));
 sg13g2_dfrbp_1 _28583_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1903),
    .D(_00968_),
    .Q_N(_13041_),
    .Q(\atari2600.ram[53][1] ));
 sg13g2_dfrbp_1 _28584_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1902),
    .D(_00969_),
    .Q_N(_13040_),
    .Q(\atari2600.ram[53][2] ));
 sg13g2_dfrbp_1 _28585_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1901),
    .D(_00970_),
    .Q_N(_13039_),
    .Q(\atari2600.ram[53][3] ));
 sg13g2_dfrbp_1 _28586_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1900),
    .D(_00971_),
    .Q_N(_13038_),
    .Q(\atari2600.ram[53][4] ));
 sg13g2_dfrbp_1 _28587_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1899),
    .D(_00972_),
    .Q_N(_13037_),
    .Q(\atari2600.ram[53][5] ));
 sg13g2_dfrbp_1 _28588_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1898),
    .D(_00973_),
    .Q_N(_13036_),
    .Q(\atari2600.ram[53][6] ));
 sg13g2_dfrbp_1 _28589_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1897),
    .D(_00974_),
    .Q_N(_13035_),
    .Q(\atari2600.ram[53][7] ));
 sg13g2_dfrbp_1 _28590_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1896),
    .D(net2990),
    .Q_N(_13034_),
    .Q(\flash_rom.addr[12] ));
 sg13g2_dfrbp_1 _28591_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1895),
    .D(net3257),
    .Q_N(_13033_),
    .Q(\flash_rom.addr[13] ));
 sg13g2_dfrbp_1 _28592_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1894),
    .D(net3050),
    .Q_N(_13032_),
    .Q(\flash_rom.addr[14] ));
 sg13g2_dfrbp_1 _28593_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1893),
    .D(net3215),
    .Q_N(_13031_),
    .Q(\flash_rom.addr[15] ));
 sg13g2_dfrbp_1 _28594_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1892),
    .D(net7237),
    .Q_N(_13030_),
    .Q(\flash_rom.addr[20] ));
 sg13g2_dfrbp_1 _28595_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1891),
    .D(net3940),
    .Q_N(_13029_),
    .Q(\flash_rom.addr[21] ));
 sg13g2_dfrbp_1 _28596_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1890),
    .D(net4434),
    .Q_N(_13028_),
    .Q(\flash_rom.addr[22] ));
 sg13g2_dfrbp_1 _28597_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1889),
    .D(net3747),
    .Q_N(_13027_),
    .Q(\flash_rom.addr[23] ));
 sg13g2_dfrbp_1 _28598_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1888),
    .D(_00983_),
    .Q_N(_13026_),
    .Q(\atari2600.ram[30][0] ));
 sg13g2_dfrbp_1 _28599_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1887),
    .D(_00984_),
    .Q_N(_13025_),
    .Q(\atari2600.ram[30][1] ));
 sg13g2_dfrbp_1 _28600_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1886),
    .D(_00985_),
    .Q_N(_13024_),
    .Q(\atari2600.ram[30][2] ));
 sg13g2_dfrbp_1 _28601_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1885),
    .D(_00986_),
    .Q_N(_13023_),
    .Q(\atari2600.ram[30][3] ));
 sg13g2_dfrbp_1 _28602_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1884),
    .D(_00987_),
    .Q_N(_13022_),
    .Q(\atari2600.ram[30][4] ));
 sg13g2_dfrbp_1 _28603_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1883),
    .D(_00988_),
    .Q_N(_13021_),
    .Q(\atari2600.ram[30][5] ));
 sg13g2_dfrbp_1 _28604_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1882),
    .D(_00989_),
    .Q_N(_13020_),
    .Q(\atari2600.ram[30][6] ));
 sg13g2_dfrbp_1 _28605_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1881),
    .D(_00990_),
    .Q_N(_13019_),
    .Q(\atari2600.ram[30][7] ));
 sg13g2_dfrbp_1 _28606_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1880),
    .D(net4539),
    .Q_N(_00095_),
    .Q(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_dfrbp_1 _28607_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1879),
    .D(net7307),
    .Q_N(_13018_),
    .Q(\atari2600.tia.audio_left_counter[1] ));
 sg13g2_dfrbp_1 _28608_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1878),
    .D(net3399),
    .Q_N(_00097_),
    .Q(\atari2600.tia.audio_left_counter[2] ));
 sg13g2_dfrbp_1 _28609_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1877),
    .D(net3020),
    .Q_N(_00098_),
    .Q(\atari2600.tia.audio_left_counter[3] ));
 sg13g2_dfrbp_1 _28610_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1876),
    .D(net3255),
    .Q_N(_00099_),
    .Q(\atari2600.tia.audio_left_counter[4] ));
 sg13g2_dfrbp_1 _28611_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1875),
    .D(net3107),
    .Q_N(_00100_),
    .Q(\atari2600.tia.audio_left_counter[5] ));
 sg13g2_dfrbp_1 _28612_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1874),
    .D(net3138),
    .Q_N(_00102_),
    .Q(\atari2600.tia.audio_left_counter[6] ));
 sg13g2_dfrbp_1 _28613_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1873),
    .D(net3263),
    .Q_N(_00103_),
    .Q(\atari2600.tia.audio_left_counter[7] ));
 sg13g2_dfrbp_1 _28614_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1872),
    .D(net3829),
    .Q_N(_00104_),
    .Q(\atari2600.tia.audio_left_counter[8] ));
 sg13g2_dfrbp_1 _28615_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1871),
    .D(net3119),
    .Q_N(_00105_),
    .Q(\atari2600.tia.audio_left_counter[9] ));
 sg13g2_dfrbp_1 _28616_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1870),
    .D(net3778),
    .Q_N(_00106_),
    .Q(\atari2600.tia.audio_left_counter[10] ));
 sg13g2_dfrbp_1 _28617_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1869),
    .D(net2987),
    .Q_N(_00107_),
    .Q(\atari2600.tia.audio_left_counter[11] ));
 sg13g2_dfrbp_1 _28618_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1868),
    .D(net3606),
    .Q_N(_00108_),
    .Q(\atari2600.tia.audio_left_counter[12] ));
 sg13g2_dfrbp_1 _28619_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1867),
    .D(net3213),
    .Q_N(_00109_),
    .Q(\atari2600.tia.audio_left_counter[13] ));
 sg13g2_dfrbp_1 _28620_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1866),
    .D(net2966),
    .Q_N(_00110_),
    .Q(\atari2600.tia.audio_left_counter[14] ));
 sg13g2_dfrbp_1 _28621_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1865),
    .D(net2953),
    .Q_N(_00111_),
    .Q(\atari2600.tia.audio_left_counter[15] ));
 sg13g2_dfrbp_1 _28622_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1864),
    .D(net7352),
    .Q_N(_00156_),
    .Q(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_dfrbp_1 _28623_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1863),
    .D(net7310),
    .Q_N(_13017_),
    .Q(\atari2600.tia.audio_right_counter[1] ));
 sg13g2_dfrbp_1 _28624_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1862),
    .D(net4211),
    .Q_N(_00113_),
    .Q(\atari2600.tia.audio_right_counter[2] ));
 sg13g2_dfrbp_1 _28625_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1861),
    .D(net3092),
    .Q_N(_00114_),
    .Q(\atari2600.tia.audio_right_counter[3] ));
 sg13g2_dfrbp_1 _28626_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1860),
    .D(net3364),
    .Q_N(_00115_),
    .Q(\atari2600.tia.audio_right_counter[4] ));
 sg13g2_dfrbp_1 _28627_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1859),
    .D(net3028),
    .Q_N(_00116_),
    .Q(\atari2600.tia.audio_right_counter[5] ));
 sg13g2_dfrbp_1 _28628_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1858),
    .D(net3800),
    .Q_N(_00117_),
    .Q(\atari2600.tia.audio_right_counter[6] ));
 sg13g2_dfrbp_1 _28629_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1857),
    .D(net2958),
    .Q_N(_00118_),
    .Q(\atari2600.tia.audio_right_counter[7] ));
 sg13g2_dfrbp_1 _28630_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1856),
    .D(net3044),
    .Q_N(_00119_),
    .Q(\atari2600.tia.audio_right_counter[8] ));
 sg13g2_dfrbp_1 _28631_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1855),
    .D(net2997),
    .Q_N(_00120_),
    .Q(\atari2600.tia.audio_right_counter[9] ));
 sg13g2_dfrbp_1 _28632_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1854),
    .D(net3844),
    .Q_N(_00121_),
    .Q(\atari2600.tia.audio_right_counter[10] ));
 sg13g2_dfrbp_1 _28633_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1853),
    .D(net3003),
    .Q_N(_00122_),
    .Q(\atari2600.tia.audio_right_counter[11] ));
 sg13g2_dfrbp_1 _28634_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1852),
    .D(net3176),
    .Q_N(_00123_),
    .Q(\atari2600.tia.audio_right_counter[12] ));
 sg13g2_dfrbp_1 _28635_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1851),
    .D(net2975),
    .Q_N(_00124_),
    .Q(\atari2600.tia.audio_right_counter[13] ));
 sg13g2_dfrbp_1 _28636_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1850),
    .D(net3012),
    .Q_N(_00125_),
    .Q(\atari2600.tia.audio_right_counter[14] ));
 sg13g2_dfrbp_1 _28637_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1849),
    .D(net2944),
    .Q_N(_00126_),
    .Q(\atari2600.tia.audio_right_counter[15] ));
 sg13g2_dfrbp_1 _28638_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1847),
    .D(net7462),
    .Q_N(_00155_),
    .Q(\atari2600.tia.audio_l ));
 sg13g2_dfrbp_1 _28639_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1845),
    .D(_01024_),
    .Q_N(_00154_),
    .Q(\atari2600.tia.audio_r ));
 sg13g2_dfrbp_1 _28640_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net806),
    .D(_01025_),
    .Q_N(_13843_),
    .Q(\atari2600.tia.vid_vsync ));
 sg13g2_dfrbp_1 _28641_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net807),
    .D(_00038_),
    .Q_N(_00153_),
    .Q(\atari2600.tia.vid_xpos[0] ));
 sg13g2_dfrbp_1 _28642_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net808),
    .D(_00039_),
    .Q_N(_00152_),
    .Q(\atari2600.tia.vid_xpos[1] ));
 sg13g2_dfrbp_1 _28643_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net809),
    .D(_00040_),
    .Q_N(_00140_),
    .Q(\atari2600.tia.vid_xpos[2] ));
 sg13g2_dfrbp_1 _28644_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net810),
    .D(_00041_),
    .Q_N(_00141_),
    .Q(\atari2600.tia.vid_xpos[3] ));
 sg13g2_dfrbp_1 _28645_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net811),
    .D(_00042_),
    .Q_N(_00145_),
    .Q(\atari2600.tia.vid_xpos[4] ));
 sg13g2_dfrbp_1 _28646_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net812),
    .D(_00043_),
    .Q_N(_00142_),
    .Q(\atari2600.tia.vid_xpos[5] ));
 sg13g2_dfrbp_1 _28647_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net813),
    .D(_00044_),
    .Q_N(_00143_),
    .Q(\atari2600.tia.vid_xpos[6] ));
 sg13g2_dfrbp_1 _28648_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net814),
    .D(_00045_),
    .Q_N(_00139_),
    .Q(\atari2600.tia.vid_xpos[7] ));
 sg13g2_dfrbp_1 _28649_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net815),
    .D(_00046_),
    .Q_N(_00157_),
    .Q(\atari2600.tia.vid_ypos[0] ));
 sg13g2_dfrbp_1 _28650_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net816),
    .D(net2950),
    .Q_N(_00158_),
    .Q(\atari2600.tia.vid_ypos[1] ));
 sg13g2_dfrbp_1 _28651_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net817),
    .D(net3115),
    .Q_N(_00159_),
    .Q(\atari2600.tia.vid_ypos[2] ));
 sg13g2_dfrbp_1 _28652_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net818),
    .D(_00049_),
    .Q_N(_00131_),
    .Q(\atari2600.tia.vid_ypos[3] ));
 sg13g2_dfrbp_1 _28653_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net819),
    .D(_00050_),
    .Q_N(_00160_),
    .Q(\atari2600.tia.vid_ypos[4] ));
 sg13g2_dfrbp_1 _28654_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net820),
    .D(net3457),
    .Q_N(_00070_),
    .Q(\atari2600.tia.vid_ypos[5] ));
 sg13g2_dfrbp_1 _28655_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net821),
    .D(_00052_),
    .Q_N(_00161_),
    .Q(\atari2600.tia.vid_ypos[6] ));
 sg13g2_dfrbp_1 _28656_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net964),
    .D(net2964),
    .Q_N(_00162_),
    .Q(\atari2600.tia.vid_ypos[7] ));
 sg13g2_dfrbp_1 _28657_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1843),
    .D(_00054_),
    .Q_N(_00130_),
    .Q(\atari2600.tia.vid_ypos[8] ));
 sg13g2_dfrbp_1 _28658_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1841),
    .D(_01026_),
    .Q_N(_13016_),
    .Q(\atari2600.tia.vblank ));
 sg13g2_dfrbp_1 _28659_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1839),
    .D(_01027_),
    .Q_N(_13015_),
    .Q(\atari2600.stall_cpu ));
 sg13g2_dfrbp_1 _28660_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1837),
    .D(_01028_),
    .Q_N(_13014_),
    .Q(\atari2600.pia.swb_dir[2] ));
 sg13g2_dfrbp_1 _28661_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1836),
    .D(_01029_),
    .Q_N(_13013_),
    .Q(\atari2600.pia.swb_dir[4] ));
 sg13g2_dfrbp_1 _28662_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1835),
    .D(_01030_),
    .Q_N(_13012_),
    .Q(\atari2600.pia.swb_dir[5] ));
 sg13g2_dfrbp_1 _28663_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1834),
    .D(_01031_),
    .Q_N(_13011_),
    .Q(\atari2600.tia.colubk[0] ));
 sg13g2_dfrbp_1 _28664_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1832),
    .D(_01032_),
    .Q_N(_13010_),
    .Q(\atari2600.tia.colubk[1] ));
 sg13g2_dfrbp_1 _28665_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1831),
    .D(_01033_),
    .Q_N(_13009_),
    .Q(\atari2600.tia.colubk[2] ));
 sg13g2_dfrbp_1 _28666_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1830),
    .D(_01034_),
    .Q_N(_13008_),
    .Q(\atari2600.tia.colubk[3] ));
 sg13g2_dfrbp_1 _28667_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1829),
    .D(_01035_),
    .Q_N(_13007_),
    .Q(\atari2600.tia.colubk[4] ));
 sg13g2_dfrbp_1 _28668_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1828),
    .D(_01036_),
    .Q_N(_13006_),
    .Q(\atari2600.tia.colubk[5] ));
 sg13g2_dfrbp_1 _28669_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1827),
    .D(_01037_),
    .Q_N(_13005_),
    .Q(\atari2600.tia.colubk[6] ));
 sg13g2_dfrbp_1 _28670_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1826),
    .D(_01038_),
    .Q_N(_13004_),
    .Q(\atari2600.tia.colup0[0] ));
 sg13g2_dfrbp_1 _28671_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1825),
    .D(_01039_),
    .Q_N(_13003_),
    .Q(\atari2600.tia.colup0[1] ));
 sg13g2_dfrbp_1 _28672_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1824),
    .D(_01040_),
    .Q_N(_13002_),
    .Q(\atari2600.tia.colup0[2] ));
 sg13g2_dfrbp_1 _28673_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1823),
    .D(_01041_),
    .Q_N(_13001_),
    .Q(\atari2600.tia.colup0[3] ));
 sg13g2_dfrbp_1 _28674_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1822),
    .D(_01042_),
    .Q_N(_13000_),
    .Q(\atari2600.tia.colup0[4] ));
 sg13g2_dfrbp_1 _28675_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1821),
    .D(_01043_),
    .Q_N(_12999_),
    .Q(\atari2600.tia.colup0[5] ));
 sg13g2_dfrbp_1 _28676_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1820),
    .D(_01044_),
    .Q_N(_12998_),
    .Q(\atari2600.tia.colup0[6] ));
 sg13g2_dfrbp_1 _28677_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1819),
    .D(_01045_),
    .Q_N(_12997_),
    .Q(\atari2600.tia.colup1[0] ));
 sg13g2_dfrbp_1 _28678_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1818),
    .D(_01046_),
    .Q_N(_12996_),
    .Q(\atari2600.tia.colup1[1] ));
 sg13g2_dfrbp_1 _28679_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1817),
    .D(_01047_),
    .Q_N(_12995_),
    .Q(\atari2600.tia.colup1[2] ));
 sg13g2_dfrbp_1 _28680_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1816),
    .D(_01048_),
    .Q_N(_12994_),
    .Q(\atari2600.tia.colup1[3] ));
 sg13g2_dfrbp_1 _28681_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1815),
    .D(_01049_),
    .Q_N(_12993_),
    .Q(\atari2600.tia.colup1[4] ));
 sg13g2_dfrbp_1 _28682_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1814),
    .D(_01050_),
    .Q_N(_12992_),
    .Q(\atari2600.tia.colup1[5] ));
 sg13g2_dfrbp_1 _28683_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1813),
    .D(_01051_),
    .Q_N(_12991_),
    .Q(\atari2600.tia.colup1[6] ));
 sg13g2_dfrbp_1 _28684_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1812),
    .D(_01052_),
    .Q_N(_12990_),
    .Q(\atari2600.tia.colupf[0] ));
 sg13g2_dfrbp_1 _28685_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1811),
    .D(_01053_),
    .Q_N(_12989_),
    .Q(\atari2600.tia.colupf[1] ));
 sg13g2_dfrbp_1 _28686_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1810),
    .D(_01054_),
    .Q_N(_12988_),
    .Q(\atari2600.tia.colupf[2] ));
 sg13g2_dfrbp_1 _28687_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1809),
    .D(_01055_),
    .Q_N(_12987_),
    .Q(\atari2600.tia.colupf[3] ));
 sg13g2_dfrbp_1 _28688_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1808),
    .D(_01056_),
    .Q_N(_12986_),
    .Q(\atari2600.tia.colupf[4] ));
 sg13g2_dfrbp_1 _28689_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1807),
    .D(_01057_),
    .Q_N(_12985_),
    .Q(\atari2600.tia.colupf[5] ));
 sg13g2_dfrbp_1 _28690_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1806),
    .D(_01058_),
    .Q_N(_12984_),
    .Q(\atari2600.tia.colupf[6] ));
 sg13g2_dfrbp_1 _28691_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1805),
    .D(_01059_),
    .Q_N(_12983_),
    .Q(\atari2600.tia.enam0 ));
 sg13g2_dfrbp_1 _28692_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1804),
    .D(_01060_),
    .Q_N(_12982_),
    .Q(\atari2600.tia.enam1 ));
 sg13g2_dfrbp_1 _28693_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1803),
    .D(_01061_),
    .Q_N(_12981_),
    .Q(\atari2600.tia.enabl ));
 sg13g2_dfrbp_1 _28694_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1802),
    .D(_01062_),
    .Q_N(_12980_),
    .Q(\atari2600.tia.vdelp0 ));
 sg13g2_dfrbp_1 _28695_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1801),
    .D(_01063_),
    .Q_N(_12979_),
    .Q(\atari2600.tia.vdelp1 ));
 sg13g2_dfrbp_1 _28696_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1800),
    .D(_01064_),
    .Q_N(_00151_),
    .Q(\atari2600.tia.refp0 ));
 sg13g2_dfrbp_1 _28697_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1799),
    .D(_01065_),
    .Q_N(_00148_),
    .Q(\atari2600.tia.refp1 ));
 sg13g2_dfrbp_1 _28698_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1798),
    .D(_01066_),
    .Q_N(_12978_),
    .Q(\atari2600.tia.refpf ));
 sg13g2_dfrbp_1 _28699_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1797),
    .D(_01067_),
    .Q_N(_12977_),
    .Q(\atari2600.tia.scorepf ));
 sg13g2_dfrbp_1 _28700_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1796),
    .D(_01068_),
    .Q_N(_12976_),
    .Q(\atari2600.tia.pf_priority ));
 sg13g2_dfrbp_1 _28701_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1795),
    .D(_01069_),
    .Q_N(_12975_),
    .Q(\atari2600.tia.diag[104] ));
 sg13g2_dfrbp_1 _28702_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1794),
    .D(_01070_),
    .Q_N(_12974_),
    .Q(\atari2600.tia.diag[105] ));
 sg13g2_dfrbp_1 _28703_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net1793),
    .D(_01071_),
    .Q_N(_12973_),
    .Q(\atari2600.tia.diag[106] ));
 sg13g2_dfrbp_1 _28704_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1792),
    .D(_01072_),
    .Q_N(_12972_),
    .Q(\atari2600.tia.diag[107] ));
 sg13g2_dfrbp_1 _28705_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1791),
    .D(_01073_),
    .Q_N(_12971_),
    .Q(\atari2600.tia.diag[108] ));
 sg13g2_dfrbp_1 _28706_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1790),
    .D(_01074_),
    .Q_N(_12970_),
    .Q(\atari2600.tia.diag[109] ));
 sg13g2_dfrbp_1 _28707_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1789),
    .D(_01075_),
    .Q_N(_12969_),
    .Q(\atari2600.tia.diag[110] ));
 sg13g2_dfrbp_1 _28708_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1788),
    .D(_01076_),
    .Q_N(_12968_),
    .Q(\atari2600.tia.diag[111] ));
 sg13g2_dfrbp_1 _28709_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1787),
    .D(_01077_),
    .Q_N(_12967_),
    .Q(\atari2600.tia.diag[96] ));
 sg13g2_dfrbp_1 _28710_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1786),
    .D(_01078_),
    .Q_N(_12966_),
    .Q(\atari2600.tia.diag[97] ));
 sg13g2_dfrbp_1 _28711_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1785),
    .D(_01079_),
    .Q_N(_12965_),
    .Q(\atari2600.tia.diag[98] ));
 sg13g2_dfrbp_1 _28712_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1784),
    .D(_01080_),
    .Q_N(_12964_),
    .Q(\atari2600.tia.diag[99] ));
 sg13g2_dfrbp_1 _28713_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1783),
    .D(_01081_),
    .Q_N(_12963_),
    .Q(\atari2600.tia.diag[100] ));
 sg13g2_dfrbp_1 _28714_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1782),
    .D(_01082_),
    .Q_N(_12962_),
    .Q(\atari2600.tia.diag[101] ));
 sg13g2_dfrbp_1 _28715_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1781),
    .D(_01083_),
    .Q_N(_12961_),
    .Q(\atari2600.tia.diag[102] ));
 sg13g2_dfrbp_1 _28716_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1780),
    .D(_01084_),
    .Q_N(_12960_),
    .Q(\atari2600.tia.diag[103] ));
 sg13g2_dfrbp_1 _28717_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1779),
    .D(_01085_),
    .Q_N(_12959_),
    .Q(\atari2600.tia.vid_out[0] ));
 sg13g2_dfrbp_1 _28718_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1778),
    .D(_01086_),
    .Q_N(_12958_),
    .Q(\atari2600.tia.vid_out[1] ));
 sg13g2_dfrbp_1 _28719_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1777),
    .D(_01087_),
    .Q_N(_12957_),
    .Q(\atari2600.tia.vid_out[2] ));
 sg13g2_dfrbp_1 _28720_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1776),
    .D(_01088_),
    .Q_N(_12956_),
    .Q(\atari2600.tia.vid_out[3] ));
 sg13g2_dfrbp_1 _28721_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1775),
    .D(_01089_),
    .Q_N(_12955_),
    .Q(\atari2600.tia.vid_out[4] ));
 sg13g2_dfrbp_1 _28722_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1774),
    .D(_01090_),
    .Q_N(_12954_),
    .Q(\atari2600.tia.vid_out[5] ));
 sg13g2_dfrbp_1 _28723_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1773),
    .D(_01091_),
    .Q_N(_12953_),
    .Q(\atari2600.tia.vid_out[6] ));
 sg13g2_dfrbp_1 _28724_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1772),
    .D(net3640),
    .Q_N(_12952_),
    .Q(\atari2600.tia.old_grp0[0] ));
 sg13g2_dfrbp_1 _28725_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1771),
    .D(net3919),
    .Q_N(_12951_),
    .Q(\atari2600.tia.old_grp0[1] ));
 sg13g2_dfrbp_1 _28726_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1770),
    .D(net3657),
    .Q_N(_12950_),
    .Q(\atari2600.tia.old_grp0[2] ));
 sg13g2_dfrbp_1 _28727_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1769),
    .D(net3813),
    .Q_N(_12949_),
    .Q(\atari2600.tia.old_grp0[3] ));
 sg13g2_dfrbp_1 _28728_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1768),
    .D(net3666),
    .Q_N(_12948_),
    .Q(\atari2600.tia.old_grp0[4] ));
 sg13g2_dfrbp_1 _28729_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1767),
    .D(net4190),
    .Q_N(_12947_),
    .Q(\atari2600.tia.old_grp0[5] ));
 sg13g2_dfrbp_1 _28730_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1766),
    .D(net3534),
    .Q_N(_12946_),
    .Q(\atari2600.tia.old_grp0[6] ));
 sg13g2_dfrbp_1 _28731_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1765),
    .D(net3537),
    .Q_N(_12945_),
    .Q(\atari2600.tia.old_grp0[7] ));
 sg13g2_dfrbp_1 _28732_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1764),
    .D(net7482),
    .Q_N(_12944_),
    .Q(\atari2600.tia.diag[64] ));
 sg13g2_dfrbp_1 _28733_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1763),
    .D(net7537),
    .Q_N(_12943_),
    .Q(\atari2600.tia.diag[65] ));
 sg13g2_dfrbp_1 _28734_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1762),
    .D(_01102_),
    .Q_N(_12942_),
    .Q(\atari2600.tia.diag[66] ));
 sg13g2_dfrbp_1 _28735_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1761),
    .D(_01103_),
    .Q_N(_12941_),
    .Q(\atari2600.tia.diag[67] ));
 sg13g2_dfrbp_1 _28736_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1760),
    .D(_01104_),
    .Q_N(_12940_),
    .Q(\atari2600.tia.diag[68] ));
 sg13g2_dfrbp_1 _28737_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1759),
    .D(_01105_),
    .Q_N(_00150_),
    .Q(\atari2600.tia.diag[69] ));
 sg13g2_dfrbp_1 _28738_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1758),
    .D(_01106_),
    .Q_N(_00149_),
    .Q(\atari2600.tia.diag[70] ));
 sg13g2_dfrbp_1 _28739_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1757),
    .D(_01107_),
    .Q_N(_12939_),
    .Q(\atari2600.tia.diag[71] ));
 sg13g2_dfrbp_1 _28740_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1756),
    .D(_01108_),
    .Q_N(_12938_),
    .Q(\atari2600.tia.diag[56] ));
 sg13g2_dfrbp_1 _28741_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1755),
    .D(_01109_),
    .Q_N(_12937_),
    .Q(\atari2600.tia.diag[57] ));
 sg13g2_dfrbp_1 _28742_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1754),
    .D(_01110_),
    .Q_N(_12936_),
    .Q(\atari2600.tia.diag[58] ));
 sg13g2_dfrbp_1 _28743_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1752),
    .D(_01111_),
    .Q_N(_12935_),
    .Q(\atari2600.tia.diag[59] ));
 sg13g2_dfrbp_1 _28744_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1750),
    .D(_01112_),
    .Q_N(_12934_),
    .Q(\atari2600.tia.diag[60] ));
 sg13g2_dfrbp_1 _28745_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1748),
    .D(_01113_),
    .Q_N(_00146_),
    .Q(\atari2600.tia.diag[61] ));
 sg13g2_dfrbp_1 _28746_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1746),
    .D(_01114_),
    .Q_N(_00144_),
    .Q(\atari2600.tia.diag[62] ));
 sg13g2_dfrbp_1 _28747_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1744),
    .D(_01115_),
    .Q_N(_00147_),
    .Q(\atari2600.tia.diag[63] ));
 sg13g2_dfrbp_1 _28748_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1742),
    .D(_01116_),
    .Q_N(_12933_),
    .Q(\atari2600.tia.diag[48] ));
 sg13g2_dfrbp_1 _28749_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1740),
    .D(_01117_),
    .Q_N(_12932_),
    .Q(\atari2600.tia.diag[49] ));
 sg13g2_dfrbp_1 _28750_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1739),
    .D(net7521),
    .Q_N(_12931_),
    .Q(\atari2600.tia.diag[50] ));
 sg13g2_dfrbp_1 _28751_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1738),
    .D(_01119_),
    .Q_N(_12930_),
    .Q(\atari2600.tia.diag[51] ));
 sg13g2_dfrbp_1 _28752_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1737),
    .D(net7511),
    .Q_N(_12929_),
    .Q(\atari2600.tia.diag[52] ));
 sg13g2_dfrbp_1 _28753_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1736),
    .D(_01121_),
    .Q_N(_12928_),
    .Q(\atari2600.tia.diag[53] ));
 sg13g2_dfrbp_1 _28754_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1735),
    .D(_01122_),
    .Q_N(_12927_),
    .Q(\atari2600.tia.diag[54] ));
 sg13g2_dfrbp_1 _28755_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1734),
    .D(_01123_),
    .Q_N(_12926_),
    .Q(\atari2600.tia.diag[55] ));
 sg13g2_dfrbp_1 _28756_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1733),
    .D(_01124_),
    .Q_N(_12925_),
    .Q(\atari2600.tia.diag[40] ));
 sg13g2_dfrbp_1 _28757_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1732),
    .D(net7573),
    .Q_N(_12924_),
    .Q(\atari2600.tia.diag[41] ));
 sg13g2_dfrbp_1 _28758_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1731),
    .D(_01126_),
    .Q_N(_12923_),
    .Q(\atari2600.tia.diag[42] ));
 sg13g2_dfrbp_1 _28759_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1730),
    .D(_01127_),
    .Q_N(_12922_),
    .Q(\atari2600.tia.diag[43] ));
 sg13g2_dfrbp_1 _28760_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1729),
    .D(_01128_),
    .Q_N(_12921_),
    .Q(\atari2600.tia.diag[44] ));
 sg13g2_dfrbp_1 _28761_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1728),
    .D(_01129_),
    .Q_N(_12920_),
    .Q(\atari2600.tia.diag[45] ));
 sg13g2_dfrbp_1 _28762_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1727),
    .D(_01130_),
    .Q_N(_12919_),
    .Q(\atari2600.tia.diag[46] ));
 sg13g2_dfrbp_1 _28763_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1726),
    .D(net7493),
    .Q_N(_12918_),
    .Q(\atari2600.tia.diag[47] ));
 sg13g2_dfrbp_1 _28764_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1725),
    .D(_01132_),
    .Q_N(_12917_),
    .Q(\atari2600.tia.diag[32] ));
 sg13g2_dfrbp_1 _28765_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1724),
    .D(net7568),
    .Q_N(_12916_),
    .Q(\atari2600.tia.diag[33] ));
 sg13g2_dfrbp_1 _28766_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1723),
    .D(_01134_),
    .Q_N(_12915_),
    .Q(\atari2600.tia.diag[34] ));
 sg13g2_dfrbp_1 _28767_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1722),
    .D(_01135_),
    .Q_N(_12914_),
    .Q(\atari2600.tia.diag[35] ));
 sg13g2_dfrbp_1 _28768_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1721),
    .D(_01136_),
    .Q_N(_12913_),
    .Q(\atari2600.tia.diag[36] ));
 sg13g2_dfrbp_1 _28769_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1720),
    .D(_01137_),
    .Q_N(_12912_),
    .Q(\atari2600.tia.diag[37] ));
 sg13g2_dfrbp_1 _28770_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1719),
    .D(_01138_),
    .Q_N(_12911_),
    .Q(\atari2600.tia.diag[38] ));
 sg13g2_dfrbp_1 _28771_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1718),
    .D(_01139_),
    .Q_N(_12910_),
    .Q(\atari2600.tia.diag[39] ));
 sg13g2_dfrbp_1 _28772_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1717),
    .D(_01140_),
    .Q_N(_12909_),
    .Q(\atari2600.tia.diag[88] ));
 sg13g2_dfrbp_1 _28773_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1716),
    .D(_01141_),
    .Q_N(_12908_),
    .Q(\atari2600.tia.diag[89] ));
 sg13g2_dfrbp_1 _28774_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1715),
    .D(_01142_),
    .Q_N(_12907_),
    .Q(\atari2600.tia.diag[90] ));
 sg13g2_dfrbp_1 _28775_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1714),
    .D(_01143_),
    .Q_N(_12906_),
    .Q(\atari2600.tia.diag[91] ));
 sg13g2_dfrbp_1 _28776_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1713),
    .D(_01144_),
    .Q_N(_12905_),
    .Q(\atari2600.tia.diag[92] ));
 sg13g2_dfrbp_1 _28777_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1712),
    .D(_01145_),
    .Q_N(_12904_),
    .Q(\atari2600.tia.diag[93] ));
 sg13g2_dfrbp_1 _28778_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1711),
    .D(_01146_),
    .Q_N(_12903_),
    .Q(\atari2600.tia.diag[94] ));
 sg13g2_dfrbp_1 _28779_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1710),
    .D(_01147_),
    .Q_N(_12902_),
    .Q(\atari2600.tia.diag[95] ));
 sg13g2_dfrbp_1 _28780_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1709),
    .D(_01148_),
    .Q_N(_12901_),
    .Q(\atari2600.tia.hmp0[0] ));
 sg13g2_dfrbp_1 _28781_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1708),
    .D(_01149_),
    .Q_N(_12900_),
    .Q(\atari2600.tia.hmp0[1] ));
 sg13g2_dfrbp_1 _28782_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1707),
    .D(_01150_),
    .Q_N(_12899_),
    .Q(\atari2600.tia.hmp0[2] ));
 sg13g2_dfrbp_1 _28783_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1706),
    .D(_01151_),
    .Q_N(_12898_),
    .Q(\atari2600.tia.hmp0[3] ));
 sg13g2_dfrbp_1 _28784_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1705),
    .D(_01152_),
    .Q_N(_12897_),
    .Q(\atari2600.tia.hmp1[0] ));
 sg13g2_dfrbp_1 _28785_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1704),
    .D(_01153_),
    .Q_N(_12896_),
    .Q(\atari2600.tia.hmp1[1] ));
 sg13g2_dfrbp_1 _28786_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1703),
    .D(_01154_),
    .Q_N(_12895_),
    .Q(\atari2600.tia.hmp1[2] ));
 sg13g2_dfrbp_1 _28787_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1702),
    .D(_01155_),
    .Q_N(_12894_),
    .Q(\atari2600.tia.hmp1[3] ));
 sg13g2_dfrbp_1 _28788_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1701),
    .D(_01156_),
    .Q_N(_12893_),
    .Q(\atari2600.tia.hmm0[0] ));
 sg13g2_dfrbp_1 _28789_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1700),
    .D(_01157_),
    .Q_N(_12892_),
    .Q(\atari2600.tia.hmm0[1] ));
 sg13g2_dfrbp_1 _28790_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1699),
    .D(_01158_),
    .Q_N(_12891_),
    .Q(\atari2600.tia.hmm0[2] ));
 sg13g2_dfrbp_1 _28791_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1698),
    .D(_01159_),
    .Q_N(_12890_),
    .Q(\atari2600.tia.hmm0[3] ));
 sg13g2_dfrbp_1 _28792_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1697),
    .D(_01160_),
    .Q_N(_12889_),
    .Q(\atari2600.tia.hmm1[0] ));
 sg13g2_dfrbp_1 _28793_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1696),
    .D(_01161_),
    .Q_N(_12888_),
    .Q(\atari2600.tia.hmm1[1] ));
 sg13g2_dfrbp_1 _28794_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1695),
    .D(_01162_),
    .Q_N(_12887_),
    .Q(\atari2600.tia.hmm1[2] ));
 sg13g2_dfrbp_1 _28795_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1694),
    .D(_01163_),
    .Q_N(_12886_),
    .Q(\atari2600.tia.hmm1[3] ));
 sg13g2_dfrbp_1 _28796_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1693),
    .D(_01164_),
    .Q_N(_12885_),
    .Q(\atari2600.tia.hmbl[0] ));
 sg13g2_dfrbp_1 _28797_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1692),
    .D(_01165_),
    .Q_N(_12884_),
    .Q(\atari2600.tia.hmbl[1] ));
 sg13g2_dfrbp_1 _28798_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1691),
    .D(_01166_),
    .Q_N(_12883_),
    .Q(\atari2600.tia.hmbl[2] ));
 sg13g2_dfrbp_1 _28799_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net965),
    .D(_01167_),
    .Q_N(_13844_),
    .Q(\atari2600.tia.hmbl[3] ));
 sg13g2_dfrbp_1 _28800_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net966),
    .D(_00023_),
    .Q_N(_13845_),
    .Q(\atari2600.tia.cx[0] ));
 sg13g2_dfrbp_1 _28801_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net967),
    .D(_00029_),
    .Q_N(_13846_),
    .Q(\atari2600.tia.cx[1] ));
 sg13g2_dfrbp_1 _28802_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net968),
    .D(net2982),
    .Q_N(_13847_),
    .Q(\atari2600.tia.cx[2] ));
 sg13g2_dfrbp_1 _28803_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net969),
    .D(net3075),
    .Q_N(_13848_),
    .Q(\atari2600.tia.cx[3] ));
 sg13g2_dfrbp_1 _28804_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net970),
    .D(_00032_),
    .Q_N(_13849_),
    .Q(\atari2600.tia.cx[4] ));
 sg13g2_dfrbp_1 _28805_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net971),
    .D(_00033_),
    .Q_N(_13850_),
    .Q(\atari2600.tia.cx[5] ));
 sg13g2_dfrbp_1 _28806_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net972),
    .D(_00034_),
    .Q_N(_13851_),
    .Q(\atari2600.tia.cx[6] ));
 sg13g2_dfrbp_1 _28807_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net973),
    .D(net2973),
    .Q_N(_13852_),
    .Q(\atari2600.tia.cx[7] ));
 sg13g2_dfrbp_1 _28808_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net974),
    .D(_00036_),
    .Q_N(_13853_),
    .Q(\atari2600.tia.cx[8] ));
 sg13g2_dfrbp_1 _28809_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net975),
    .D(net2993),
    .Q_N(_13854_),
    .Q(\atari2600.tia.cx[9] ));
 sg13g2_dfrbp_1 _28810_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net976),
    .D(_00024_),
    .Q_N(_13855_),
    .Q(\atari2600.tia.cx[10] ));
 sg13g2_dfrbp_1 _28811_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net977),
    .D(_00025_),
    .Q_N(_13856_),
    .Q(\atari2600.tia.cx[11] ));
 sg13g2_dfrbp_1 _28812_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net978),
    .D(_00026_),
    .Q_N(_13857_),
    .Q(\atari2600.tia.cx[12] ));
 sg13g2_dfrbp_1 _28813_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1151),
    .D(_00027_),
    .Q_N(_13858_),
    .Q(\atari2600.tia.cx[13] ));
 sg13g2_dfrbp_1 _28814_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1690),
    .D(_00028_),
    .Q_N(_12882_),
    .Q(\atari2600.tia.cx[14] ));
 sg13g2_dfrbp_1 _28815_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1689),
    .D(_01168_),
    .Q_N(_12881_),
    .Q(\atari2600.tia.cx_clr ));
 sg13g2_dfrbp_1 _28816_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1688),
    .D(_01169_),
    .Q_N(_12880_),
    .Q(\atari2600.tia.audc0[0] ));
 sg13g2_dfrbp_1 _28817_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1687),
    .D(_01170_),
    .Q_N(_12879_),
    .Q(\atari2600.tia.audc0[1] ));
 sg13g2_dfrbp_1 _28818_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1686),
    .D(_01171_),
    .Q_N(_12878_),
    .Q(\atari2600.tia.audc0[2] ));
 sg13g2_dfrbp_1 _28819_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1685),
    .D(_01172_),
    .Q_N(_12877_),
    .Q(\atari2600.tia.audc0[3] ));
 sg13g2_dfrbp_1 _28820_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1684),
    .D(_01173_),
    .Q_N(_12876_),
    .Q(\atari2600.tia.audc1[0] ));
 sg13g2_dfrbp_1 _28821_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1683),
    .D(_01174_),
    .Q_N(_12875_),
    .Q(\atari2600.tia.audc1[1] ));
 sg13g2_dfrbp_1 _28822_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1682),
    .D(_01175_),
    .Q_N(_12874_),
    .Q(\atari2600.tia.audc1[2] ));
 sg13g2_dfrbp_1 _28823_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1681),
    .D(_01176_),
    .Q_N(_12873_),
    .Q(\atari2600.tia.audc1[3] ));
 sg13g2_dfrbp_1 _28824_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1680),
    .D(_01177_),
    .Q_N(_12872_),
    .Q(\atari2600.tia.audv0[0] ));
 sg13g2_dfrbp_1 _28825_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1679),
    .D(_01178_),
    .Q_N(_12871_),
    .Q(\atari2600.tia.audv0[1] ));
 sg13g2_dfrbp_1 _28826_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1678),
    .D(_01179_),
    .Q_N(_12870_),
    .Q(\atari2600.tia.audv0[2] ));
 sg13g2_dfrbp_1 _28827_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1677),
    .D(_01180_),
    .Q_N(_12869_),
    .Q(\atari2600.tia.audv0[3] ));
 sg13g2_dfrbp_1 _28828_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1675),
    .D(_01181_),
    .Q_N(_12868_),
    .Q(\atari2600.tia.audv1[0] ));
 sg13g2_dfrbp_1 _28829_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1673),
    .D(_01182_),
    .Q_N(_12867_),
    .Q(\atari2600.tia.audv1[1] ));
 sg13g2_dfrbp_1 _28830_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1671),
    .D(_01183_),
    .Q_N(_12866_),
    .Q(\atari2600.tia.audv1[2] ));
 sg13g2_dfrbp_1 _28831_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1669),
    .D(_01184_),
    .Q_N(_12865_),
    .Q(\atari2600.tia.audv1[3] ));
 sg13g2_dfrbp_1 _28832_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1667),
    .D(_01185_),
    .Q_N(_00096_),
    .Q(\atari2600.tia.audf0[0] ));
 sg13g2_dfrbp_1 _28833_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1665),
    .D(_01186_),
    .Q_N(_12864_),
    .Q(\atari2600.tia.audf0[1] ));
 sg13g2_dfrbp_1 _28834_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1663),
    .D(_01187_),
    .Q_N(_12863_),
    .Q(\atari2600.tia.audf0[2] ));
 sg13g2_dfrbp_1 _28835_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1662),
    .D(_01188_),
    .Q_N(_12862_),
    .Q(\atari2600.tia.audf0[3] ));
 sg13g2_dfrbp_1 _28836_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1661),
    .D(_01189_),
    .Q_N(_00101_),
    .Q(\atari2600.tia.audf0[4] ));
 sg13g2_dfrbp_1 _28837_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1660),
    .D(_01190_),
    .Q_N(_00127_),
    .Q(\atari2600.tia.audf1[0] ));
 sg13g2_dfrbp_1 _28838_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1659),
    .D(_01191_),
    .Q_N(_12861_),
    .Q(\atari2600.tia.audf1[1] ));
 sg13g2_dfrbp_1 _28839_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1658),
    .D(_01192_),
    .Q_N(_12860_),
    .Q(\atari2600.tia.audf1[2] ));
 sg13g2_dfrbp_1 _28840_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1657),
    .D(_01193_),
    .Q_N(_12859_),
    .Q(\atari2600.tia.audf1[3] ));
 sg13g2_dfrbp_1 _28841_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1656),
    .D(_01194_),
    .Q_N(_00128_),
    .Q(\atari2600.tia.audf1[4] ));
 sg13g2_dfrbp_1 _28842_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1655),
    .D(net7373),
    .Q_N(_12858_),
    .Q(\atari2600.tia.p4_l ));
 sg13g2_dfrbp_1 _28843_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1654),
    .D(net6874),
    .Q_N(_12857_),
    .Q(\atari2600.tia.poly4_l.x[1] ));
 sg13g2_dfrbp_1 _28844_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1653),
    .D(_01197_),
    .Q_N(_12856_),
    .Q(\atari2600.tia.poly4_l.x[2] ));
 sg13g2_dfrbp_1 _28845_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1652),
    .D(net7137),
    .Q_N(_12855_),
    .Q(\atari2600.tia.poly4_l.x[3] ));
 sg13g2_dfrbp_1 _28846_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1651),
    .D(net4457),
    .Q_N(_12854_),
    .Q(\atari2600.tia.p5_l ));
 sg13g2_dfrbp_1 _28847_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1650),
    .D(_01200_),
    .Q_N(_12853_),
    .Q(\atari2600.tia.poly5_l.x[1] ));
 sg13g2_dfrbp_1 _28848_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1649),
    .D(_01201_),
    .Q_N(_12852_),
    .Q(\atari2600.tia.poly5_l.x[2] ));
 sg13g2_dfrbp_1 _28849_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1648),
    .D(_01202_),
    .Q_N(_12851_),
    .Q(\atari2600.tia.poly5_l.x[3] ));
 sg13g2_dfrbp_1 _28850_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1647),
    .D(_01203_),
    .Q_N(_12850_),
    .Q(\atari2600.tia.poly5_l.x[4] ));
 sg13g2_dfrbp_1 _28851_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1646),
    .D(net7226),
    .Q_N(_12849_),
    .Q(\atari2600.tia.p9_l ));
 sg13g2_dfrbp_1 _28852_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1645),
    .D(_01205_),
    .Q_N(_12848_),
    .Q(\atari2600.tia.poly9_l.x[1] ));
 sg13g2_dfrbp_1 _28853_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1644),
    .D(net7154),
    .Q_N(_12847_),
    .Q(\atari2600.tia.poly9_l.x[2] ));
 sg13g2_dfrbp_1 _28854_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1643),
    .D(_01207_),
    .Q_N(_12846_),
    .Q(\atari2600.tia.poly9_l.x[3] ));
 sg13g2_dfrbp_1 _28855_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1642),
    .D(net7163),
    .Q_N(_12845_),
    .Q(\atari2600.tia.poly9_l.x[4] ));
 sg13g2_dfrbp_1 _28856_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1641),
    .D(net6946),
    .Q_N(_12844_),
    .Q(\atari2600.tia.poly9_l.x[5] ));
 sg13g2_dfrbp_1 _28857_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1640),
    .D(_01210_),
    .Q_N(_12843_),
    .Q(\atari2600.tia.poly9_l.x[6] ));
 sg13g2_dfrbp_1 _28858_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1639),
    .D(net4512),
    .Q_N(_12842_),
    .Q(\atari2600.tia.poly9_l.x[7] ));
 sg13g2_dfrbp_1 _28859_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1638),
    .D(_01212_),
    .Q_N(_12841_),
    .Q(\atari2600.tia.poly9_l.x[8] ));
 sg13g2_dfrbp_1 _28860_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1637),
    .D(net7326),
    .Q_N(_12840_),
    .Q(\atari2600.tia.p4_r ));
 sg13g2_dfrbp_1 _28861_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1636),
    .D(net7245),
    .Q_N(_12839_),
    .Q(\atari2600.tia.poly4_r.x[1] ));
 sg13g2_dfrbp_1 _28862_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1635),
    .D(_01215_),
    .Q_N(_12838_),
    .Q(\atari2600.tia.poly4_r.x[2] ));
 sg13g2_dfrbp_1 _28863_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1634),
    .D(net4436),
    .Q_N(_12837_),
    .Q(\atari2600.tia.poly4_r.x[3] ));
 sg13g2_dfrbp_1 _28864_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1633),
    .D(net6816),
    .Q_N(_12836_),
    .Q(\atari2600.tia.p5_r ));
 sg13g2_dfrbp_1 _28865_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1632),
    .D(net7202),
    .Q_N(_12835_),
    .Q(\atari2600.tia.poly5_r.x[1] ));
 sg13g2_dfrbp_1 _28866_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1631),
    .D(net4867),
    .Q_N(_12834_),
    .Q(\atari2600.tia.poly5_r.x[2] ));
 sg13g2_dfrbp_1 _28867_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1630),
    .D(_01220_),
    .Q_N(_12833_),
    .Q(\atari2600.tia.poly5_r.x[3] ));
 sg13g2_dfrbp_1 _28868_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1629),
    .D(net6985),
    .Q_N(_12832_),
    .Q(\atari2600.tia.poly5_r.x[4] ));
 sg13g2_dfrbp_1 _28869_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1628),
    .D(net7258),
    .Q_N(_12831_),
    .Q(\atari2600.tia.p9_r ));
 sg13g2_dfrbp_1 _28870_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1627),
    .D(_01223_),
    .Q_N(_12830_),
    .Q(\atari2600.tia.poly9_r.x[1] ));
 sg13g2_dfrbp_1 _28871_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1626),
    .D(_01224_),
    .Q_N(_12829_),
    .Q(\atari2600.tia.poly9_r.x[2] ));
 sg13g2_dfrbp_1 _28872_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1625),
    .D(net4442),
    .Q_N(_12828_),
    .Q(\atari2600.tia.poly9_r.x[3] ));
 sg13g2_dfrbp_1 _28873_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1624),
    .D(net7206),
    .Q_N(_12827_),
    .Q(\atari2600.tia.poly9_r.x[4] ));
 sg13g2_dfrbp_1 _28874_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1623),
    .D(_01227_),
    .Q_N(_12826_),
    .Q(\atari2600.tia.poly9_r.x[5] ));
 sg13g2_dfrbp_1 _28875_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1622),
    .D(_01228_),
    .Q_N(_12825_),
    .Q(\atari2600.tia.poly9_r.x[6] ));
 sg13g2_dfrbp_1 _28876_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1621),
    .D(_01229_),
    .Q_N(_12824_),
    .Q(\atari2600.tia.poly9_r.x[7] ));
 sg13g2_dfrbp_1 _28877_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1620),
    .D(net4411),
    .Q_N(_12823_),
    .Q(\atari2600.tia.poly9_r.x[8] ));
 sg13g2_dfrbp_1 _28878_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1619),
    .D(_01231_),
    .Q_N(_12822_),
    .Q(\atari2600.ram[72][0] ));
 sg13g2_dfrbp_1 _28879_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1618),
    .D(_01232_),
    .Q_N(_12821_),
    .Q(\atari2600.ram[72][1] ));
 sg13g2_dfrbp_1 _28880_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1617),
    .D(_01233_),
    .Q_N(_12820_),
    .Q(\atari2600.ram[72][2] ));
 sg13g2_dfrbp_1 _28881_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1616),
    .D(_01234_),
    .Q_N(_12819_),
    .Q(\atari2600.ram[72][3] ));
 sg13g2_dfrbp_1 _28882_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1615),
    .D(_01235_),
    .Q_N(_12818_),
    .Q(\atari2600.ram[72][4] ));
 sg13g2_dfrbp_1 _28883_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1614),
    .D(_01236_),
    .Q_N(_12817_),
    .Q(\atari2600.ram[72][5] ));
 sg13g2_dfrbp_1 _28884_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1613),
    .D(_01237_),
    .Q_N(_12816_),
    .Q(\atari2600.ram[72][6] ));
 sg13g2_dfrbp_1 _28885_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1612),
    .D(_01238_),
    .Q_N(_12815_),
    .Q(\atari2600.ram[72][7] ));
 sg13g2_dfrbp_1 _28886_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1611),
    .D(net7029),
    .Q_N(_12814_),
    .Q(\atari2600.pia.interval[0] ));
 sg13g2_dfrbp_1 _28887_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1610),
    .D(net3122),
    .Q_N(_12813_),
    .Q(\atari2600.pia.instat[0] ));
 sg13g2_dfrbp_1 _28888_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1609),
    .D(_01241_),
    .Q_N(_12812_),
    .Q(\atari2600.ram[52][0] ));
 sg13g2_dfrbp_1 _28889_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1608),
    .D(_01242_),
    .Q_N(_12811_),
    .Q(\atari2600.ram[52][1] ));
 sg13g2_dfrbp_1 _28890_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1607),
    .D(_01243_),
    .Q_N(_12810_),
    .Q(\atari2600.ram[52][2] ));
 sg13g2_dfrbp_1 _28891_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1606),
    .D(_01244_),
    .Q_N(_12809_),
    .Q(\atari2600.ram[52][3] ));
 sg13g2_dfrbp_1 _28892_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1605),
    .D(_01245_),
    .Q_N(_12808_),
    .Q(\atari2600.ram[52][4] ));
 sg13g2_dfrbp_1 _28893_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1604),
    .D(_01246_),
    .Q_N(_12807_),
    .Q(\atari2600.ram[52][5] ));
 sg13g2_dfrbp_1 _28894_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1603),
    .D(_01247_),
    .Q_N(_12806_),
    .Q(\atari2600.ram[52][6] ));
 sg13g2_dfrbp_1 _28895_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1602),
    .D(_01248_),
    .Q_N(_12805_),
    .Q(\atari2600.ram[52][7] ));
 sg13g2_dfrbp_1 _28896_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1601),
    .D(_01249_),
    .Q_N(_12804_),
    .Q(\atari2600.ram[51][0] ));
 sg13g2_dfrbp_1 _28897_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1600),
    .D(_01250_),
    .Q_N(_12803_),
    .Q(\atari2600.ram[51][1] ));
 sg13g2_dfrbp_1 _28898_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1599),
    .D(_01251_),
    .Q_N(_12802_),
    .Q(\atari2600.ram[51][2] ));
 sg13g2_dfrbp_1 _28899_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1598),
    .D(_01252_),
    .Q_N(_12801_),
    .Q(\atari2600.ram[51][3] ));
 sg13g2_dfrbp_1 _28900_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1597),
    .D(_01253_),
    .Q_N(_12800_),
    .Q(\atari2600.ram[51][4] ));
 sg13g2_dfrbp_1 _28901_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1596),
    .D(_01254_),
    .Q_N(_12799_),
    .Q(\atari2600.ram[51][5] ));
 sg13g2_dfrbp_1 _28902_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1595),
    .D(_01255_),
    .Q_N(_12798_),
    .Q(\atari2600.ram[51][6] ));
 sg13g2_dfrbp_1 _28903_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1594),
    .D(_01256_),
    .Q_N(_12797_),
    .Q(\atari2600.ram[51][7] ));
 sg13g2_dfrbp_1 _28904_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1593),
    .D(_01257_),
    .Q_N(_12796_),
    .Q(\atari2600.ram[50][0] ));
 sg13g2_dfrbp_1 _28905_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1592),
    .D(_01258_),
    .Q_N(_12795_),
    .Q(\atari2600.ram[50][1] ));
 sg13g2_dfrbp_1 _28906_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1591),
    .D(_01259_),
    .Q_N(_12794_),
    .Q(\atari2600.ram[50][2] ));
 sg13g2_dfrbp_1 _28907_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1582),
    .D(_01260_),
    .Q_N(_12793_),
    .Q(\atari2600.ram[50][3] ));
 sg13g2_dfrbp_1 _28908_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1581),
    .D(_01261_),
    .Q_N(_12792_),
    .Q(\atari2600.ram[50][4] ));
 sg13g2_dfrbp_1 _28909_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1580),
    .D(_01262_),
    .Q_N(_12791_),
    .Q(\atari2600.ram[50][5] ));
 sg13g2_dfrbp_1 _28910_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1579),
    .D(_01263_),
    .Q_N(_12790_),
    .Q(\atari2600.ram[50][6] ));
 sg13g2_dfrbp_1 _28911_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1578),
    .D(_01264_),
    .Q_N(_12789_),
    .Q(\atari2600.ram[50][7] ));
 sg13g2_dfrbp_1 _28912_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1577),
    .D(_01265_),
    .Q_N(_12788_),
    .Q(\atari2600.ram[4][0] ));
 sg13g2_dfrbp_1 _28913_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1576),
    .D(_01266_),
    .Q_N(_12787_),
    .Q(\atari2600.ram[4][1] ));
 sg13g2_dfrbp_1 _28914_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1575),
    .D(_01267_),
    .Q_N(_12786_),
    .Q(\atari2600.ram[4][2] ));
 sg13g2_dfrbp_1 _28915_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1574),
    .D(_01268_),
    .Q_N(_12785_),
    .Q(\atari2600.ram[4][3] ));
 sg13g2_dfrbp_1 _28916_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1573),
    .D(_01269_),
    .Q_N(_12784_),
    .Q(\atari2600.ram[4][4] ));
 sg13g2_dfrbp_1 _28917_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1572),
    .D(_01270_),
    .Q_N(_12783_),
    .Q(\atari2600.ram[4][5] ));
 sg13g2_dfrbp_1 _28918_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1571),
    .D(_01271_),
    .Q_N(_12782_),
    .Q(\atari2600.ram[4][6] ));
 sg13g2_dfrbp_1 _28919_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1570),
    .D(_01272_),
    .Q_N(_12781_),
    .Q(\atari2600.ram[4][7] ));
 sg13g2_dfrbp_1 _28920_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1569),
    .D(_01273_),
    .Q_N(_12780_),
    .Q(\atari2600.ram[48][0] ));
 sg13g2_dfrbp_1 _28921_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1568),
    .D(_01274_),
    .Q_N(_12779_),
    .Q(\atari2600.ram[48][1] ));
 sg13g2_dfrbp_1 _28922_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1567),
    .D(_01275_),
    .Q_N(_12778_),
    .Q(\atari2600.ram[48][2] ));
 sg13g2_dfrbp_1 _28923_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net1566),
    .D(_01276_),
    .Q_N(_12777_),
    .Q(\atari2600.ram[48][3] ));
 sg13g2_dfrbp_1 _28924_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1565),
    .D(_01277_),
    .Q_N(_12776_),
    .Q(\atari2600.ram[48][4] ));
 sg13g2_dfrbp_1 _28925_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net1564),
    .D(_01278_),
    .Q_N(_12775_),
    .Q(\atari2600.ram[48][5] ));
 sg13g2_dfrbp_1 _28926_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net1563),
    .D(_01279_),
    .Q_N(_12774_),
    .Q(\atari2600.ram[48][6] ));
 sg13g2_dfrbp_1 _28927_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1562),
    .D(_01280_),
    .Q_N(_12773_),
    .Q(\atari2600.ram[48][7] ));
 sg13g2_dfrbp_1 _28928_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net1561),
    .D(_01281_),
    .Q_N(_12772_),
    .Q(\atari2600.ram[37][0] ));
 sg13g2_dfrbp_1 _28929_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net1560),
    .D(_01282_),
    .Q_N(_12771_),
    .Q(\atari2600.ram[37][1] ));
 sg13g2_dfrbp_1 _28930_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1559),
    .D(_01283_),
    .Q_N(_12770_),
    .Q(\atari2600.ram[37][2] ));
 sg13g2_dfrbp_1 _28931_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1558),
    .D(_01284_),
    .Q_N(_12769_),
    .Q(\atari2600.ram[37][3] ));
 sg13g2_dfrbp_1 _28932_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net1557),
    .D(_01285_),
    .Q_N(_12768_),
    .Q(\atari2600.ram[37][4] ));
 sg13g2_dfrbp_1 _28933_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1556),
    .D(_01286_),
    .Q_N(_12767_),
    .Q(\atari2600.ram[37][5] ));
 sg13g2_dfrbp_1 _28934_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net1555),
    .D(_01287_),
    .Q_N(_12766_),
    .Q(\atari2600.ram[37][6] ));
 sg13g2_dfrbp_1 _28935_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1554),
    .D(_01288_),
    .Q_N(_12765_),
    .Q(\atari2600.ram[37][7] ));
 sg13g2_dfrbp_1 _28936_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1553),
    .D(_01289_),
    .Q_N(_12764_),
    .Q(\atari2600.ram[47][0] ));
 sg13g2_dfrbp_1 _28937_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1552),
    .D(_01290_),
    .Q_N(_12763_),
    .Q(\atari2600.ram[47][1] ));
 sg13g2_dfrbp_1 _28938_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1551),
    .D(_01291_),
    .Q_N(_12762_),
    .Q(\atari2600.ram[47][2] ));
 sg13g2_dfrbp_1 _28939_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1550),
    .D(_01292_),
    .Q_N(_12761_),
    .Q(\atari2600.ram[47][3] ));
 sg13g2_dfrbp_1 _28940_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1549),
    .D(_01293_),
    .Q_N(_12760_),
    .Q(\atari2600.ram[47][4] ));
 sg13g2_dfrbp_1 _28941_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1548),
    .D(_01294_),
    .Q_N(_12759_),
    .Q(\atari2600.ram[47][5] ));
 sg13g2_dfrbp_1 _28942_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1547),
    .D(_01295_),
    .Q_N(_12758_),
    .Q(\atari2600.ram[47][6] ));
 sg13g2_dfrbp_1 _28943_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1546),
    .D(_01296_),
    .Q_N(_12757_),
    .Q(\atari2600.ram[47][7] ));
 sg13g2_dfrbp_1 _28944_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1545),
    .D(_01297_),
    .Q_N(_12756_),
    .Q(\atari2600.ram[32][0] ));
 sg13g2_dfrbp_1 _28945_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1544),
    .D(_01298_),
    .Q_N(_12755_),
    .Q(\atari2600.ram[32][1] ));
 sg13g2_dfrbp_1 _28946_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1543),
    .D(_01299_),
    .Q_N(_12754_),
    .Q(\atari2600.ram[32][2] ));
 sg13g2_dfrbp_1 _28947_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1542),
    .D(_01300_),
    .Q_N(_12753_),
    .Q(\atari2600.ram[32][3] ));
 sg13g2_dfrbp_1 _28948_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1541),
    .D(_01301_),
    .Q_N(_12752_),
    .Q(\atari2600.ram[32][4] ));
 sg13g2_dfrbp_1 _28949_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1540),
    .D(_01302_),
    .Q_N(_12751_),
    .Q(\atari2600.ram[32][5] ));
 sg13g2_dfrbp_1 _28950_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1539),
    .D(_01303_),
    .Q_N(_12750_),
    .Q(\atari2600.ram[32][6] ));
 sg13g2_dfrbp_1 _28951_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1538),
    .D(_01304_),
    .Q_N(_12749_),
    .Q(\atari2600.ram[32][7] ));
 sg13g2_dfrbp_1 _28952_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1537),
    .D(_01305_),
    .Q_N(_12748_),
    .Q(\atari2600.cpu.AXYS[0][0] ));
 sg13g2_dfrbp_1 _28953_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1536),
    .D(_01306_),
    .Q_N(_12747_),
    .Q(\atari2600.cpu.AXYS[0][1] ));
 sg13g2_dfrbp_1 _28954_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1535),
    .D(_01307_),
    .Q_N(_12746_),
    .Q(\atari2600.cpu.AXYS[0][2] ));
 sg13g2_dfrbp_1 _28955_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1534),
    .D(_01308_),
    .Q_N(_12745_),
    .Q(\atari2600.cpu.AXYS[0][3] ));
 sg13g2_dfrbp_1 _28956_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1533),
    .D(net4499),
    .Q_N(_12744_),
    .Q(\atari2600.cpu.AXYS[0][4] ));
 sg13g2_dfrbp_1 _28957_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1532),
    .D(_01310_),
    .Q_N(_12743_),
    .Q(\atari2600.cpu.AXYS[0][5] ));
 sg13g2_dfrbp_1 _28958_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1531),
    .D(_01311_),
    .Q_N(_12742_),
    .Q(\atari2600.cpu.AXYS[0][6] ));
 sg13g2_dfrbp_1 _28959_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1530),
    .D(_01312_),
    .Q_N(_12741_),
    .Q(\atari2600.cpu.AXYS[0][7] ));
 sg13g2_dfrbp_1 _28960_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1529),
    .D(_01313_),
    .Q_N(_12740_),
    .Q(\atari2600.tia.diag[76] ));
 sg13g2_dfrbp_1 _28961_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1528),
    .D(_01314_),
    .Q_N(_12739_),
    .Q(\atari2600.tia.diag[77] ));
 sg13g2_dfrbp_1 _28962_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1527),
    .D(_01315_),
    .Q_N(_12738_),
    .Q(\atari2600.tia.diag[78] ));
 sg13g2_dfrbp_1 _28963_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1526),
    .D(_01316_),
    .Q_N(_12737_),
    .Q(\atari2600.tia.diag[79] ));
 sg13g2_dfrbp_1 _28964_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1525),
    .D(_01317_),
    .Q_N(_12736_),
    .Q(\atari2600.tia.diag[80] ));
 sg13g2_dfrbp_1 _28965_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1524),
    .D(_01318_),
    .Q_N(_12735_),
    .Q(\atari2600.tia.diag[81] ));
 sg13g2_dfrbp_1 _28966_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1523),
    .D(_01319_),
    .Q_N(_12734_),
    .Q(\atari2600.tia.diag[82] ));
 sg13g2_dfrbp_1 _28967_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1522),
    .D(_01320_),
    .Q_N(_12733_),
    .Q(\atari2600.tia.diag[83] ));
 sg13g2_dfrbp_1 _28968_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1521),
    .D(_01321_),
    .Q_N(_12732_),
    .Q(\atari2600.tia.diag[84] ));
 sg13g2_dfrbp_1 _28969_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1520),
    .D(_01322_),
    .Q_N(_12731_),
    .Q(\atari2600.tia.diag[85] ));
 sg13g2_dfrbp_1 _28970_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1519),
    .D(_01323_),
    .Q_N(_12730_),
    .Q(\atari2600.tia.diag[86] ));
 sg13g2_dfrbp_1 _28971_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1518),
    .D(_01324_),
    .Q_N(_12729_),
    .Q(\atari2600.tia.diag[87] ));
 sg13g2_dfrbp_1 _28972_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1517),
    .D(_01325_),
    .Q_N(_12728_),
    .Q(\atari2600.ram[46][0] ));
 sg13g2_dfrbp_1 _28973_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1516),
    .D(_01326_),
    .Q_N(_12727_),
    .Q(\atari2600.ram[46][1] ));
 sg13g2_dfrbp_1 _28974_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1515),
    .D(_01327_),
    .Q_N(_12726_),
    .Q(\atari2600.ram[46][2] ));
 sg13g2_dfrbp_1 _28975_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1514),
    .D(_01328_),
    .Q_N(_12725_),
    .Q(\atari2600.ram[46][3] ));
 sg13g2_dfrbp_1 _28976_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1513),
    .D(_01329_),
    .Q_N(_12724_),
    .Q(\atari2600.ram[46][4] ));
 sg13g2_dfrbp_1 _28977_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1512),
    .D(_01330_),
    .Q_N(_12723_),
    .Q(\atari2600.ram[46][5] ));
 sg13g2_dfrbp_1 _28978_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1511),
    .D(_01331_),
    .Q_N(_12722_),
    .Q(\atari2600.ram[46][6] ));
 sg13g2_dfrbp_1 _28979_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1510),
    .D(_01332_),
    .Q_N(_12721_),
    .Q(\atari2600.ram[46][7] ));
 sg13g2_dfrbp_1 _28980_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1509),
    .D(_01333_),
    .Q_N(_12720_),
    .Q(\atari2600.ram[25][0] ));
 sg13g2_dfrbp_1 _28981_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1508),
    .D(_01334_),
    .Q_N(_12719_),
    .Q(\atari2600.ram[25][1] ));
 sg13g2_dfrbp_1 _28982_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1507),
    .D(_01335_),
    .Q_N(_12718_),
    .Q(\atari2600.ram[25][2] ));
 sg13g2_dfrbp_1 _28983_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1506),
    .D(_01336_),
    .Q_N(_12717_),
    .Q(\atari2600.ram[25][3] ));
 sg13g2_dfrbp_1 _28984_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1505),
    .D(_01337_),
    .Q_N(_12716_),
    .Q(\atari2600.ram[25][4] ));
 sg13g2_dfrbp_1 _28985_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1504),
    .D(_01338_),
    .Q_N(_12715_),
    .Q(\atari2600.ram[25][5] ));
 sg13g2_dfrbp_1 _28986_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1503),
    .D(_01339_),
    .Q_N(_12714_),
    .Q(\atari2600.ram[25][6] ));
 sg13g2_dfrbp_1 _28987_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1152),
    .D(_01340_),
    .Q_N(_13859_),
    .Q(\atari2600.ram[25][7] ));
 sg13g2_dfrbp_1 _28988_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1153),
    .D(_00019_),
    .Q_N(_13860_),
    .Q(\atari2600.tia.p1_copies[1] ));
 sg13g2_dfrbp_1 _28989_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1154),
    .D(_00020_),
    .Q_N(_13861_),
    .Q(\atari2600.tia.p1_copies[2] ));
 sg13g2_dfrbp_1 _28990_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1188),
    .D(_00017_),
    .Q_N(_13862_),
    .Q(\atari2600.tia.p0_copies[1] ));
 sg13g2_dfrbp_1 _28991_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1502),
    .D(_00018_),
    .Q_N(_12713_),
    .Q(\atari2600.tia.p0_copies[2] ));
 sg13g2_dfrbp_1 _28992_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1501),
    .D(_01341_),
    .Q_N(_00082_),
    .Q(\atari2600.cpu.DI[0] ));
 sg13g2_dfrbp_1 _28993_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1500),
    .D(_01342_),
    .Q_N(_00080_),
    .Q(\atari2600.cpu.DI[1] ));
 sg13g2_dfrbp_1 _28994_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1499),
    .D(_01343_),
    .Q_N(_12712_),
    .Q(\atari2600.cpu.DI[2] ));
 sg13g2_dfrbp_1 _28995_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1498),
    .D(_01344_),
    .Q_N(_12711_),
    .Q(\atari2600.cpu.DI[3] ));
 sg13g2_dfrbp_1 _28996_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1497),
    .D(_01345_),
    .Q_N(_12710_),
    .Q(\atari2600.cpu.DI[4] ));
 sg13g2_dfrbp_1 _28997_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1496),
    .D(_01346_),
    .Q_N(_12709_),
    .Q(\atari2600.cpu.DI[5] ));
 sg13g2_dfrbp_1 _28998_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1495),
    .D(_01347_),
    .Q_N(_12708_),
    .Q(\atari2600.cpu.DI[6] ));
 sg13g2_dfrbp_1 _28999_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1494),
    .D(net7474),
    .Q_N(_12707_),
    .Q(\atari2600.cpu.DI[7] ));
 sg13g2_dfrbp_1 _29000_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1493),
    .D(_01349_),
    .Q_N(_12706_),
    .Q(\atari2600.cpu.cond_code[0] ));
 sg13g2_dfrbp_1 _29001_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1492),
    .D(_01350_),
    .Q_N(_12705_),
    .Q(\atari2600.cpu.cond_code[1] ));
 sg13g2_dfrbp_1 _29002_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1491),
    .D(_01351_),
    .Q_N(_00056_),
    .Q(\atari2600.cpu.cond_code[2] ));
 sg13g2_dfrbp_1 _29003_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1490),
    .D(_01352_),
    .Q_N(_00134_),
    .Q(\atari2600.cpu.plp ));
 sg13g2_dfrbp_1 _29004_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1489),
    .D(_01353_),
    .Q_N(_12704_),
    .Q(\atari2600.cpu.php ));
 sg13g2_dfrbp_1 _29005_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1488),
    .D(_01354_),
    .Q_N(_00166_),
    .Q(\atari2600.cpu.clc ));
 sg13g2_dfrbp_1 _29006_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1487),
    .D(_01355_),
    .Q_N(_12703_),
    .Q(\atari2600.cpu.sec ));
 sg13g2_dfrbp_1 _29007_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1486),
    .D(_01356_),
    .Q_N(_00164_),
    .Q(\atari2600.cpu.cld ));
 sg13g2_dfrbp_1 _29008_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1485),
    .D(_01357_),
    .Q_N(_12702_),
    .Q(\atari2600.cpu.sed ));
 sg13g2_dfrbp_1 _29009_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1484),
    .D(net3008),
    .Q_N(_00165_),
    .Q(\atari2600.cpu.cli ));
 sg13g2_dfrbp_1 _29010_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1483),
    .D(net3547),
    .Q_N(_12701_),
    .Q(\atari2600.cpu.sei ));
 sg13g2_dfrbp_1 _29011_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1482),
    .D(_01360_),
    .Q_N(_12700_),
    .Q(\atari2600.cpu.clv ));
 sg13g2_dfrbp_1 _29012_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1481),
    .D(_01361_),
    .Q_N(_12699_),
    .Q(\atari2600.cpu.bit_ins ));
 sg13g2_dfrbp_1 _29013_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1480),
    .D(_01362_),
    .Q_N(_12698_),
    .Q(\atari2600.cpu.rotate ));
 sg13g2_dfrbp_1 _29014_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1479),
    .D(_01363_),
    .Q_N(_12697_),
    .Q(\atari2600.cpu.shift_right ));
 sg13g2_dfrbp_1 _29015_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1478),
    .D(_01364_),
    .Q_N(_12696_),
    .Q(\atari2600.cpu.compare ));
 sg13g2_dfrbp_1 _29016_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1477),
    .D(_01365_),
    .Q_N(_12695_),
    .Q(\atari2600.cpu.adc_bcd ));
 sg13g2_dfrbp_1 _29017_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1476),
    .D(_01366_),
    .Q_N(_12694_),
    .Q(\atari2600.cpu.shift ));
 sg13g2_dfrbp_1 _29018_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1475),
    .D(_01367_),
    .Q_N(_12693_),
    .Q(\atari2600.cpu.adc_sbc ));
 sg13g2_dfrbp_1 _29019_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1474),
    .D(_01368_),
    .Q_N(_12692_),
    .Q(\atari2600.cpu.inc ));
 sg13g2_dfrbp_1 _29020_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1473),
    .D(_01369_),
    .Q_N(_12691_),
    .Q(\atari2600.cpu.load_only ));
 sg13g2_dfrbp_1 _29021_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1472),
    .D(_01370_),
    .Q_N(_00133_),
    .Q(\atari2600.cpu.write_back ));
 sg13g2_dfrbp_1 _29022_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1471),
    .D(net7465),
    .Q_N(_12690_),
    .Q(\atari2600.cpu.store ));
 sg13g2_dfrbp_1 _29023_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1470),
    .D(_01372_),
    .Q_N(_12689_),
    .Q(\atari2600.cpu.index_y ));
 sg13g2_dfrbp_1 _29024_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1189),
    .D(_01373_),
    .Q_N(_13863_),
    .Q(\atari2600.cpu.res ));
 sg13g2_dfrbp_1 _29025_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1190),
    .D(\atari2600.cpu.DIMUX[0] ),
    .Q_N(_00081_),
    .Q(\atari2600.cpu.DIHOLD[0] ));
 sg13g2_dfrbp_1 _29026_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1191),
    .D(\atari2600.cpu.DIMUX[1] ),
    .Q_N(_00079_),
    .Q(\atari2600.cpu.DIHOLD[1] ));
 sg13g2_dfrbp_1 _29027_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1192),
    .D(net7312),
    .Q_N(_13864_),
    .Q(\atari2600.cpu.DIHOLD[2] ));
 sg13g2_dfrbp_1 _29028_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(net7268),
    .Q_N(_13865_),
    .Q(\atari2600.cpu.DIHOLD[3] ));
 sg13g2_dfrbp_1 _29029_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1194),
    .D(\atari2600.cpu.DIMUX[4] ),
    .Q_N(_13866_),
    .Q(\atari2600.cpu.DIHOLD[4] ));
 sg13g2_dfrbp_1 _29030_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1195),
    .D(\atari2600.cpu.DIMUX[5] ),
    .Q_N(_13867_),
    .Q(\atari2600.cpu.DIHOLD[5] ));
 sg13g2_dfrbp_1 _29031_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1212),
    .D(net7300),
    .Q_N(_13868_),
    .Q(\atari2600.cpu.DIHOLD[6] ));
 sg13g2_dfrbp_1 _29032_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1469),
    .D(\atari2600.cpu.DIMUX[7] ),
    .Q_N(_12688_),
    .Q(\atari2600.cpu.DIHOLD[7] ));
 sg13g2_dfrbp_1 _29033_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1468),
    .D(_01374_),
    .Q_N(_12687_),
    .Q(\atari2600.cpu.load_reg ));
 sg13g2_dfrbp_1 _29034_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1467),
    .D(_01375_),
    .Q_N(_12686_),
    .Q(\atari2600.cpu.IRHOLD_valid ));
 sg13g2_dfrbp_1 _29035_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1466),
    .D(net4641),
    .Q_N(_12685_),
    .Q(\atari2600.cpu.IRHOLD[0] ));
 sg13g2_dfrbp_1 _29036_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1465),
    .D(_01377_),
    .Q_N(_12684_),
    .Q(\atari2600.cpu.IRHOLD[1] ));
 sg13g2_dfrbp_1 _29037_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1464),
    .D(net7182),
    .Q_N(_12683_),
    .Q(\atari2600.cpu.IRHOLD[2] ));
 sg13g2_dfrbp_1 _29038_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1463),
    .D(net7188),
    .Q_N(_12682_),
    .Q(\atari2600.cpu.IRHOLD[3] ));
 sg13g2_dfrbp_1 _29039_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1462),
    .D(_01380_),
    .Q_N(_12681_),
    .Q(\atari2600.cpu.IRHOLD[4] ));
 sg13g2_dfrbp_1 _29040_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1461),
    .D(_01381_),
    .Q_N(_12680_),
    .Q(\atari2600.cpu.IRHOLD[5] ));
 sg13g2_dfrbp_1 _29041_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1460),
    .D(net7251),
    .Q_N(_12679_),
    .Q(\atari2600.cpu.IRHOLD[6] ));
 sg13g2_dfrbp_1 _29042_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1459),
    .D(_01383_),
    .Q_N(_12678_),
    .Q(\atari2600.cpu.IRHOLD[7] ));
 sg13g2_dfrbp_1 _29043_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1458),
    .D(net2947),
    .Q_N(_00136_),
    .Q(\atari2600.cpu.D ));
 sg13g2_dfrbp_1 _29044_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1457),
    .D(net7192),
    .Q_N(_00075_),
    .Q(\atari2600.cpu.I ));
 sg13g2_dfrbp_1 _29045_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1456),
    .D(net7219),
    .Q_N(_00137_),
    .Q(\atari2600.cpu.V ));
 sg13g2_dfrbp_1 _29046_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1455),
    .D(_01387_),
    .Q_N(_00138_),
    .Q(\atari2600.cpu.N ));
 sg13g2_dfrbp_1 _29047_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1454),
    .D(net7120),
    .Q_N(_00073_),
    .Q(\atari2600.cpu.Z ));
 sg13g2_dfrbp_1 _29048_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1287),
    .D(net7518),
    .Q_N(_00077_),
    .Q(\atari2600.cpu.C ));
 sg13g2_dfrbp_1 _29049_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1453),
    .D(net4938),
    .Q_N(_00163_),
    .Q(\atari2600.cpu.adj_bcd ));
 sg13g2_dfrbp_1 _29050_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1452),
    .D(net7144),
    .Q_N(_12677_),
    .Q(\atari2600.cpu.backwards ));
 sg13g2_dfrbp_1 _29051_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1451),
    .D(net7097),
    .Q_N(_12676_),
    .Q(\atari2600.cpu.ABL[0] ));
 sg13g2_dfrbp_1 _29052_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1450),
    .D(net7249),
    .Q_N(_12675_),
    .Q(\atari2600.cpu.ABL[1] ));
 sg13g2_dfrbp_1 _29053_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1449),
    .D(net7004),
    .Q_N(_12674_),
    .Q(\atari2600.cpu.ABL[2] ));
 sg13g2_dfrbp_1 _29054_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1448),
    .D(net7060),
    .Q_N(_12673_),
    .Q(\atari2600.cpu.ABL[3] ));
 sg13g2_dfrbp_1 _29055_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1447),
    .D(net7151),
    .Q_N(_12672_),
    .Q(\atari2600.cpu.ABL[4] ));
 sg13g2_dfrbp_1 _29056_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1446),
    .D(_01396_),
    .Q_N(_12671_),
    .Q(\atari2600.cpu.ABL[5] ));
 sg13g2_dfrbp_1 _29057_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1445),
    .D(_01397_),
    .Q_N(_12670_),
    .Q(\atari2600.cpu.ABL[6] ));
 sg13g2_dfrbp_1 _29058_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1444),
    .D(_01398_),
    .Q_N(_12669_),
    .Q(\atari2600.cpu.ABL[7] ));
 sg13g2_dfrbp_1 _29059_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1443),
    .D(_01399_),
    .Q_N(_12668_),
    .Q(\atari2600.cpu.ALU.AI7 ));
 sg13g2_dfrbp_1 _29060_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1442),
    .D(_01400_),
    .Q_N(_12667_),
    .Q(\atari2600.cpu.ADD[0] ));
 sg13g2_dfrbp_1 _29061_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1441),
    .D(_01401_),
    .Q_N(_00074_),
    .Q(\atari2600.cpu.ADD[1] ));
 sg13g2_dfrbp_1 _29062_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1440),
    .D(_01402_),
    .Q_N(_00076_),
    .Q(\atari2600.cpu.ADD[2] ));
 sg13g2_dfrbp_1 _29063_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1439),
    .D(_01403_),
    .Q_N(_00090_),
    .Q(\atari2600.cpu.ADD[3] ));
 sg13g2_dfrbp_1 _29064_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1438),
    .D(_01404_),
    .Q_N(_12666_),
    .Q(\atari2600.cpu.ADD[4] ));
 sg13g2_dfrbp_1 _29065_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1437),
    .D(_01405_),
    .Q_N(_00086_),
    .Q(\atari2600.cpu.ADD[5] ));
 sg13g2_dfrbp_1 _29066_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1436),
    .D(_01406_),
    .Q_N(_00092_),
    .Q(\atari2600.cpu.ADD[6] ));
 sg13g2_dfrbp_1 _29067_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1435),
    .D(_01407_),
    .Q_N(_00091_),
    .Q(\atari2600.cpu.ADD[7] ));
 sg13g2_dfrbp_1 _29068_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1434),
    .D(_01408_),
    .Q_N(_12665_),
    .Q(\atari2600.cpu.ALU.HC ));
 sg13g2_dfrbp_1 _29069_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1433),
    .D(_01409_),
    .Q_N(_12664_),
    .Q(\atari2600.cpu.ALU.CO ));
 sg13g2_dfrbp_1 _29070_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1432),
    .D(_01410_),
    .Q_N(_00087_),
    .Q(\atari2600.cpu.PC[0] ));
 sg13g2_dfrbp_1 _29071_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1431),
    .D(net4444),
    .Q_N(_00088_),
    .Q(\atari2600.cpu.PC[1] ));
 sg13g2_dfrbp_1 _29072_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1430),
    .D(net3643),
    .Q_N(_00078_),
    .Q(\atari2600.cpu.PC[2] ));
 sg13g2_dfrbp_1 _29073_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1429),
    .D(_01413_),
    .Q_N(_00089_),
    .Q(\atari2600.cpu.PC[3] ));
 sg13g2_dfrbp_1 _29074_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1428),
    .D(net7009),
    .Q_N(_00085_),
    .Q(\atari2600.cpu.PC[4] ));
 sg13g2_dfrbp_1 _29075_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1427),
    .D(net7242),
    .Q_N(_00060_),
    .Q(\atari2600.cpu.PC[5] ));
 sg13g2_dfrbp_1 _29076_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1426),
    .D(net7146),
    .Q_N(_00061_),
    .Q(\atari2600.cpu.PC[6] ));
 sg13g2_dfrbp_1 _29077_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1425),
    .D(net7197),
    .Q_N(_00062_),
    .Q(\atari2600.cpu.PC[7] ));
 sg13g2_dfrbp_1 _29078_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1424),
    .D(net6865),
    .Q_N(_00063_),
    .Q(\atari2600.cpu.PC[8] ));
 sg13g2_dfrbp_1 _29079_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1423),
    .D(net7262),
    .Q_N(_00064_),
    .Q(\atari2600.cpu.PC[9] ));
 sg13g2_dfrbp_1 _29080_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1422),
    .D(net4481),
    .Q_N(_00065_),
    .Q(\atari2600.cpu.PC[10] ));
 sg13g2_dfrbp_1 _29081_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1421),
    .D(net7117),
    .Q_N(_00066_),
    .Q(\atari2600.cpu.PC[11] ));
 sg13g2_dfrbp_1 _29082_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1420),
    .D(net7176),
    .Q_N(_00067_),
    .Q(\atari2600.cpu.PC[12] ));
 sg13g2_dfrbp_1 _29083_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1419),
    .D(net7215),
    .Q_N(_00068_),
    .Q(\atari2600.cpu.PC[13] ));
 sg13g2_dfrbp_1 _29084_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1418),
    .D(_01424_),
    .Q_N(_12663_),
    .Q(\atari2600.cpu.PC[14] ));
 sg13g2_dfrbp_1 _29085_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1417),
    .D(_01425_),
    .Q_N(_12662_),
    .Q(\atari2600.cpu.PC[15] ));
 sg13g2_dfrbp_1 _29086_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1416),
    .D(_01426_),
    .Q_N(_12661_),
    .Q(\atari2600.ram[45][0] ));
 sg13g2_dfrbp_1 _29087_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1415),
    .D(_01427_),
    .Q_N(_12660_),
    .Q(\atari2600.ram[45][1] ));
 sg13g2_dfrbp_1 _29088_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1414),
    .D(_01428_),
    .Q_N(_12659_),
    .Q(\atari2600.ram[45][2] ));
 sg13g2_dfrbp_1 _29089_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1413),
    .D(_01429_),
    .Q_N(_12658_),
    .Q(\atari2600.ram[45][3] ));
 sg13g2_dfrbp_1 _29090_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1412),
    .D(_01430_),
    .Q_N(_12657_),
    .Q(\atari2600.ram[45][4] ));
 sg13g2_dfrbp_1 _29091_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1411),
    .D(_01431_),
    .Q_N(_12656_),
    .Q(\atari2600.ram[45][5] ));
 sg13g2_dfrbp_1 _29092_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1410),
    .D(_01432_),
    .Q_N(_12655_),
    .Q(\atari2600.ram[45][6] ));
 sg13g2_dfrbp_1 _29093_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1409),
    .D(_01433_),
    .Q_N(_12654_),
    .Q(\atari2600.ram[45][7] ));
 sg13g2_dfrbp_1 _29094_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1408),
    .D(_01434_),
    .Q_N(_12653_),
    .Q(\atari2600.ram[44][0] ));
 sg13g2_dfrbp_1 _29095_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1407),
    .D(_01435_),
    .Q_N(_12652_),
    .Q(\atari2600.ram[44][1] ));
 sg13g2_dfrbp_1 _29096_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1406),
    .D(_01436_),
    .Q_N(_12651_),
    .Q(\atari2600.ram[44][2] ));
 sg13g2_dfrbp_1 _29097_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1405),
    .D(_01437_),
    .Q_N(_12650_),
    .Q(\atari2600.ram[44][3] ));
 sg13g2_dfrbp_1 _29098_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1404),
    .D(_01438_),
    .Q_N(_12649_),
    .Q(\atari2600.ram[44][4] ));
 sg13g2_dfrbp_1 _29099_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1403),
    .D(_01439_),
    .Q_N(_12648_),
    .Q(\atari2600.ram[44][5] ));
 sg13g2_dfrbp_1 _29100_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1402),
    .D(_01440_),
    .Q_N(_12647_),
    .Q(\atari2600.ram[44][6] ));
 sg13g2_dfrbp_1 _29101_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1401),
    .D(_01441_),
    .Q_N(_12646_),
    .Q(\atari2600.ram[44][7] ));
 sg13g2_dfrbp_1 _29102_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1400),
    .D(_01442_),
    .Q_N(_12645_),
    .Q(\atari2600.clk_counter[0] ));
 sg13g2_dfrbp_1 _29103_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1399),
    .D(_01443_),
    .Q_N(_12644_),
    .Q(\atari2600.clk_counter[1] ));
 sg13g2_dfrbp_1 _29104_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1398),
    .D(_01444_),
    .Q_N(_12643_),
    .Q(\atari2600.clk_counter[2] ));
 sg13g2_dfrbp_1 _29105_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1396),
    .D(_01445_),
    .Q_N(_12642_),
    .Q(\atari2600.clk_counter[3] ));
 sg13g2_dfrbp_1 _29106_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1394),
    .D(_01446_),
    .Q_N(_12641_),
    .Q(\atari2600.clk_counter[4] ));
 sg13g2_dfrbp_1 _29107_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1392),
    .D(_01447_),
    .Q_N(_12640_),
    .Q(\atari2600.clk_counter[5] ));
 sg13g2_dfrbp_1 _29108_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1390),
    .D(_01448_),
    .Q_N(_12639_),
    .Q(\atari2600.clk_counter[6] ));
 sg13g2_dfrbp_1 _29109_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1388),
    .D(_01449_),
    .Q_N(_12638_),
    .Q(\atari2600.clk_counter[7] ));
 sg13g2_dfrbp_1 _29110_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1386),
    .D(net3067),
    .Q_N(_00129_),
    .Q(\atari2600.clk_counter[8] ));
 sg13g2_dfrbp_1 _29111_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1384),
    .D(_01451_),
    .Q_N(_12637_),
    .Q(\atari2600.ram[91][0] ));
 sg13g2_dfrbp_1 _29112_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1383),
    .D(_01452_),
    .Q_N(_12636_),
    .Q(\atari2600.ram[91][1] ));
 sg13g2_dfrbp_1 _29113_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1382),
    .D(_01453_),
    .Q_N(_12635_),
    .Q(\atari2600.ram[91][2] ));
 sg13g2_dfrbp_1 _29114_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1381),
    .D(_01454_),
    .Q_N(_12634_),
    .Q(\atari2600.ram[91][3] ));
 sg13g2_dfrbp_1 _29115_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1380),
    .D(_01455_),
    .Q_N(_12633_),
    .Q(\atari2600.ram[91][4] ));
 sg13g2_dfrbp_1 _29116_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1379),
    .D(_01456_),
    .Q_N(_12632_),
    .Q(\atari2600.ram[91][5] ));
 sg13g2_dfrbp_1 _29117_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1378),
    .D(_01457_),
    .Q_N(_12631_),
    .Q(\atari2600.ram[91][6] ));
 sg13g2_dfrbp_1 _29118_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1377),
    .D(_01458_),
    .Q_N(_12630_),
    .Q(\atari2600.ram[91][7] ));
 sg13g2_dfrbp_1 _29119_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1376),
    .D(_01459_),
    .Q_N(_12629_),
    .Q(\atari2600.ram[21][0] ));
 sg13g2_dfrbp_1 _29120_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1375),
    .D(_01460_),
    .Q_N(_12628_),
    .Q(\atari2600.ram[21][1] ));
 sg13g2_dfrbp_1 _29121_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1374),
    .D(_01461_),
    .Q_N(_12627_),
    .Q(\atari2600.ram[21][2] ));
 sg13g2_dfrbp_1 _29122_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1373),
    .D(_01462_),
    .Q_N(_12626_),
    .Q(\atari2600.ram[21][3] ));
 sg13g2_dfrbp_1 _29123_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1372),
    .D(_01463_),
    .Q_N(_12625_),
    .Q(\atari2600.ram[21][4] ));
 sg13g2_dfrbp_1 _29124_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1371),
    .D(_01464_),
    .Q_N(_12624_),
    .Q(\atari2600.ram[21][5] ));
 sg13g2_dfrbp_1 _29125_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1370),
    .D(_01465_),
    .Q_N(_12623_),
    .Q(\atari2600.ram[21][6] ));
 sg13g2_dfrbp_1 _29126_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1369),
    .D(_01466_),
    .Q_N(_12622_),
    .Q(\atari2600.ram[21][7] ));
 sg13g2_dfrbp_1 _29127_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1368),
    .D(_01467_),
    .Q_N(_12621_),
    .Q(\atari2600.ram[24][0] ));
 sg13g2_dfrbp_1 _29128_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1367),
    .D(_01468_),
    .Q_N(_12620_),
    .Q(\atari2600.ram[24][1] ));
 sg13g2_dfrbp_1 _29129_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1366),
    .D(_01469_),
    .Q_N(_12619_),
    .Q(\atari2600.ram[24][2] ));
 sg13g2_dfrbp_1 _29130_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1365),
    .D(_01470_),
    .Q_N(_12618_),
    .Q(\atari2600.ram[24][3] ));
 sg13g2_dfrbp_1 _29131_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1364),
    .D(_01471_),
    .Q_N(_12617_),
    .Q(\atari2600.ram[24][4] ));
 sg13g2_dfrbp_1 _29132_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1363),
    .D(_01472_),
    .Q_N(_12616_),
    .Q(\atari2600.ram[24][5] ));
 sg13g2_dfrbp_1 _29133_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1362),
    .D(_01473_),
    .Q_N(_12615_),
    .Q(\atari2600.ram[24][6] ));
 sg13g2_dfrbp_1 _29134_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1361),
    .D(_01474_),
    .Q_N(_12614_),
    .Q(\atari2600.ram[24][7] ));
 sg13g2_dfrbp_1 _29135_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1288),
    .D(_01475_),
    .Q_N(_13869_),
    .Q(\flash_rom.data_ready ));
 sg13g2_dfrbp_1 _29136_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1318),
    .D(net2929),
    .Q_N(_13870_),
    .Q(\gamepad_pmod.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _29137_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1360),
    .D(net2928),
    .Q_N(_12613_),
    .Q(\gamepad_pmod.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _29138_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1359),
    .D(net2956),
    .Q_N(_12612_),
    .Q(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _29139_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1358),
    .D(net6925),
    .Q_N(_12611_),
    .Q(\gamepad_pmod.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _29140_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1357),
    .D(net7095),
    .Q_N(_12610_),
    .Q(\gamepad_pmod.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _29141_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1356),
    .D(net7232),
    .Q_N(_12609_),
    .Q(\gamepad_pmod.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _29142_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1355),
    .D(net6710),
    .Q_N(_12608_),
    .Q(\gamepad_pmod.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _29143_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1354),
    .D(net6679),
    .Q_N(_12607_),
    .Q(\gamepad_pmod.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _29144_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1353),
    .D(_01482_),
    .Q_N(_12606_),
    .Q(\gamepad_pmod.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _29145_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1352),
    .D(_01483_),
    .Q_N(_12605_),
    .Q(\gamepad_pmod.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _29146_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1351),
    .D(net7084),
    .Q_N(_12604_),
    .Q(\gamepad_pmod.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _29147_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1350),
    .D(net7228),
    .Q_N(_12603_),
    .Q(\gamepad_pmod.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _29148_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1349),
    .D(net6810),
    .Q_N(_12602_),
    .Q(\gamepad_pmod.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _29149_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1348),
    .D(net4535),
    .Q_N(_12601_),
    .Q(\gamepad_pmod.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _29150_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1347),
    .D(_01488_),
    .Q_N(_12600_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _29151_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1346),
    .D(_01489_),
    .Q_N(_12599_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _29152_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1345),
    .D(_01490_),
    .Q_N(_12598_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _29153_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1344),
    .D(_01491_),
    .Q_N(_12597_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _29154_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1343),
    .D(_01492_),
    .Q_N(_12596_),
    .Q(\atari2600.ram[88][0] ));
 sg13g2_dfrbp_1 _29155_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1342),
    .D(_01493_),
    .Q_N(_12595_),
    .Q(\atari2600.ram[88][1] ));
 sg13g2_dfrbp_1 _29156_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1341),
    .D(_01494_),
    .Q_N(_12594_),
    .Q(\atari2600.ram[88][2] ));
 sg13g2_dfrbp_1 _29157_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1340),
    .D(_01495_),
    .Q_N(_12593_),
    .Q(\atari2600.ram[88][3] ));
 sg13g2_dfrbp_1 _29158_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1339),
    .D(_01496_),
    .Q_N(_12592_),
    .Q(\atari2600.ram[88][4] ));
 sg13g2_dfrbp_1 _29159_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1338),
    .D(_01497_),
    .Q_N(_12591_),
    .Q(\atari2600.ram[88][5] ));
 sg13g2_dfrbp_1 _29160_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1337),
    .D(_01498_),
    .Q_N(_12590_),
    .Q(\atari2600.ram[88][6] ));
 sg13g2_dfrbp_1 _29161_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1336),
    .D(_01499_),
    .Q_N(_12589_),
    .Q(\atari2600.ram[88][7] ));
 sg13g2_dfrbp_1 _29162_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1335),
    .D(_01500_),
    .Q_N(_12588_),
    .Q(\atari2600.ram[8][0] ));
 sg13g2_dfrbp_1 _29163_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1334),
    .D(_01501_),
    .Q_N(_12587_),
    .Q(\atari2600.ram[8][1] ));
 sg13g2_dfrbp_1 _29164_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1333),
    .D(_01502_),
    .Q_N(_12586_),
    .Q(\atari2600.ram[8][2] ));
 sg13g2_dfrbp_1 _29165_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1332),
    .D(_01503_),
    .Q_N(_12585_),
    .Q(\atari2600.ram[8][3] ));
 sg13g2_dfrbp_1 _29166_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1331),
    .D(_01504_),
    .Q_N(_12584_),
    .Q(\atari2600.ram[8][4] ));
 sg13g2_dfrbp_1 _29167_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1330),
    .D(_01505_),
    .Q_N(_12583_),
    .Q(\atari2600.ram[8][5] ));
 sg13g2_dfrbp_1 _29168_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1329),
    .D(_01506_),
    .Q_N(_12582_),
    .Q(\atari2600.ram[8][6] ));
 sg13g2_dfrbp_1 _29169_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1324),
    .D(_01507_),
    .Q_N(_13871_),
    .Q(\atari2600.ram[8][7] ));
 sg13g2_dfrbp_1 _29170_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1328),
    .D(net7596),
    .Q_N(_12581_),
    .Q(\hvsync_gen.vga.vsync ));
 sg13g2_dfrbp_1 _29171_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1327),
    .D(net2936),
    .Q_N(_00168_),
    .Q(\hvsync_gen.vga.vpos[0] ));
 sg13g2_dfrbp_1 _29172_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1326),
    .D(net7322),
    .Q_N(_12580_),
    .Q(\hvsync_gen.vga.vpos[1] ));
 sg13g2_dfrbp_1 _29173_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1325),
    .D(_01510_),
    .Q_N(_12579_),
    .Q(\hvsync_gen.vga.vpos[2] ));
 sg13g2_dfrbp_1 _29174_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1323),
    .D(_01511_),
    .Q_N(_12578_),
    .Q(\hvsync_gen.vga.vpos[3] ));
 sg13g2_dfrbp_1 _29175_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1322),
    .D(_01512_),
    .Q_N(_12577_),
    .Q(\hvsync_gen.vga.vpos[4] ));
 sg13g2_dfrbp_1 _29176_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1321),
    .D(net7180),
    .Q_N(_12576_),
    .Q(\hvsync_gen.vga.vpos[5] ));
 sg13g2_dfrbp_1 _29177_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1320),
    .D(_01514_),
    .Q_N(_12575_),
    .Q(\hvsync_gen.vga.vpos[6] ));
 sg13g2_dfrbp_1 _29178_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1319),
    .D(_01515_),
    .Q_N(_12574_),
    .Q(\hvsync_gen.vga.vpos[7] ));
 sg13g2_dfrbp_1 _29179_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1317),
    .D(_01516_),
    .Q_N(_12573_),
    .Q(\hvsync_gen.vga.vpos[8] ));
 sg13g2_dfrbp_1 _29180_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1583),
    .D(net7132),
    .Q_N(_13872_),
    .Q(\hvsync_gen.vga.vpos[9] ));
 sg13g2_dfrbp_1 _29181_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1316),
    .D(_00055_),
    .Q_N(_12572_),
    .Q(hsync));
 sg13g2_dfrbp_1 _29182_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1315),
    .D(_01518_),
    .Q_N(_12571_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _29183_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1314),
    .D(_01519_),
    .Q_N(_12570_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _29184_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1313),
    .D(_01520_),
    .Q_N(_12569_),
    .Q(\atari2600.ram[23][0] ));
 sg13g2_dfrbp_1 _29185_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1312),
    .D(_01521_),
    .Q_N(_12568_),
    .Q(\atari2600.ram[23][1] ));
 sg13g2_dfrbp_1 _29186_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1311),
    .D(_01522_),
    .Q_N(_12567_),
    .Q(\atari2600.ram[23][2] ));
 sg13g2_dfrbp_1 _29187_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1310),
    .D(_01523_),
    .Q_N(_12566_),
    .Q(\atari2600.ram[23][3] ));
 sg13g2_dfrbp_1 _29188_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1309),
    .D(_01524_),
    .Q_N(_12565_),
    .Q(\atari2600.ram[23][4] ));
 sg13g2_dfrbp_1 _29189_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1308),
    .D(_01525_),
    .Q_N(_12564_),
    .Q(\atari2600.ram[23][5] ));
 sg13g2_dfrbp_1 _29190_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1307),
    .D(_01526_),
    .Q_N(_12563_),
    .Q(\atari2600.ram[23][6] ));
 sg13g2_dfrbp_1 _29191_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1306),
    .D(_01527_),
    .Q_N(_12562_),
    .Q(\atari2600.ram[23][7] ));
 sg13g2_dfrbp_1 _29192_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1305),
    .D(_01528_),
    .Q_N(_12561_),
    .Q(\atari2600.ram[33][0] ));
 sg13g2_dfrbp_1 _29193_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1304),
    .D(_01529_),
    .Q_N(_12560_),
    .Q(\atari2600.ram[33][1] ));
 sg13g2_dfrbp_1 _29194_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1303),
    .D(_01530_),
    .Q_N(_12559_),
    .Q(\atari2600.ram[33][2] ));
 sg13g2_dfrbp_1 _29195_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1302),
    .D(_01531_),
    .Q_N(_12558_),
    .Q(\atari2600.ram[33][3] ));
 sg13g2_dfrbp_1 _29196_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1301),
    .D(_01532_),
    .Q_N(_12557_),
    .Q(\atari2600.ram[33][4] ));
 sg13g2_dfrbp_1 _29197_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1300),
    .D(_01533_),
    .Q_N(_12556_),
    .Q(\atari2600.ram[33][5] ));
 sg13g2_dfrbp_1 _29198_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net1299),
    .D(_01534_),
    .Q_N(_12555_),
    .Q(\atari2600.ram[33][6] ));
 sg13g2_dfrbp_1 _29199_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1298),
    .D(_01535_),
    .Q_N(_12554_),
    .Q(\atari2600.ram[33][7] ));
 sg13g2_dfrbp_1 _29200_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1297),
    .D(_01536_),
    .Q_N(_12553_),
    .Q(\atari2600.ram[28][0] ));
 sg13g2_dfrbp_1 _29201_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1296),
    .D(_01537_),
    .Q_N(_12552_),
    .Q(\atari2600.ram[28][1] ));
 sg13g2_dfrbp_1 _29202_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1295),
    .D(_01538_),
    .Q_N(_12551_),
    .Q(\atari2600.ram[28][2] ));
 sg13g2_dfrbp_1 _29203_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1294),
    .D(_01539_),
    .Q_N(_12550_),
    .Q(\atari2600.ram[28][3] ));
 sg13g2_dfrbp_1 _29204_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1293),
    .D(_01540_),
    .Q_N(_12549_),
    .Q(\atari2600.ram[28][4] ));
 sg13g2_dfrbp_1 _29205_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1292),
    .D(_01541_),
    .Q_N(_12548_),
    .Q(\atari2600.ram[28][5] ));
 sg13g2_dfrbp_1 _29206_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1291),
    .D(_01542_),
    .Q_N(_12547_),
    .Q(\atari2600.ram[28][6] ));
 sg13g2_dfrbp_1 _29207_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1290),
    .D(_01543_),
    .Q_N(_12546_),
    .Q(\atari2600.ram[28][7] ));
 sg13g2_dfrbp_1 _29208_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1289),
    .D(_01544_),
    .Q_N(_12545_),
    .Q(\atari2600.ram[34][0] ));
 sg13g2_dfrbp_1 _29209_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1286),
    .D(_01545_),
    .Q_N(_12544_),
    .Q(\atari2600.ram[34][1] ));
 sg13g2_dfrbp_1 _29210_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1285),
    .D(_01546_),
    .Q_N(_12543_),
    .Q(\atari2600.ram[34][2] ));
 sg13g2_dfrbp_1 _29211_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1284),
    .D(_01547_),
    .Q_N(_12542_),
    .Q(\atari2600.ram[34][3] ));
 sg13g2_dfrbp_1 _29212_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1283),
    .D(_01548_),
    .Q_N(_12541_),
    .Q(\atari2600.ram[34][4] ));
 sg13g2_dfrbp_1 _29213_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1282),
    .D(_01549_),
    .Q_N(_12540_),
    .Q(\atari2600.ram[34][5] ));
 sg13g2_dfrbp_1 _29214_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net1281),
    .D(_01550_),
    .Q_N(_12539_),
    .Q(\atari2600.ram[34][6] ));
 sg13g2_dfrbp_1 _29215_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1280),
    .D(_01551_),
    .Q_N(_12538_),
    .Q(\atari2600.ram[34][7] ));
 sg13g2_dfrbp_1 _29216_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1279),
    .D(net3226),
    .Q_N(_12537_),
    .Q(\gamepad_pmod.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _29217_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1278),
    .D(_01553_),
    .Q_N(_12536_),
    .Q(\gamepad_pmod.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _29218_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1277),
    .D(net4422),
    .Q_N(_12535_),
    .Q(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _29219_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1276),
    .D(net4808),
    .Q_N(_12534_),
    .Q(\gamepad_pmod.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _29220_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1275),
    .D(net3787),
    .Q_N(_12533_),
    .Q(\gamepad_pmod.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _29221_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1274),
    .D(net4451),
    .Q_N(_12532_),
    .Q(\gamepad_pmod.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _29222_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1273),
    .D(net4104),
    .Q_N(_12531_),
    .Q(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _29223_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1272),
    .D(net4351),
    .Q_N(_12530_),
    .Q(\gamepad_pmod.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _29224_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1271),
    .D(net4484),
    .Q_N(_12529_),
    .Q(\gamepad_pmod.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _29225_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1270),
    .D(net6846),
    .Q_N(_12528_),
    .Q(\gamepad_pmod.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _29226_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1269),
    .D(net4432),
    .Q_N(_12527_),
    .Q(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _29227_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1268),
    .D(net3423),
    .Q_N(_12526_),
    .Q(\gamepad_pmod.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _29228_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1267),
    .D(_01564_),
    .Q_N(_12525_),
    .Q(\atari2600.ram[27][0] ));
 sg13g2_dfrbp_1 _29229_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1266),
    .D(_01565_),
    .Q_N(_12524_),
    .Q(\atari2600.ram[27][1] ));
 sg13g2_dfrbp_1 _29230_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1265),
    .D(_01566_),
    .Q_N(_12523_),
    .Q(\atari2600.ram[27][2] ));
 sg13g2_dfrbp_1 _29231_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1264),
    .D(_01567_),
    .Q_N(_12522_),
    .Q(\atari2600.ram[27][3] ));
 sg13g2_dfrbp_1 _29232_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1263),
    .D(_01568_),
    .Q_N(_12521_),
    .Q(\atari2600.ram[27][4] ));
 sg13g2_dfrbp_1 _29233_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1262),
    .D(_01569_),
    .Q_N(_12520_),
    .Q(\atari2600.ram[27][5] ));
 sg13g2_dfrbp_1 _29234_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1261),
    .D(_01570_),
    .Q_N(_12519_),
    .Q(\atari2600.ram[27][6] ));
 sg13g2_dfrbp_1 _29235_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1260),
    .D(_01571_),
    .Q_N(_12518_),
    .Q(\atari2600.ram[27][7] ));
 sg13g2_dfrbp_1 _29236_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1259),
    .D(_01572_),
    .Q_N(_12517_),
    .Q(\atari2600.ram[31][0] ));
 sg13g2_dfrbp_1 _29237_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1258),
    .D(_01573_),
    .Q_N(_12516_),
    .Q(\atari2600.ram[31][1] ));
 sg13g2_dfrbp_1 _29238_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1257),
    .D(_01574_),
    .Q_N(_12515_),
    .Q(\atari2600.ram[31][2] ));
 sg13g2_dfrbp_1 _29239_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1256),
    .D(_01575_),
    .Q_N(_12514_),
    .Q(\atari2600.ram[31][3] ));
 sg13g2_dfrbp_1 _29240_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1255),
    .D(_01576_),
    .Q_N(_12513_),
    .Q(\atari2600.ram[31][4] ));
 sg13g2_dfrbp_1 _29241_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1254),
    .D(_01577_),
    .Q_N(_12512_),
    .Q(\atari2600.ram[31][5] ));
 sg13g2_dfrbp_1 _29242_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1253),
    .D(_01578_),
    .Q_N(_12511_),
    .Q(\atari2600.ram[31][6] ));
 sg13g2_dfrbp_1 _29243_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1252),
    .D(_01579_),
    .Q_N(_12510_),
    .Q(\atari2600.ram[31][7] ));
 sg13g2_dfrbp_1 _29244_ (.CLK(clknet_leaf_364_clk),
    .RESET_B(net1251),
    .D(_01580_),
    .Q_N(_12509_),
    .Q(\atari2600.ram[36][0] ));
 sg13g2_dfrbp_1 _29245_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1250),
    .D(_01581_),
    .Q_N(_12508_),
    .Q(\atari2600.ram[36][1] ));
 sg13g2_dfrbp_1 _29246_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1249),
    .D(_01582_),
    .Q_N(_12507_),
    .Q(\atari2600.ram[36][2] ));
 sg13g2_dfrbp_1 _29247_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1248),
    .D(_01583_),
    .Q_N(_12506_),
    .Q(\atari2600.ram[36][3] ));
 sg13g2_dfrbp_1 _29248_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1247),
    .D(_01584_),
    .Q_N(_12505_),
    .Q(\atari2600.ram[36][4] ));
 sg13g2_dfrbp_1 _29249_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1246),
    .D(_01585_),
    .Q_N(_12504_),
    .Q(\atari2600.ram[36][5] ));
 sg13g2_dfrbp_1 _29250_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1245),
    .D(_01586_),
    .Q_N(_12503_),
    .Q(\atari2600.ram[36][6] ));
 sg13g2_dfrbp_1 _29251_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1244),
    .D(_01587_),
    .Q_N(_12502_),
    .Q(\atari2600.ram[36][7] ));
 sg13g2_dfrbp_1 _29252_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1243),
    .D(_01588_),
    .Q_N(_12501_),
    .Q(\atari2600.cpu.AXYS[2][0] ));
 sg13g2_dfrbp_1 _29253_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1242),
    .D(_01589_),
    .Q_N(_12500_),
    .Q(\atari2600.cpu.AXYS[2][1] ));
 sg13g2_dfrbp_1 _29254_ (.CLK(clknet_leaf_365_clk),
    .RESET_B(net1241),
    .D(_01590_),
    .Q_N(_12499_),
    .Q(\atari2600.cpu.AXYS[2][2] ));
 sg13g2_dfrbp_1 _29255_ (.CLK(clknet_leaf_365_clk),
    .RESET_B(net1240),
    .D(_01591_),
    .Q_N(_12498_),
    .Q(\atari2600.cpu.AXYS[2][3] ));
 sg13g2_dfrbp_1 _29256_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1239),
    .D(net3895),
    .Q_N(_12497_),
    .Q(\atari2600.cpu.AXYS[2][4] ));
 sg13g2_dfrbp_1 _29257_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1238),
    .D(_01593_),
    .Q_N(_12496_),
    .Q(\atari2600.cpu.AXYS[2][5] ));
 sg13g2_dfrbp_1 _29258_ (.CLK(clknet_leaf_365_clk),
    .RESET_B(net1237),
    .D(_01594_),
    .Q_N(_12495_),
    .Q(\atari2600.cpu.AXYS[2][6] ));
 sg13g2_dfrbp_1 _29259_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1236),
    .D(_01595_),
    .Q_N(_12494_),
    .Q(\atari2600.cpu.AXYS[2][7] ));
 sg13g2_dfrbp_1 _29260_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1235),
    .D(_01596_),
    .Q_N(_12493_),
    .Q(\atari2600.cpu.AXYS[1][0] ));
 sg13g2_dfrbp_1 _29261_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1234),
    .D(_01597_),
    .Q_N(_12492_),
    .Q(\atari2600.cpu.AXYS[1][1] ));
 sg13g2_dfrbp_1 _29262_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1233),
    .D(_01598_),
    .Q_N(_12491_),
    .Q(\atari2600.cpu.AXYS[1][2] ));
 sg13g2_dfrbp_1 _29263_ (.CLK(clknet_leaf_365_clk),
    .RESET_B(net1232),
    .D(_01599_),
    .Q_N(_12490_),
    .Q(\atari2600.cpu.AXYS[1][3] ));
 sg13g2_dfrbp_1 _29264_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1231),
    .D(net3438),
    .Q_N(_12489_),
    .Q(\atari2600.cpu.AXYS[1][4] ));
 sg13g2_dfrbp_1 _29265_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1230),
    .D(_01601_),
    .Q_N(_12488_),
    .Q(\atari2600.cpu.AXYS[1][5] ));
 sg13g2_dfrbp_1 _29266_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1229),
    .D(_01602_),
    .Q_N(_12487_),
    .Q(\atari2600.cpu.AXYS[1][6] ));
 sg13g2_dfrbp_1 _29267_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1228),
    .D(_01603_),
    .Q_N(_12486_),
    .Q(\atari2600.cpu.AXYS[1][7] ));
 sg13g2_dfrbp_1 _29268_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1227),
    .D(_01604_),
    .Q_N(_12485_),
    .Q(\atari2600.ram[54][0] ));
 sg13g2_dfrbp_1 _29269_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net1226),
    .D(_01605_),
    .Q_N(_12484_),
    .Q(\atari2600.ram[54][1] ));
 sg13g2_dfrbp_1 _29270_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1225),
    .D(_01606_),
    .Q_N(_12483_),
    .Q(\atari2600.ram[54][2] ));
 sg13g2_dfrbp_1 _29271_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1224),
    .D(_01607_),
    .Q_N(_12482_),
    .Q(\atari2600.ram[54][3] ));
 sg13g2_dfrbp_1 _29272_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1223),
    .D(_01608_),
    .Q_N(_12481_),
    .Q(\atari2600.ram[54][4] ));
 sg13g2_dfrbp_1 _29273_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1222),
    .D(_01609_),
    .Q_N(_12480_),
    .Q(\atari2600.ram[54][5] ));
 sg13g2_dfrbp_1 _29274_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1221),
    .D(_01610_),
    .Q_N(_12479_),
    .Q(\atari2600.ram[54][6] ));
 sg13g2_dfrbp_1 _29275_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1220),
    .D(_01611_),
    .Q_N(_12478_),
    .Q(\atari2600.ram[54][7] ));
 sg13g2_dfrbp_1 _29276_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1219),
    .D(_01612_),
    .Q_N(_12477_),
    .Q(\atari2600.ram[55][0] ));
 sg13g2_dfrbp_1 _29277_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1218),
    .D(_01613_),
    .Q_N(_12476_),
    .Q(\atari2600.ram[55][1] ));
 sg13g2_dfrbp_1 _29278_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1217),
    .D(_01614_),
    .Q_N(_12475_),
    .Q(\atari2600.ram[55][2] ));
 sg13g2_dfrbp_1 _29279_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1216),
    .D(_01615_),
    .Q_N(_12474_),
    .Q(\atari2600.ram[55][3] ));
 sg13g2_dfrbp_1 _29280_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net1215),
    .D(_01616_),
    .Q_N(_12473_),
    .Q(\atari2600.ram[55][4] ));
 sg13g2_dfrbp_1 _29281_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1214),
    .D(_01617_),
    .Q_N(_12472_),
    .Q(\atari2600.ram[55][5] ));
 sg13g2_dfrbp_1 _29282_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1213),
    .D(_01618_),
    .Q_N(_12471_),
    .Q(\atari2600.ram[55][6] ));
 sg13g2_dfrbp_1 _29283_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1211),
    .D(_01619_),
    .Q_N(_12470_),
    .Q(\atari2600.ram[55][7] ));
 sg13g2_dfrbp_1 _29284_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1210),
    .D(_01620_),
    .Q_N(_12469_),
    .Q(\atari2600.ram[56][0] ));
 sg13g2_dfrbp_1 _29285_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1209),
    .D(_01621_),
    .Q_N(_12468_),
    .Q(\atari2600.ram[56][1] ));
 sg13g2_dfrbp_1 _29286_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1208),
    .D(_01622_),
    .Q_N(_12467_),
    .Q(\atari2600.ram[56][2] ));
 sg13g2_dfrbp_1 _29287_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1207),
    .D(_01623_),
    .Q_N(_12466_),
    .Q(\atari2600.ram[56][3] ));
 sg13g2_dfrbp_1 _29288_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1206),
    .D(_01624_),
    .Q_N(_12465_),
    .Q(\atari2600.ram[56][4] ));
 sg13g2_dfrbp_1 _29289_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1205),
    .D(_01625_),
    .Q_N(_12464_),
    .Q(\atari2600.ram[56][5] ));
 sg13g2_dfrbp_1 _29290_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1204),
    .D(_01626_),
    .Q_N(_12463_),
    .Q(\atari2600.ram[56][6] ));
 sg13g2_dfrbp_1 _29291_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1203),
    .D(_01627_),
    .Q_N(_12462_),
    .Q(\atari2600.ram[56][7] ));
 sg13g2_dfrbp_1 _29292_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1202),
    .D(_01628_),
    .Q_N(_12461_),
    .Q(\atari2600.ram[57][0] ));
 sg13g2_dfrbp_1 _29293_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1201),
    .D(_01629_),
    .Q_N(_12460_),
    .Q(\atari2600.ram[57][1] ));
 sg13g2_dfrbp_1 _29294_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1200),
    .D(_01630_),
    .Q_N(_12459_),
    .Q(\atari2600.ram[57][2] ));
 sg13g2_dfrbp_1 _29295_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1199),
    .D(_01631_),
    .Q_N(_12458_),
    .Q(\atari2600.ram[57][3] ));
 sg13g2_dfrbp_1 _29296_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1198),
    .D(_01632_),
    .Q_N(_12457_),
    .Q(\atari2600.ram[57][4] ));
 sg13g2_dfrbp_1 _29297_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1197),
    .D(_01633_),
    .Q_N(_12456_),
    .Q(\atari2600.ram[57][5] ));
 sg13g2_dfrbp_1 _29298_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1196),
    .D(_01634_),
    .Q_N(_12455_),
    .Q(\atari2600.ram[57][6] ));
 sg13g2_dfrbp_1 _29299_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1187),
    .D(_01635_),
    .Q_N(_12454_),
    .Q(\atari2600.ram[57][7] ));
 sg13g2_dfrbp_1 _29300_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1186),
    .D(_01636_),
    .Q_N(_12453_),
    .Q(\atari2600.ram[58][0] ));
 sg13g2_dfrbp_1 _29301_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1185),
    .D(_01637_),
    .Q_N(_12452_),
    .Q(\atari2600.ram[58][1] ));
 sg13g2_dfrbp_1 _29302_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1184),
    .D(_01638_),
    .Q_N(_12451_),
    .Q(\atari2600.ram[58][2] ));
 sg13g2_dfrbp_1 _29303_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1183),
    .D(_01639_),
    .Q_N(_12450_),
    .Q(\atari2600.ram[58][3] ));
 sg13g2_dfrbp_1 _29304_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1182),
    .D(_01640_),
    .Q_N(_12449_),
    .Q(\atari2600.ram[58][4] ));
 sg13g2_dfrbp_1 _29305_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1181),
    .D(_01641_),
    .Q_N(_12448_),
    .Q(\atari2600.ram[58][5] ));
 sg13g2_dfrbp_1 _29306_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1180),
    .D(_01642_),
    .Q_N(_12447_),
    .Q(\atari2600.ram[58][6] ));
 sg13g2_dfrbp_1 _29307_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1179),
    .D(_01643_),
    .Q_N(_12446_),
    .Q(\atari2600.ram[58][7] ));
 sg13g2_dfrbp_1 _29308_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1178),
    .D(_01644_),
    .Q_N(_12445_),
    .Q(\atari2600.ram[5][0] ));
 sg13g2_dfrbp_1 _29309_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1177),
    .D(_01645_),
    .Q_N(_12444_),
    .Q(\atari2600.ram[5][1] ));
 sg13g2_dfrbp_1 _29310_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1176),
    .D(_01646_),
    .Q_N(_12443_),
    .Q(\atari2600.ram[5][2] ));
 sg13g2_dfrbp_1 _29311_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1175),
    .D(_01647_),
    .Q_N(_12442_),
    .Q(\atari2600.ram[5][3] ));
 sg13g2_dfrbp_1 _29312_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1174),
    .D(_01648_),
    .Q_N(_12441_),
    .Q(\atari2600.ram[5][4] ));
 sg13g2_dfrbp_1 _29313_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1173),
    .D(_01649_),
    .Q_N(_12440_),
    .Q(\atari2600.ram[5][5] ));
 sg13g2_dfrbp_1 _29314_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1172),
    .D(_01650_),
    .Q_N(_12439_),
    .Q(\atari2600.ram[5][6] ));
 sg13g2_dfrbp_1 _29315_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1171),
    .D(_01651_),
    .Q_N(_12438_),
    .Q(\atari2600.ram[5][7] ));
 sg13g2_dfrbp_1 _29316_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1170),
    .D(_01652_),
    .Q_N(_12437_),
    .Q(\atari2600.ram[60][0] ));
 sg13g2_dfrbp_1 _29317_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1169),
    .D(_01653_),
    .Q_N(_12436_),
    .Q(\atari2600.ram[60][1] ));
 sg13g2_dfrbp_1 _29318_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1168),
    .D(_01654_),
    .Q_N(_12435_),
    .Q(\atari2600.ram[60][2] ));
 sg13g2_dfrbp_1 _29319_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net1167),
    .D(_01655_),
    .Q_N(_12434_),
    .Q(\atari2600.ram[60][3] ));
 sg13g2_dfrbp_1 _29320_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net1166),
    .D(_01656_),
    .Q_N(_12433_),
    .Q(\atari2600.ram[60][4] ));
 sg13g2_dfrbp_1 _29321_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1165),
    .D(_01657_),
    .Q_N(_12432_),
    .Q(\atari2600.ram[60][5] ));
 sg13g2_dfrbp_1 _29322_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net1164),
    .D(_01658_),
    .Q_N(_12431_),
    .Q(\atari2600.ram[60][6] ));
 sg13g2_dfrbp_1 _29323_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1163),
    .D(_01659_),
    .Q_N(_12430_),
    .Q(\atari2600.ram[60][7] ));
 sg13g2_dfrbp_1 _29324_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1162),
    .D(_01660_),
    .Q_N(_12429_),
    .Q(\atari2600.ram[61][0] ));
 sg13g2_dfrbp_1 _29325_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1161),
    .D(_01661_),
    .Q_N(_12428_),
    .Q(\atari2600.ram[61][1] ));
 sg13g2_dfrbp_1 _29326_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1160),
    .D(_01662_),
    .Q_N(_12427_),
    .Q(\atari2600.ram[61][2] ));
 sg13g2_dfrbp_1 _29327_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net1159),
    .D(_01663_),
    .Q_N(_12426_),
    .Q(\atari2600.ram[61][3] ));
 sg13g2_dfrbp_1 _29328_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net1158),
    .D(_01664_),
    .Q_N(_12425_),
    .Q(\atari2600.ram[61][4] ));
 sg13g2_dfrbp_1 _29329_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1157),
    .D(_01665_),
    .Q_N(_12424_),
    .Q(\atari2600.ram[61][5] ));
 sg13g2_dfrbp_1 _29330_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1156),
    .D(_01666_),
    .Q_N(_12423_),
    .Q(\atari2600.ram[61][6] ));
 sg13g2_dfrbp_1 _29331_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net1155),
    .D(_01667_),
    .Q_N(_12422_),
    .Q(\atari2600.ram[61][7] ));
 sg13g2_dfrbp_1 _29332_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net1150),
    .D(_01668_),
    .Q_N(_12421_),
    .Q(\atari2600.ram[62][0] ));
 sg13g2_dfrbp_1 _29333_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1149),
    .D(_01669_),
    .Q_N(_12420_),
    .Q(\atari2600.ram[62][1] ));
 sg13g2_dfrbp_1 _29334_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1148),
    .D(_01670_),
    .Q_N(_12419_),
    .Q(\atari2600.ram[62][2] ));
 sg13g2_dfrbp_1 _29335_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1147),
    .D(_01671_),
    .Q_N(_12418_),
    .Q(\atari2600.ram[62][3] ));
 sg13g2_dfrbp_1 _29336_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1146),
    .D(_01672_),
    .Q_N(_12417_),
    .Q(\atari2600.ram[62][4] ));
 sg13g2_dfrbp_1 _29337_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net1145),
    .D(_01673_),
    .Q_N(_12416_),
    .Q(\atari2600.ram[62][5] ));
 sg13g2_dfrbp_1 _29338_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net1144),
    .D(_01674_),
    .Q_N(_12415_),
    .Q(\atari2600.ram[62][6] ));
 sg13g2_dfrbp_1 _29339_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net1143),
    .D(_01675_),
    .Q_N(_12414_),
    .Q(\atari2600.ram[62][7] ));
 sg13g2_dfrbp_1 _29340_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1142),
    .D(_01676_),
    .Q_N(_12413_),
    .Q(\atari2600.ram[63][0] ));
 sg13g2_dfrbp_1 _29341_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1141),
    .D(_01677_),
    .Q_N(_12412_),
    .Q(\atari2600.ram[63][1] ));
 sg13g2_dfrbp_1 _29342_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1140),
    .D(_01678_),
    .Q_N(_12411_),
    .Q(\atari2600.ram[63][2] ));
 sg13g2_dfrbp_1 _29343_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1139),
    .D(_01679_),
    .Q_N(_12410_),
    .Q(\atari2600.ram[63][3] ));
 sg13g2_dfrbp_1 _29344_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1138),
    .D(_01680_),
    .Q_N(_12409_),
    .Q(\atari2600.ram[63][4] ));
 sg13g2_dfrbp_1 _29345_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1137),
    .D(_01681_),
    .Q_N(_12408_),
    .Q(\atari2600.ram[63][5] ));
 sg13g2_dfrbp_1 _29346_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1136),
    .D(_01682_),
    .Q_N(_12407_),
    .Q(\atari2600.ram[63][6] ));
 sg13g2_dfrbp_1 _29347_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net1135),
    .D(_01683_),
    .Q_N(_12406_),
    .Q(\atari2600.ram[63][7] ));
 sg13g2_dfrbp_1 _29348_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1134),
    .D(_01684_),
    .Q_N(_12405_),
    .Q(\atari2600.ram[64][0] ));
 sg13g2_dfrbp_1 _29349_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1133),
    .D(_01685_),
    .Q_N(_12404_),
    .Q(\atari2600.ram[64][1] ));
 sg13g2_dfrbp_1 _29350_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1132),
    .D(_01686_),
    .Q_N(_12403_),
    .Q(\atari2600.ram[64][2] ));
 sg13g2_dfrbp_1 _29351_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1131),
    .D(_01687_),
    .Q_N(_12402_),
    .Q(\atari2600.ram[64][3] ));
 sg13g2_dfrbp_1 _29352_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1130),
    .D(_01688_),
    .Q_N(_12401_),
    .Q(\atari2600.ram[64][4] ));
 sg13g2_dfrbp_1 _29353_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1129),
    .D(_01689_),
    .Q_N(_12400_),
    .Q(\atari2600.ram[64][5] ));
 sg13g2_dfrbp_1 _29354_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1128),
    .D(_01690_),
    .Q_N(_12399_),
    .Q(\atari2600.ram[64][6] ));
 sg13g2_dfrbp_1 _29355_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1127),
    .D(_01691_),
    .Q_N(_12398_),
    .Q(\atari2600.ram[64][7] ));
 sg13g2_dfrbp_1 _29356_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1126),
    .D(_01692_),
    .Q_N(_12397_),
    .Q(\atari2600.ram[65][0] ));
 sg13g2_dfrbp_1 _29357_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1125),
    .D(_01693_),
    .Q_N(_12396_),
    .Q(\atari2600.ram[65][1] ));
 sg13g2_dfrbp_1 _29358_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1124),
    .D(_01694_),
    .Q_N(_12395_),
    .Q(\atari2600.ram[65][2] ));
 sg13g2_dfrbp_1 _29359_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1123),
    .D(_01695_),
    .Q_N(_12394_),
    .Q(\atari2600.ram[65][3] ));
 sg13g2_dfrbp_1 _29360_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1122),
    .D(_01696_),
    .Q_N(_12393_),
    .Q(\atari2600.ram[65][4] ));
 sg13g2_dfrbp_1 _29361_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1121),
    .D(_01697_),
    .Q_N(_12392_),
    .Q(\atari2600.ram[65][5] ));
 sg13g2_dfrbp_1 _29362_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1120),
    .D(_01698_),
    .Q_N(_12391_),
    .Q(\atari2600.ram[65][6] ));
 sg13g2_dfrbp_1 _29363_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1119),
    .D(_01699_),
    .Q_N(_12390_),
    .Q(\atari2600.ram[65][7] ));
 sg13g2_dfrbp_1 _29364_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1118),
    .D(_01700_),
    .Q_N(_12389_),
    .Q(\atari2600.ram[66][0] ));
 sg13g2_dfrbp_1 _29365_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1117),
    .D(_01701_),
    .Q_N(_12388_),
    .Q(\atari2600.ram[66][1] ));
 sg13g2_dfrbp_1 _29366_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1116),
    .D(_01702_),
    .Q_N(_12387_),
    .Q(\atari2600.ram[66][2] ));
 sg13g2_dfrbp_1 _29367_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1115),
    .D(_01703_),
    .Q_N(_12386_),
    .Q(\atari2600.ram[66][3] ));
 sg13g2_dfrbp_1 _29368_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1114),
    .D(_01704_),
    .Q_N(_12385_),
    .Q(\atari2600.ram[66][4] ));
 sg13g2_dfrbp_1 _29369_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1113),
    .D(_01705_),
    .Q_N(_12384_),
    .Q(\atari2600.ram[66][5] ));
 sg13g2_dfrbp_1 _29370_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1112),
    .D(_01706_),
    .Q_N(_12383_),
    .Q(\atari2600.ram[66][6] ));
 sg13g2_dfrbp_1 _29371_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1111),
    .D(_01707_),
    .Q_N(_12382_),
    .Q(\atari2600.ram[66][7] ));
 sg13g2_dfrbp_1 _29372_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1110),
    .D(_01708_),
    .Q_N(_12381_),
    .Q(\atari2600.ram[67][0] ));
 sg13g2_dfrbp_1 _29373_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1109),
    .D(_01709_),
    .Q_N(_12380_),
    .Q(\atari2600.ram[67][1] ));
 sg13g2_dfrbp_1 _29374_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1108),
    .D(_01710_),
    .Q_N(_12379_),
    .Q(\atari2600.ram[67][2] ));
 sg13g2_dfrbp_1 _29375_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1107),
    .D(_01711_),
    .Q_N(_12378_),
    .Q(\atari2600.ram[67][3] ));
 sg13g2_dfrbp_1 _29376_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1106),
    .D(_01712_),
    .Q_N(_12377_),
    .Q(\atari2600.ram[67][4] ));
 sg13g2_dfrbp_1 _29377_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1105),
    .D(_01713_),
    .Q_N(_12376_),
    .Q(\atari2600.ram[67][5] ));
 sg13g2_dfrbp_1 _29378_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1104),
    .D(_01714_),
    .Q_N(_12375_),
    .Q(\atari2600.ram[67][6] ));
 sg13g2_dfrbp_1 _29379_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1103),
    .D(_01715_),
    .Q_N(_12374_),
    .Q(\atari2600.ram[67][7] ));
 sg13g2_dfrbp_1 _29380_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1102),
    .D(_01716_),
    .Q_N(_12373_),
    .Q(\atari2600.ram[68][0] ));
 sg13g2_dfrbp_1 _29381_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1101),
    .D(_01717_),
    .Q_N(_12372_),
    .Q(\atari2600.ram[68][1] ));
 sg13g2_dfrbp_1 _29382_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1100),
    .D(_01718_),
    .Q_N(_12371_),
    .Q(\atari2600.ram[68][2] ));
 sg13g2_dfrbp_1 _29383_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1099),
    .D(_01719_),
    .Q_N(_12370_),
    .Q(\atari2600.ram[68][3] ));
 sg13g2_dfrbp_1 _29384_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1098),
    .D(_01720_),
    .Q_N(_12369_),
    .Q(\atari2600.ram[68][4] ));
 sg13g2_dfrbp_1 _29385_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1097),
    .D(_01721_),
    .Q_N(_12368_),
    .Q(\atari2600.ram[68][5] ));
 sg13g2_dfrbp_1 _29386_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1096),
    .D(_01722_),
    .Q_N(_12367_),
    .Q(\atari2600.ram[68][6] ));
 sg13g2_dfrbp_1 _29387_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1095),
    .D(_01723_),
    .Q_N(_12366_),
    .Q(\atari2600.ram[68][7] ));
 sg13g2_dfrbp_1 _29388_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1094),
    .D(_01724_),
    .Q_N(_12365_),
    .Q(\atari2600.ram[6][0] ));
 sg13g2_dfrbp_1 _29389_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1093),
    .D(_01725_),
    .Q_N(_12364_),
    .Q(\atari2600.ram[6][1] ));
 sg13g2_dfrbp_1 _29390_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1092),
    .D(_01726_),
    .Q_N(_12363_),
    .Q(\atari2600.ram[6][2] ));
 sg13g2_dfrbp_1 _29391_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1091),
    .D(_01727_),
    .Q_N(_12362_),
    .Q(\atari2600.ram[6][3] ));
 sg13g2_dfrbp_1 _29392_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1090),
    .D(_01728_),
    .Q_N(_12361_),
    .Q(\atari2600.ram[6][4] ));
 sg13g2_dfrbp_1 _29393_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1089),
    .D(_01729_),
    .Q_N(_12360_),
    .Q(\atari2600.ram[6][5] ));
 sg13g2_dfrbp_1 _29394_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1088),
    .D(_01730_),
    .Q_N(_12359_),
    .Q(\atari2600.ram[6][6] ));
 sg13g2_dfrbp_1 _29395_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1087),
    .D(_01731_),
    .Q_N(_12358_),
    .Q(\atari2600.ram[6][7] ));
 sg13g2_dfrbp_1 _29396_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1086),
    .D(_01732_),
    .Q_N(_12357_),
    .Q(\atari2600.ram[70][0] ));
 sg13g2_dfrbp_1 _29397_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1085),
    .D(_01733_),
    .Q_N(_12356_),
    .Q(\atari2600.ram[70][1] ));
 sg13g2_dfrbp_1 _29398_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1084),
    .D(_01734_),
    .Q_N(_12355_),
    .Q(\atari2600.ram[70][2] ));
 sg13g2_dfrbp_1 _29399_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1083),
    .D(_01735_),
    .Q_N(_12354_),
    .Q(\atari2600.ram[70][3] ));
 sg13g2_dfrbp_1 _29400_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1082),
    .D(_01736_),
    .Q_N(_12353_),
    .Q(\atari2600.ram[70][4] ));
 sg13g2_dfrbp_1 _29401_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1081),
    .D(_01737_),
    .Q_N(_12352_),
    .Q(\atari2600.ram[70][5] ));
 sg13g2_dfrbp_1 _29402_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1080),
    .D(_01738_),
    .Q_N(_12351_),
    .Q(\atari2600.ram[70][6] ));
 sg13g2_dfrbp_1 _29403_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1079),
    .D(_01739_),
    .Q_N(_12350_),
    .Q(\atari2600.ram[70][7] ));
 sg13g2_dfrbp_1 _29404_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1078),
    .D(_01740_),
    .Q_N(_12349_),
    .Q(\atari2600.ram[20][0] ));
 sg13g2_dfrbp_1 _29405_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1077),
    .D(_01741_),
    .Q_N(_12348_),
    .Q(\atari2600.ram[20][1] ));
 sg13g2_dfrbp_1 _29406_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1076),
    .D(_01742_),
    .Q_N(_12347_),
    .Q(\atari2600.ram[20][2] ));
 sg13g2_dfrbp_1 _29407_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1075),
    .D(_01743_),
    .Q_N(_12346_),
    .Q(\atari2600.ram[20][3] ));
 sg13g2_dfrbp_1 _29408_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1074),
    .D(_01744_),
    .Q_N(_12345_),
    .Q(\atari2600.ram[20][4] ));
 sg13g2_dfrbp_1 _29409_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1073),
    .D(_01745_),
    .Q_N(_12344_),
    .Q(\atari2600.ram[20][5] ));
 sg13g2_dfrbp_1 _29410_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1072),
    .D(_01746_),
    .Q_N(_12343_),
    .Q(\atari2600.ram[20][6] ));
 sg13g2_dfrbp_1 _29411_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1071),
    .D(_01747_),
    .Q_N(_12342_),
    .Q(\atari2600.ram[20][7] ));
 sg13g2_dfrbp_1 _29412_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1070),
    .D(_01748_),
    .Q_N(_12341_),
    .Q(\atari2600.ram[1][0] ));
 sg13g2_dfrbp_1 _29413_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1069),
    .D(_01749_),
    .Q_N(_12340_),
    .Q(\atari2600.ram[1][1] ));
 sg13g2_dfrbp_1 _29414_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1068),
    .D(_01750_),
    .Q_N(_12339_),
    .Q(\atari2600.ram[1][2] ));
 sg13g2_dfrbp_1 _29415_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1067),
    .D(_01751_),
    .Q_N(_12338_),
    .Q(\atari2600.ram[1][3] ));
 sg13g2_dfrbp_1 _29416_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1066),
    .D(_01752_),
    .Q_N(_12337_),
    .Q(\atari2600.ram[1][4] ));
 sg13g2_dfrbp_1 _29417_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1065),
    .D(_01753_),
    .Q_N(_12336_),
    .Q(\atari2600.ram[1][5] ));
 sg13g2_dfrbp_1 _29418_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1064),
    .D(_01754_),
    .Q_N(_12335_),
    .Q(\atari2600.ram[1][6] ));
 sg13g2_dfrbp_1 _29419_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1063),
    .D(_01755_),
    .Q_N(_12334_),
    .Q(\atari2600.ram[1][7] ));
 sg13g2_dfrbp_1 _29420_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1062),
    .D(_01756_),
    .Q_N(_12333_),
    .Q(\atari2600.ram[18][0] ));
 sg13g2_dfrbp_1 _29421_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1061),
    .D(_01757_),
    .Q_N(_12332_),
    .Q(\atari2600.ram[18][1] ));
 sg13g2_dfrbp_1 _29422_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1060),
    .D(_01758_),
    .Q_N(_12331_),
    .Q(\atari2600.ram[18][2] ));
 sg13g2_dfrbp_1 _29423_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1059),
    .D(_01759_),
    .Q_N(_12330_),
    .Q(\atari2600.ram[18][3] ));
 sg13g2_dfrbp_1 _29424_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1058),
    .D(_01760_),
    .Q_N(_12329_),
    .Q(\atari2600.ram[18][4] ));
 sg13g2_dfrbp_1 _29425_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1057),
    .D(_01761_),
    .Q_N(_12328_),
    .Q(\atari2600.ram[18][5] ));
 sg13g2_dfrbp_1 _29426_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1056),
    .D(_01762_),
    .Q_N(_12327_),
    .Q(\atari2600.ram[18][6] ));
 sg13g2_dfrbp_1 _29427_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1055),
    .D(_01763_),
    .Q_N(_12326_),
    .Q(\atari2600.ram[18][7] ));
 sg13g2_dfrbp_1 _29428_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1054),
    .D(_01764_),
    .Q_N(_12325_),
    .Q(\atari2600.ram[17][0] ));
 sg13g2_dfrbp_1 _29429_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1053),
    .D(_01765_),
    .Q_N(_12324_),
    .Q(\atari2600.ram[17][1] ));
 sg13g2_dfrbp_1 _29430_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1052),
    .D(_01766_),
    .Q_N(_12323_),
    .Q(\atari2600.ram[17][2] ));
 sg13g2_dfrbp_1 _29431_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1051),
    .D(_01767_),
    .Q_N(_12322_),
    .Q(\atari2600.ram[17][3] ));
 sg13g2_dfrbp_1 _29432_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1050),
    .D(_01768_),
    .Q_N(_12321_),
    .Q(\atari2600.ram[17][4] ));
 sg13g2_dfrbp_1 _29433_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1049),
    .D(_01769_),
    .Q_N(_12320_),
    .Q(\atari2600.ram[17][5] ));
 sg13g2_dfrbp_1 _29434_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1048),
    .D(_01770_),
    .Q_N(_12319_),
    .Q(\atari2600.ram[17][6] ));
 sg13g2_dfrbp_1 _29435_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1047),
    .D(_01771_),
    .Q_N(_12318_),
    .Q(\atari2600.ram[17][7] ));
 sg13g2_dfrbp_1 _29436_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1046),
    .D(_01772_),
    .Q_N(_12317_),
    .Q(\atari2600.address_bus_r[0] ));
 sg13g2_dfrbp_1 _29437_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1045),
    .D(_01773_),
    .Q_N(_12316_),
    .Q(\atari2600.address_bus_r[1] ));
 sg13g2_dfrbp_1 _29438_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1044),
    .D(_01774_),
    .Q_N(_12315_),
    .Q(\atari2600.address_bus_r[2] ));
 sg13g2_dfrbp_1 _29439_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1043),
    .D(_01775_),
    .Q_N(_12314_),
    .Q(\atari2600.address_bus_r[3] ));
 sg13g2_dfrbp_1 _29440_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1042),
    .D(_01776_),
    .Q_N(_12313_),
    .Q(\atari2600.address_bus_r[4] ));
 sg13g2_dfrbp_1 _29441_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1041),
    .D(_01777_),
    .Q_N(_12312_),
    .Q(\atari2600.address_bus_r[5] ));
 sg13g2_dfrbp_1 _29442_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1040),
    .D(_01778_),
    .Q_N(_12311_),
    .Q(\atari2600.address_bus_r[6] ));
 sg13g2_dfrbp_1 _29443_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1039),
    .D(_01779_),
    .Q_N(_12310_),
    .Q(\atari2600.address_bus_r[7] ));
 sg13g2_dfrbp_1 _29444_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1038),
    .D(_01780_),
    .Q_N(_12309_),
    .Q(\atari2600.address_bus_r[8] ));
 sg13g2_dfrbp_1 _29445_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1037),
    .D(_01781_),
    .Q_N(_12308_),
    .Q(\atari2600.address_bus_r[9] ));
 sg13g2_dfrbp_1 _29446_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1036),
    .D(_01782_),
    .Q_N(_12307_),
    .Q(\atari2600.address_bus_r[10] ));
 sg13g2_dfrbp_1 _29447_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1035),
    .D(_01783_),
    .Q_N(_12306_),
    .Q(\atari2600.address_bus_r[11] ));
 sg13g2_dfrbp_1 _29448_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1034),
    .D(_01784_),
    .Q_N(_12305_),
    .Q(\atari2600.address_bus_r[12] ));
 sg13g2_dfrbp_1 _29449_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1033),
    .D(_01785_),
    .Q_N(_12304_),
    .Q(\atari2600.ram[16][0] ));
 sg13g2_dfrbp_1 _29450_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1032),
    .D(_01786_),
    .Q_N(_12303_),
    .Q(\atari2600.ram[16][1] ));
 sg13g2_dfrbp_1 _29451_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1031),
    .D(_01787_),
    .Q_N(_12302_),
    .Q(\atari2600.ram[16][2] ));
 sg13g2_dfrbp_1 _29452_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1030),
    .D(_01788_),
    .Q_N(_12301_),
    .Q(\atari2600.ram[16][3] ));
 sg13g2_dfrbp_1 _29453_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1029),
    .D(_01789_),
    .Q_N(_12300_),
    .Q(\atari2600.ram[16][4] ));
 sg13g2_dfrbp_1 _29454_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1028),
    .D(_01790_),
    .Q_N(_12299_),
    .Q(\atari2600.ram[16][5] ));
 sg13g2_dfrbp_1 _29455_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1027),
    .D(_01791_),
    .Q_N(_12298_),
    .Q(\atari2600.ram[16][6] ));
 sg13g2_dfrbp_1 _29456_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1026),
    .D(_01792_),
    .Q_N(_12297_),
    .Q(\atari2600.ram[16][7] ));
 sg13g2_dfrbp_1 _29457_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1025),
    .D(_01793_),
    .Q_N(_12296_),
    .Q(\atari2600.ram[15][0] ));
 sg13g2_dfrbp_1 _29458_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1024),
    .D(_01794_),
    .Q_N(_12295_),
    .Q(\atari2600.ram[15][1] ));
 sg13g2_dfrbp_1 _29459_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1023),
    .D(_01795_),
    .Q_N(_12294_),
    .Q(\atari2600.ram[15][2] ));
 sg13g2_dfrbp_1 _29460_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1022),
    .D(_01796_),
    .Q_N(_12293_),
    .Q(\atari2600.ram[15][3] ));
 sg13g2_dfrbp_1 _29461_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1021),
    .D(_01797_),
    .Q_N(_12292_),
    .Q(\atari2600.ram[15][4] ));
 sg13g2_dfrbp_1 _29462_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1020),
    .D(_01798_),
    .Q_N(_12291_),
    .Q(\atari2600.ram[15][5] ));
 sg13g2_dfrbp_1 _29463_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1019),
    .D(_01799_),
    .Q_N(_12290_),
    .Q(\atari2600.ram[15][6] ));
 sg13g2_dfrbp_1 _29464_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1018),
    .D(_01800_),
    .Q_N(_12289_),
    .Q(\atari2600.ram[15][7] ));
 sg13g2_dfrbp_1 _29465_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1017),
    .D(_01801_),
    .Q_N(_12288_),
    .Q(\atari2600.ram[14][0] ));
 sg13g2_dfrbp_1 _29466_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1016),
    .D(_01802_),
    .Q_N(_12287_),
    .Q(\atari2600.ram[14][1] ));
 sg13g2_dfrbp_1 _29467_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1015),
    .D(_01803_),
    .Q_N(_12286_),
    .Q(\atari2600.ram[14][2] ));
 sg13g2_dfrbp_1 _29468_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1014),
    .D(_01804_),
    .Q_N(_12285_),
    .Q(\atari2600.ram[14][3] ));
 sg13g2_dfrbp_1 _29469_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1013),
    .D(_01805_),
    .Q_N(_12284_),
    .Q(\atari2600.ram[14][4] ));
 sg13g2_dfrbp_1 _29470_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1012),
    .D(_01806_),
    .Q_N(_12283_),
    .Q(\atari2600.ram[14][5] ));
 sg13g2_dfrbp_1 _29471_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1011),
    .D(_01807_),
    .Q_N(_12282_),
    .Q(\atari2600.ram[14][6] ));
 sg13g2_dfrbp_1 _29472_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1584),
    .D(_01808_),
    .Q_N(_13873_),
    .Q(\atari2600.ram[14][7] ));
 sg13g2_dfrbp_1 _29473_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1585),
    .D(_00001_),
    .Q_N(_13874_),
    .Q(\atari2600.ram_data[0] ));
 sg13g2_dfrbp_1 _29474_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1586),
    .D(_00002_),
    .Q_N(_13875_),
    .Q(\atari2600.ram_data[1] ));
 sg13g2_dfrbp_1 _29475_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1587),
    .D(_00003_),
    .Q_N(_13876_),
    .Q(\atari2600.ram_data[2] ));
 sg13g2_dfrbp_1 _29476_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1588),
    .D(_00004_),
    .Q_N(_13877_),
    .Q(\atari2600.ram_data[3] ));
 sg13g2_dfrbp_1 _29477_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1589),
    .D(_00005_),
    .Q_N(_13878_),
    .Q(\atari2600.ram_data[4] ));
 sg13g2_dfrbp_1 _29478_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1590),
    .D(_00006_),
    .Q_N(_13879_),
    .Q(\atari2600.ram_data[5] ));
 sg13g2_dfrbp_1 _29479_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net989),
    .D(_00007_),
    .Q_N(_13880_),
    .Q(\atari2600.ram_data[6] ));
 sg13g2_dfrbp_1 _29480_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1010),
    .D(_00008_),
    .Q_N(_12281_),
    .Q(\atari2600.ram_data[7] ));
 sg13g2_dfrbp_1 _29481_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1009),
    .D(net7394),
    .Q_N(_12280_),
    .Q(\flash_rom.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _29482_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1008),
    .D(net7476),
    .Q_N(_12279_),
    .Q(\flash_rom.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _29483_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1006),
    .D(_01811_),
    .Q_N(_12278_),
    .Q(\flash_rom.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _29484_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1004),
    .D(net4156),
    .Q_N(_00132_),
    .Q(\flash_rom.fsm_state[0] ));
 sg13g2_dfrbp_1 _29485_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1002),
    .D(_01813_),
    .Q_N(_12277_),
    .Q(\flash_rom.fsm_state[1] ));
 sg13g2_dfrbp_1 _29486_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1000),
    .D(_01814_),
    .Q_N(_00094_),
    .Q(\flash_rom.fsm_state[2] ));
 sg13g2_dfrbp_1 _29487_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net998),
    .D(_01815_),
    .Q_N(_12276_),
    .Q(\external_rom_data[0] ));
 sg13g2_dfrbp_1 _29488_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net997),
    .D(net7403),
    .Q_N(_12275_),
    .Q(\external_rom_data[1] ));
 sg13g2_dfrbp_1 _29489_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net996),
    .D(_01817_),
    .Q_N(_12274_),
    .Q(\external_rom_data[2] ));
 sg13g2_dfrbp_1 _29490_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net995),
    .D(_01818_),
    .Q_N(_12273_),
    .Q(\external_rom_data[3] ));
 sg13g2_dfrbp_1 _29491_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net994),
    .D(net3489),
    .Q_N(_12272_),
    .Q(\external_rom_data[4] ));
 sg13g2_dfrbp_1 _29492_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net993),
    .D(net3357),
    .Q_N(_12271_),
    .Q(\external_rom_data[5] ));
 sg13g2_dfrbp_1 _29493_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net992),
    .D(net4166),
    .Q_N(_12270_),
    .Q(\external_rom_data[6] ));
 sg13g2_dfrbp_1 _29494_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net991),
    .D(net4381),
    .Q_N(_12269_),
    .Q(\external_rom_data[7] ));
 sg13g2_dfrbp_1 _29495_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net990),
    .D(_01823_),
    .Q_N(_00112_),
    .Q(\flash_rom.spi_clk_out ));
 sg13g2_dfrbp_1 _29496_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net988),
    .D(net7298),
    .Q_N(_12268_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _29497_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net986),
    .D(net7305),
    .Q_N(_12267_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _29498_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net984),
    .D(_01826_),
    .Q_N(_12266_),
    .Q(\atari2600.tia.p1_spacing[4] ));
 sg13g2_dfrbp_1 _29499_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net982),
    .D(_01827_),
    .Q_N(_12265_),
    .Q(\atari2600.tia.p1_spacing[5] ));
 sg13g2_dfrbp_1 _29500_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net980),
    .D(_01828_),
    .Q_N(_12264_),
    .Q(\atari2600.tia.p1_spacing[6] ));
 sg13g2_dfrbp_1 _29501_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net963),
    .D(_01829_),
    .Q_N(_12263_),
    .Q(\atari2600.ram[42][0] ));
 sg13g2_dfrbp_1 _29502_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net962),
    .D(_01830_),
    .Q_N(_12262_),
    .Q(\atari2600.ram[42][1] ));
 sg13g2_dfrbp_1 _29503_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net961),
    .D(_01831_),
    .Q_N(_12261_),
    .Q(\atari2600.ram[42][2] ));
 sg13g2_dfrbp_1 _29504_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net960),
    .D(_01832_),
    .Q_N(_12260_),
    .Q(\atari2600.ram[42][3] ));
 sg13g2_dfrbp_1 _29505_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net959),
    .D(_01833_),
    .Q_N(_12259_),
    .Q(\atari2600.ram[42][4] ));
 sg13g2_dfrbp_1 _29506_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net958),
    .D(_01834_),
    .Q_N(_12258_),
    .Q(\atari2600.ram[42][5] ));
 sg13g2_dfrbp_1 _29507_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net957),
    .D(_01835_),
    .Q_N(_12257_),
    .Q(\atari2600.ram[42][6] ));
 sg13g2_dfrbp_1 _29508_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net956),
    .D(_01836_),
    .Q_N(_12256_),
    .Q(\atari2600.ram[42][7] ));
 sg13g2_dfrbp_1 _29509_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net955),
    .D(_01837_),
    .Q_N(_12255_),
    .Q(\atari2600.ram[43][0] ));
 sg13g2_dfrbp_1 _29510_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net954),
    .D(_01838_),
    .Q_N(_12254_),
    .Q(\atari2600.ram[43][1] ));
 sg13g2_dfrbp_1 _29511_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net953),
    .D(_01839_),
    .Q_N(_12253_),
    .Q(\atari2600.ram[43][2] ));
 sg13g2_dfrbp_1 _29512_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net952),
    .D(_01840_),
    .Q_N(_12252_),
    .Q(\atari2600.ram[43][3] ));
 sg13g2_dfrbp_1 _29513_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net951),
    .D(_01841_),
    .Q_N(_12251_),
    .Q(\atari2600.ram[43][4] ));
 sg13g2_dfrbp_1 _29514_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net950),
    .D(_01842_),
    .Q_N(_12250_),
    .Q(\atari2600.ram[43][5] ));
 sg13g2_dfrbp_1 _29515_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net949),
    .D(_01843_),
    .Q_N(_12249_),
    .Q(\atari2600.ram[43][6] ));
 sg13g2_dfrbp_1 _29516_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net948),
    .D(_01844_),
    .Q_N(_12248_),
    .Q(\atari2600.ram[43][7] ));
 sg13g2_dfrbp_1 _29517_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net947),
    .D(_01845_),
    .Q_N(_12247_),
    .Q(\atari2600.ram[41][0] ));
 sg13g2_dfrbp_1 _29518_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net946),
    .D(_01846_),
    .Q_N(_12246_),
    .Q(\atari2600.ram[41][1] ));
 sg13g2_dfrbp_1 _29519_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net945),
    .D(_01847_),
    .Q_N(_12245_),
    .Q(\atari2600.ram[41][2] ));
 sg13g2_dfrbp_1 _29520_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net944),
    .D(_01848_),
    .Q_N(_12244_),
    .Q(\atari2600.ram[41][3] ));
 sg13g2_dfrbp_1 _29521_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net943),
    .D(_01849_),
    .Q_N(_12243_),
    .Q(\atari2600.ram[41][4] ));
 sg13g2_dfrbp_1 _29522_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net942),
    .D(_01850_),
    .Q_N(_12242_),
    .Q(\atari2600.ram[41][5] ));
 sg13g2_dfrbp_1 _29523_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net941),
    .D(_01851_),
    .Q_N(_12241_),
    .Q(\atari2600.ram[41][6] ));
 sg13g2_dfrbp_1 _29524_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net940),
    .D(_01852_),
    .Q_N(_12240_),
    .Q(\atari2600.ram[41][7] ));
 sg13g2_dfrbp_1 _29525_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net939),
    .D(_01853_),
    .Q_N(_12239_),
    .Q(\atari2600.ram[40][0] ));
 sg13g2_dfrbp_1 _29526_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net938),
    .D(_01854_),
    .Q_N(_12238_),
    .Q(\atari2600.ram[40][1] ));
 sg13g2_dfrbp_1 _29527_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net937),
    .D(_01855_),
    .Q_N(_12237_),
    .Q(\atari2600.ram[40][2] ));
 sg13g2_dfrbp_1 _29528_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net936),
    .D(_01856_),
    .Q_N(_12236_),
    .Q(\atari2600.ram[40][3] ));
 sg13g2_dfrbp_1 _29529_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net935),
    .D(_01857_),
    .Q_N(_12235_),
    .Q(\atari2600.ram[40][4] ));
 sg13g2_dfrbp_1 _29530_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net934),
    .D(_01858_),
    .Q_N(_12234_),
    .Q(\atari2600.ram[40][5] ));
 sg13g2_dfrbp_1 _29531_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net933),
    .D(_01859_),
    .Q_N(_12233_),
    .Q(\atari2600.ram[40][6] ));
 sg13g2_dfrbp_1 _29532_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net932),
    .D(_01860_),
    .Q_N(_12232_),
    .Q(\atari2600.ram[40][7] ));
 sg13g2_dfrbp_1 _29533_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net931),
    .D(_01861_),
    .Q_N(_12231_),
    .Q(\atari2600.ram[3][0] ));
 sg13g2_dfrbp_1 _29534_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net930),
    .D(_01862_),
    .Q_N(_12230_),
    .Q(\atari2600.ram[3][1] ));
 sg13g2_dfrbp_1 _29535_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net929),
    .D(_01863_),
    .Q_N(_12229_),
    .Q(\atari2600.ram[3][2] ));
 sg13g2_dfrbp_1 _29536_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net928),
    .D(_01864_),
    .Q_N(_12228_),
    .Q(\atari2600.ram[3][3] ));
 sg13g2_dfrbp_1 _29537_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net927),
    .D(_01865_),
    .Q_N(_12227_),
    .Q(\atari2600.ram[3][4] ));
 sg13g2_dfrbp_1 _29538_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net926),
    .D(_01866_),
    .Q_N(_12226_),
    .Q(\atari2600.ram[3][5] ));
 sg13g2_dfrbp_1 _29539_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net925),
    .D(_01867_),
    .Q_N(_12225_),
    .Q(\atari2600.ram[3][6] ));
 sg13g2_dfrbp_1 _29540_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net924),
    .D(_01868_),
    .Q_N(_12224_),
    .Q(\atari2600.ram[3][7] ));
 sg13g2_dfrbp_1 _29541_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net923),
    .D(_01869_),
    .Q_N(_12223_),
    .Q(\atari2600.ram[38][0] ));
 sg13g2_dfrbp_1 _29542_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net922),
    .D(_01870_),
    .Q_N(_12222_),
    .Q(\atari2600.ram[38][1] ));
 sg13g2_dfrbp_1 _29543_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net921),
    .D(_01871_),
    .Q_N(_12221_),
    .Q(\atari2600.ram[38][2] ));
 sg13g2_dfrbp_1 _29544_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net920),
    .D(_01872_),
    .Q_N(_12220_),
    .Q(\atari2600.ram[38][3] ));
 sg13g2_dfrbp_1 _29545_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net919),
    .D(_01873_),
    .Q_N(_12219_),
    .Q(\atari2600.ram[38][4] ));
 sg13g2_dfrbp_1 _29546_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net918),
    .D(_01874_),
    .Q_N(_12218_),
    .Q(\atari2600.ram[38][5] ));
 sg13g2_dfrbp_1 _29547_ (.CLK(clknet_leaf_364_clk),
    .RESET_B(net917),
    .D(_01875_),
    .Q_N(_12217_),
    .Q(\atari2600.ram[38][6] ));
 sg13g2_dfrbp_1 _29548_ (.CLK(clknet_leaf_363_clk),
    .RESET_B(net916),
    .D(_01876_),
    .Q_N(_12216_),
    .Q(\atari2600.ram[38][7] ));
 sg13g2_dfrbp_1 _29549_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net915),
    .D(net7126),
    .Q_N(_12215_),
    .Q(\atari2600.cpu.ABH[5] ));
 sg13g2_dfrbp_1 _29550_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net914),
    .D(net4387),
    .Q_N(_12214_),
    .Q(\atari2600.cpu.ABH[6] ));
 sg13g2_dfrbp_1 _29551_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net913),
    .D(net4453),
    .Q_N(_12213_),
    .Q(\atari2600.cpu.ABH[7] ));
 sg13g2_dfrbp_1 _29552_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net912),
    .D(_01880_),
    .Q_N(_12212_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _29553_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net911),
    .D(_01881_),
    .Q_N(_12211_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _29554_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net910),
    .D(_01882_),
    .Q_N(_00057_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _29555_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net909),
    .D(_01883_),
    .Q_N(_12210_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _29556_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net908),
    .D(_01884_),
    .Q_N(_00058_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _29557_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net907),
    .D(_01885_),
    .Q_N(_12209_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _29558_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net906),
    .D(_01886_),
    .Q_N(_00059_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _29559_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net905),
    .D(net7255),
    .Q_N(_00135_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _29560_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net904),
    .D(_01888_),
    .Q_N(_12208_),
    .Q(\atari2600.ram[9][0] ));
 sg13g2_dfrbp_1 _29561_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net903),
    .D(_01889_),
    .Q_N(_12207_),
    .Q(\atari2600.ram[9][1] ));
 sg13g2_dfrbp_1 _29562_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net902),
    .D(_01890_),
    .Q_N(_12206_),
    .Q(\atari2600.ram[9][2] ));
 sg13g2_dfrbp_1 _29563_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net901),
    .D(_01891_),
    .Q_N(_12205_),
    .Q(\atari2600.ram[9][3] ));
 sg13g2_dfrbp_1 _29564_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net900),
    .D(_01892_),
    .Q_N(_12204_),
    .Q(\atari2600.ram[9][4] ));
 sg13g2_dfrbp_1 _29565_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net899),
    .D(_01893_),
    .Q_N(_12203_),
    .Q(\atari2600.ram[9][5] ));
 sg13g2_dfrbp_1 _29566_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net898),
    .D(_01894_),
    .Q_N(_12202_),
    .Q(\atari2600.ram[9][6] ));
 sg13g2_dfrbp_1 _29567_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net897),
    .D(_01895_),
    .Q_N(_12201_),
    .Q(\atari2600.ram[9][7] ));
 sg13g2_dfrbp_1 _29568_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net896),
    .D(_01896_),
    .Q_N(_12200_),
    .Q(\scanline[19][0] ));
 sg13g2_dfrbp_1 _29569_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net895),
    .D(_01897_),
    .Q_N(_12199_),
    .Q(\scanline[19][1] ));
 sg13g2_dfrbp_1 _29570_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net894),
    .D(_01898_),
    .Q_N(_12198_),
    .Q(\scanline[19][2] ));
 sg13g2_dfrbp_1 _29571_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net893),
    .D(_01899_),
    .Q_N(_12197_),
    .Q(\scanline[19][3] ));
 sg13g2_dfrbp_1 _29572_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net892),
    .D(_01900_),
    .Q_N(_12196_),
    .Q(\scanline[19][4] ));
 sg13g2_dfrbp_1 _29573_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net891),
    .D(_01901_),
    .Q_N(_12195_),
    .Q(\scanline[19][5] ));
 sg13g2_dfrbp_1 _29574_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net890),
    .D(_01902_),
    .Q_N(_12194_),
    .Q(\scanline[19][6] ));
 sg13g2_dfrbp_1 _29575_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net889),
    .D(_01903_),
    .Q_N(_12193_),
    .Q(\scanline[29][0] ));
 sg13g2_dfrbp_1 _29576_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net888),
    .D(_01904_),
    .Q_N(_12192_),
    .Q(\scanline[29][1] ));
 sg13g2_dfrbp_1 _29577_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net887),
    .D(_01905_),
    .Q_N(_12191_),
    .Q(\scanline[29][2] ));
 sg13g2_dfrbp_1 _29578_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net886),
    .D(_01906_),
    .Q_N(_12190_),
    .Q(\scanline[29][3] ));
 sg13g2_dfrbp_1 _29579_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net885),
    .D(_01907_),
    .Q_N(_12189_),
    .Q(\scanline[29][4] ));
 sg13g2_dfrbp_1 _29580_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net884),
    .D(_01908_),
    .Q_N(_12188_),
    .Q(\scanline[29][5] ));
 sg13g2_dfrbp_1 _29581_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net883),
    .D(_01909_),
    .Q_N(_12187_),
    .Q(\scanline[29][6] ));
 sg13g2_dfrbp_1 _29582_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net882),
    .D(_01910_),
    .Q_N(_12186_),
    .Q(\scanline[39][0] ));
 sg13g2_dfrbp_1 _29583_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net881),
    .D(_01911_),
    .Q_N(_12185_),
    .Q(\scanline[39][1] ));
 sg13g2_dfrbp_1 _29584_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net880),
    .D(_01912_),
    .Q_N(_12184_),
    .Q(\scanline[39][2] ));
 sg13g2_dfrbp_1 _29585_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net879),
    .D(_01913_),
    .Q_N(_12183_),
    .Q(\scanline[39][3] ));
 sg13g2_dfrbp_1 _29586_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net878),
    .D(_01914_),
    .Q_N(_12182_),
    .Q(\scanline[39][4] ));
 sg13g2_dfrbp_1 _29587_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net877),
    .D(_01915_),
    .Q_N(_12181_),
    .Q(\scanline[39][5] ));
 sg13g2_dfrbp_1 _29588_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net876),
    .D(_01916_),
    .Q_N(_12180_),
    .Q(\scanline[39][6] ));
 sg13g2_dfrbp_1 _29589_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net875),
    .D(_01917_),
    .Q_N(_12179_),
    .Q(\scanline[49][0] ));
 sg13g2_dfrbp_1 _29590_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net874),
    .D(_01918_),
    .Q_N(_12178_),
    .Q(\scanline[49][1] ));
 sg13g2_dfrbp_1 _29591_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net873),
    .D(_01919_),
    .Q_N(_12177_),
    .Q(\scanline[49][2] ));
 sg13g2_dfrbp_1 _29592_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net872),
    .D(_01920_),
    .Q_N(_12176_),
    .Q(\scanline[49][3] ));
 sg13g2_dfrbp_1 _29593_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net871),
    .D(_01921_),
    .Q_N(_12175_),
    .Q(\scanline[49][4] ));
 sg13g2_dfrbp_1 _29594_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net870),
    .D(_01922_),
    .Q_N(_12174_),
    .Q(\scanline[49][5] ));
 sg13g2_dfrbp_1 _29595_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net869),
    .D(_01923_),
    .Q_N(_12173_),
    .Q(\scanline[49][6] ));
 sg13g2_dfrbp_1 _29596_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net868),
    .D(_01924_),
    .Q_N(_12172_),
    .Q(\scanline[59][0] ));
 sg13g2_dfrbp_1 _29597_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net867),
    .D(_01925_),
    .Q_N(_12171_),
    .Q(\scanline[59][1] ));
 sg13g2_dfrbp_1 _29598_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net866),
    .D(_01926_),
    .Q_N(_12170_),
    .Q(\scanline[59][2] ));
 sg13g2_dfrbp_1 _29599_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net865),
    .D(_01927_),
    .Q_N(_12169_),
    .Q(\scanline[59][3] ));
 sg13g2_dfrbp_1 _29600_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net864),
    .D(_01928_),
    .Q_N(_12168_),
    .Q(\scanline[59][4] ));
 sg13g2_dfrbp_1 _29601_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net863),
    .D(_01929_),
    .Q_N(_12167_),
    .Q(\scanline[59][5] ));
 sg13g2_dfrbp_1 _29602_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net862),
    .D(_01930_),
    .Q_N(_12166_),
    .Q(\scanline[59][6] ));
 sg13g2_dfrbp_1 _29603_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net861),
    .D(_01931_),
    .Q_N(_12165_),
    .Q(\scanline[69][0] ));
 sg13g2_dfrbp_1 _29604_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net860),
    .D(_01932_),
    .Q_N(_12164_),
    .Q(\scanline[69][1] ));
 sg13g2_dfrbp_1 _29605_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net859),
    .D(_01933_),
    .Q_N(_12163_),
    .Q(\scanline[69][2] ));
 sg13g2_dfrbp_1 _29606_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net858),
    .D(_01934_),
    .Q_N(_12162_),
    .Q(\scanline[69][3] ));
 sg13g2_dfrbp_1 _29607_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net857),
    .D(_01935_),
    .Q_N(_12161_),
    .Q(\scanline[69][4] ));
 sg13g2_dfrbp_1 _29608_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net856),
    .D(_01936_),
    .Q_N(_12160_),
    .Q(\scanline[69][5] ));
 sg13g2_dfrbp_1 _29609_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net855),
    .D(_01937_),
    .Q_N(_12159_),
    .Q(\scanline[69][6] ));
 sg13g2_dfrbp_1 _29610_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net854),
    .D(_01938_),
    .Q_N(_12158_),
    .Q(\scanline[79][0] ));
 sg13g2_dfrbp_1 _29611_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net853),
    .D(_01939_),
    .Q_N(_12157_),
    .Q(\scanline[79][1] ));
 sg13g2_dfrbp_1 _29612_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net852),
    .D(_01940_),
    .Q_N(_12156_),
    .Q(\scanline[79][2] ));
 sg13g2_dfrbp_1 _29613_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net851),
    .D(_01941_),
    .Q_N(_12155_),
    .Q(\scanline[79][3] ));
 sg13g2_dfrbp_1 _29614_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net850),
    .D(_01942_),
    .Q_N(_12154_),
    .Q(\scanline[79][4] ));
 sg13g2_dfrbp_1 _29615_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net849),
    .D(_01943_),
    .Q_N(_12153_),
    .Q(\scanline[79][5] ));
 sg13g2_dfrbp_1 _29616_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net848),
    .D(_01944_),
    .Q_N(_12152_),
    .Q(\scanline[79][6] ));
 sg13g2_dfrbp_1 _29617_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net847),
    .D(_01945_),
    .Q_N(_12151_),
    .Q(\scanline[89][0] ));
 sg13g2_dfrbp_1 _29618_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net846),
    .D(_01946_),
    .Q_N(_12150_),
    .Q(\scanline[89][1] ));
 sg13g2_dfrbp_1 _29619_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net845),
    .D(_01947_),
    .Q_N(_12149_),
    .Q(\scanline[89][2] ));
 sg13g2_dfrbp_1 _29620_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net844),
    .D(_01948_),
    .Q_N(_12148_),
    .Q(\scanline[89][3] ));
 sg13g2_dfrbp_1 _29621_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net843),
    .D(_01949_),
    .Q_N(_12147_),
    .Q(\scanline[89][4] ));
 sg13g2_dfrbp_1 _29622_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net842),
    .D(_01950_),
    .Q_N(_12146_),
    .Q(\scanline[89][5] ));
 sg13g2_dfrbp_1 _29623_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net841),
    .D(_01951_),
    .Q_N(_12145_),
    .Q(\scanline[89][6] ));
 sg13g2_dfrbp_1 _29624_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net840),
    .D(_01952_),
    .Q_N(_12144_),
    .Q(\scanline[99][0] ));
 sg13g2_dfrbp_1 _29625_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net839),
    .D(_01953_),
    .Q_N(_12143_),
    .Q(\scanline[99][1] ));
 sg13g2_dfrbp_1 _29626_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net838),
    .D(_01954_),
    .Q_N(_12142_),
    .Q(\scanline[99][2] ));
 sg13g2_dfrbp_1 _29627_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net837),
    .D(_01955_),
    .Q_N(_12141_),
    .Q(\scanline[99][3] ));
 sg13g2_dfrbp_1 _29628_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net836),
    .D(_01956_),
    .Q_N(_12140_),
    .Q(\scanline[99][4] ));
 sg13g2_dfrbp_1 _29629_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net835),
    .D(_01957_),
    .Q_N(_12139_),
    .Q(\scanline[99][5] ));
 sg13g2_dfrbp_1 _29630_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net834),
    .D(_01958_),
    .Q_N(_12138_),
    .Q(\scanline[99][6] ));
 sg13g2_dfrbp_1 _29631_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net833),
    .D(_01959_),
    .Q_N(_12137_),
    .Q(\scanline[109][0] ));
 sg13g2_dfrbp_1 _29632_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net832),
    .D(_01960_),
    .Q_N(_12136_),
    .Q(\scanline[109][1] ));
 sg13g2_dfrbp_1 _29633_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net831),
    .D(_01961_),
    .Q_N(_12135_),
    .Q(\scanline[109][2] ));
 sg13g2_dfrbp_1 _29634_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net830),
    .D(_01962_),
    .Q_N(_12134_),
    .Q(\scanline[109][3] ));
 sg13g2_dfrbp_1 _29635_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net829),
    .D(_01963_),
    .Q_N(_12133_),
    .Q(\scanline[109][4] ));
 sg13g2_dfrbp_1 _29636_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net828),
    .D(_01964_),
    .Q_N(_12132_),
    .Q(\scanline[109][5] ));
 sg13g2_dfrbp_1 _29637_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net827),
    .D(_01965_),
    .Q_N(_12131_),
    .Q(\scanline[109][6] ));
 sg13g2_dfrbp_1 _29638_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net826),
    .D(_01966_),
    .Q_N(_12130_),
    .Q(\scanline[119][0] ));
 sg13g2_dfrbp_1 _29639_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net825),
    .D(_01967_),
    .Q_N(_12129_),
    .Q(\scanline[119][1] ));
 sg13g2_dfrbp_1 _29640_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net824),
    .D(_01968_),
    .Q_N(_12128_),
    .Q(\scanline[119][2] ));
 sg13g2_dfrbp_1 _29641_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net823),
    .D(_01969_),
    .Q_N(_12127_),
    .Q(\scanline[119][3] ));
 sg13g2_dfrbp_1 _29642_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net822),
    .D(_01970_),
    .Q_N(_12126_),
    .Q(\scanline[119][4] ));
 sg13g2_dfrbp_1 _29643_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net804),
    .D(_01971_),
    .Q_N(_12125_),
    .Q(\scanline[119][5] ));
 sg13g2_dfrbp_1 _29644_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net803),
    .D(_01972_),
    .Q_N(_12124_),
    .Q(\scanline[119][6] ));
 sg13g2_dfrbp_1 _29645_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net802),
    .D(_01973_),
    .Q_N(_12123_),
    .Q(\scanline[129][0] ));
 sg13g2_dfrbp_1 _29646_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net801),
    .D(_01974_),
    .Q_N(_12122_),
    .Q(\scanline[129][1] ));
 sg13g2_dfrbp_1 _29647_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net800),
    .D(_01975_),
    .Q_N(_12121_),
    .Q(\scanline[129][2] ));
 sg13g2_dfrbp_1 _29648_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net799),
    .D(_01976_),
    .Q_N(_12120_),
    .Q(\scanline[129][3] ));
 sg13g2_dfrbp_1 _29649_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net798),
    .D(_01977_),
    .Q_N(_12119_),
    .Q(\scanline[129][4] ));
 sg13g2_dfrbp_1 _29650_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net797),
    .D(_01978_),
    .Q_N(_12118_),
    .Q(\scanline[129][5] ));
 sg13g2_dfrbp_1 _29651_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net796),
    .D(_01979_),
    .Q_N(_12117_),
    .Q(\scanline[129][6] ));
 sg13g2_dfrbp_1 _29652_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net795),
    .D(_01980_),
    .Q_N(_12116_),
    .Q(\scanline[139][0] ));
 sg13g2_dfrbp_1 _29653_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net794),
    .D(_01981_),
    .Q_N(_12115_),
    .Q(\scanline[139][1] ));
 sg13g2_dfrbp_1 _29654_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net793),
    .D(_01982_),
    .Q_N(_12114_),
    .Q(\scanline[139][2] ));
 sg13g2_dfrbp_1 _29655_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net792),
    .D(_01983_),
    .Q_N(_12113_),
    .Q(\scanline[139][3] ));
 sg13g2_dfrbp_1 _29656_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net791),
    .D(_01984_),
    .Q_N(_12112_),
    .Q(\scanline[139][4] ));
 sg13g2_dfrbp_1 _29657_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net790),
    .D(_01985_),
    .Q_N(_12111_),
    .Q(\scanline[139][5] ));
 sg13g2_dfrbp_1 _29658_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net789),
    .D(_01986_),
    .Q_N(_12110_),
    .Q(\scanline[139][6] ));
 sg13g2_dfrbp_1 _29659_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net788),
    .D(_01987_),
    .Q_N(_12109_),
    .Q(\scanline[149][0] ));
 sg13g2_dfrbp_1 _29660_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net787),
    .D(_01988_),
    .Q_N(_12108_),
    .Q(\scanline[149][1] ));
 sg13g2_dfrbp_1 _29661_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net786),
    .D(_01989_),
    .Q_N(_12107_),
    .Q(\scanline[149][2] ));
 sg13g2_dfrbp_1 _29662_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net785),
    .D(_01990_),
    .Q_N(_12106_),
    .Q(\scanline[149][3] ));
 sg13g2_dfrbp_1 _29663_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net784),
    .D(_01991_),
    .Q_N(_12105_),
    .Q(\scanline[149][4] ));
 sg13g2_dfrbp_1 _29664_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net783),
    .D(_01992_),
    .Q_N(_12104_),
    .Q(\scanline[149][5] ));
 sg13g2_dfrbp_1 _29665_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net782),
    .D(_01993_),
    .Q_N(_12103_),
    .Q(\scanline[149][6] ));
 sg13g2_dfrbp_1 _29666_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net781),
    .D(_01994_),
    .Q_N(_12102_),
    .Q(\scanline[159][0] ));
 sg13g2_dfrbp_1 _29667_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net780),
    .D(_01995_),
    .Q_N(_12101_),
    .Q(\scanline[159][1] ));
 sg13g2_dfrbp_1 _29668_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net779),
    .D(_01996_),
    .Q_N(_12100_),
    .Q(\scanline[159][2] ));
 sg13g2_dfrbp_1 _29669_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net778),
    .D(_01997_),
    .Q_N(_12099_),
    .Q(\scanline[159][3] ));
 sg13g2_dfrbp_1 _29670_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net777),
    .D(_01998_),
    .Q_N(_12098_),
    .Q(\scanline[159][4] ));
 sg13g2_dfrbp_1 _29671_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net776),
    .D(_01999_),
    .Q_N(_12097_),
    .Q(\scanline[159][5] ));
 sg13g2_dfrbp_1 _29672_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net775),
    .D(_02000_),
    .Q_N(_12096_),
    .Q(\scanline[159][6] ));
 sg13g2_dfrbp_1 _29673_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net774),
    .D(_02001_),
    .Q_N(_12095_),
    .Q(\scanline[25][0] ));
 sg13g2_dfrbp_1 _29674_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net773),
    .D(_02002_),
    .Q_N(_12094_),
    .Q(\scanline[25][1] ));
 sg13g2_dfrbp_1 _29675_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net772),
    .D(_02003_),
    .Q_N(_12093_),
    .Q(\scanline[25][2] ));
 sg13g2_dfrbp_1 _29676_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net771),
    .D(_02004_),
    .Q_N(_12092_),
    .Q(\scanline[25][3] ));
 sg13g2_dfrbp_1 _29677_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net770),
    .D(_02005_),
    .Q_N(_12091_),
    .Q(\scanline[25][4] ));
 sg13g2_dfrbp_1 _29678_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net769),
    .D(_02006_),
    .Q_N(_12090_),
    .Q(\scanline[25][5] ));
 sg13g2_dfrbp_1 _29679_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net768),
    .D(_02007_),
    .Q_N(_12089_),
    .Q(\scanline[25][6] ));
 sg13g2_dfrbp_1 _29680_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net767),
    .D(_02008_),
    .Q_N(_12088_),
    .Q(\scanline[26][0] ));
 sg13g2_dfrbp_1 _29681_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net766),
    .D(_02009_),
    .Q_N(_12087_),
    .Q(\scanline[26][1] ));
 sg13g2_dfrbp_1 _29682_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net765),
    .D(_02010_),
    .Q_N(_12086_),
    .Q(\scanline[26][2] ));
 sg13g2_dfrbp_1 _29683_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net764),
    .D(_02011_),
    .Q_N(_12085_),
    .Q(\scanline[26][3] ));
 sg13g2_dfrbp_1 _29684_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net763),
    .D(_02012_),
    .Q_N(_12084_),
    .Q(\scanline[26][4] ));
 sg13g2_dfrbp_1 _29685_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net762),
    .D(_02013_),
    .Q_N(_12083_),
    .Q(\scanline[26][5] ));
 sg13g2_dfrbp_1 _29686_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net761),
    .D(_02014_),
    .Q_N(_12082_),
    .Q(\scanline[26][6] ));
 sg13g2_dfrbp_1 _29687_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net760),
    .D(_02015_),
    .Q_N(_12081_),
    .Q(\scanline[27][0] ));
 sg13g2_dfrbp_1 _29688_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net759),
    .D(_02016_),
    .Q_N(_12080_),
    .Q(\scanline[27][1] ));
 sg13g2_dfrbp_1 _29689_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net758),
    .D(_02017_),
    .Q_N(_12079_),
    .Q(\scanline[27][2] ));
 sg13g2_dfrbp_1 _29690_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net757),
    .D(_02018_),
    .Q_N(_12078_),
    .Q(\scanline[27][3] ));
 sg13g2_dfrbp_1 _29691_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net756),
    .D(_02019_),
    .Q_N(_12077_),
    .Q(\scanline[27][4] ));
 sg13g2_dfrbp_1 _29692_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net755),
    .D(_02020_),
    .Q_N(_12076_),
    .Q(\scanline[27][5] ));
 sg13g2_dfrbp_1 _29693_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net754),
    .D(_02021_),
    .Q_N(_12075_),
    .Q(\scanline[27][6] ));
 sg13g2_dfrbp_1 _29694_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net753),
    .D(_02022_),
    .Q_N(_12074_),
    .Q(\scanline[28][0] ));
 sg13g2_dfrbp_1 _29695_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net752),
    .D(_02023_),
    .Q_N(_12073_),
    .Q(\scanline[28][1] ));
 sg13g2_dfrbp_1 _29696_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net751),
    .D(_02024_),
    .Q_N(_12072_),
    .Q(\scanline[28][2] ));
 sg13g2_dfrbp_1 _29697_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net750),
    .D(_02025_),
    .Q_N(_12071_),
    .Q(\scanline[28][3] ));
 sg13g2_dfrbp_1 _29698_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net749),
    .D(_02026_),
    .Q_N(_12070_),
    .Q(\scanline[28][4] ));
 sg13g2_dfrbp_1 _29699_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net748),
    .D(_02027_),
    .Q_N(_12069_),
    .Q(\scanline[28][5] ));
 sg13g2_dfrbp_1 _29700_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net747),
    .D(_02028_),
    .Q_N(_12068_),
    .Q(\scanline[28][6] ));
 sg13g2_dfrbp_1 _29701_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net746),
    .D(_02029_),
    .Q_N(_12067_),
    .Q(\scanline[2][0] ));
 sg13g2_dfrbp_1 _29702_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net745),
    .D(_02030_),
    .Q_N(_12066_),
    .Q(\scanline[2][1] ));
 sg13g2_dfrbp_1 _29703_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net744),
    .D(_02031_),
    .Q_N(_12065_),
    .Q(\scanline[2][2] ));
 sg13g2_dfrbp_1 _29704_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net743),
    .D(_02032_),
    .Q_N(_12064_),
    .Q(\scanline[2][3] ));
 sg13g2_dfrbp_1 _29705_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net742),
    .D(_02033_),
    .Q_N(_12063_),
    .Q(\scanline[2][4] ));
 sg13g2_dfrbp_1 _29706_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net741),
    .D(_02034_),
    .Q_N(_12062_),
    .Q(\scanline[2][5] ));
 sg13g2_dfrbp_1 _29707_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net740),
    .D(_02035_),
    .Q_N(_12061_),
    .Q(\scanline[2][6] ));
 sg13g2_dfrbp_1 _29708_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net739),
    .D(_02036_),
    .Q_N(_12060_),
    .Q(\scanline[30][0] ));
 sg13g2_dfrbp_1 _29709_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net738),
    .D(_02037_),
    .Q_N(_12059_),
    .Q(\scanline[30][1] ));
 sg13g2_dfrbp_1 _29710_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net737),
    .D(_02038_),
    .Q_N(_12058_),
    .Q(\scanline[30][2] ));
 sg13g2_dfrbp_1 _29711_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net736),
    .D(_02039_),
    .Q_N(_12057_),
    .Q(\scanline[30][3] ));
 sg13g2_dfrbp_1 _29712_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net735),
    .D(_02040_),
    .Q_N(_12056_),
    .Q(\scanline[30][4] ));
 sg13g2_dfrbp_1 _29713_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net734),
    .D(_02041_),
    .Q_N(_12055_),
    .Q(\scanline[30][5] ));
 sg13g2_dfrbp_1 _29714_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net733),
    .D(_02042_),
    .Q_N(_12054_),
    .Q(\scanline[30][6] ));
 sg13g2_dfrbp_1 _29715_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net732),
    .D(_02043_),
    .Q_N(_12053_),
    .Q(\scanline[31][0] ));
 sg13g2_dfrbp_1 _29716_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net731),
    .D(_02044_),
    .Q_N(_12052_),
    .Q(\scanline[31][1] ));
 sg13g2_dfrbp_1 _29717_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net730),
    .D(_02045_),
    .Q_N(_12051_),
    .Q(\scanline[31][2] ));
 sg13g2_dfrbp_1 _29718_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net729),
    .D(_02046_),
    .Q_N(_12050_),
    .Q(\scanline[31][3] ));
 sg13g2_dfrbp_1 _29719_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net728),
    .D(_02047_),
    .Q_N(_12049_),
    .Q(\scanline[31][4] ));
 sg13g2_dfrbp_1 _29720_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net727),
    .D(_02048_),
    .Q_N(_12048_),
    .Q(\scanline[31][5] ));
 sg13g2_dfrbp_1 _29721_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net726),
    .D(_02049_),
    .Q_N(_12047_),
    .Q(\scanline[31][6] ));
 sg13g2_dfrbp_1 _29722_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net725),
    .D(_02050_),
    .Q_N(_12046_),
    .Q(\scanline[32][0] ));
 sg13g2_dfrbp_1 _29723_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net724),
    .D(_02051_),
    .Q_N(_12045_),
    .Q(\scanline[32][1] ));
 sg13g2_dfrbp_1 _29724_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net723),
    .D(_02052_),
    .Q_N(_12044_),
    .Q(\scanline[32][2] ));
 sg13g2_dfrbp_1 _29725_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net722),
    .D(_02053_),
    .Q_N(_12043_),
    .Q(\scanline[32][3] ));
 sg13g2_dfrbp_1 _29726_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net721),
    .D(_02054_),
    .Q_N(_12042_),
    .Q(\scanline[32][4] ));
 sg13g2_dfrbp_1 _29727_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net720),
    .D(_02055_),
    .Q_N(_12041_),
    .Q(\scanline[32][5] ));
 sg13g2_dfrbp_1 _29728_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net719),
    .D(_02056_),
    .Q_N(_12040_),
    .Q(\scanline[32][6] ));
 sg13g2_dfrbp_1 _29729_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net718),
    .D(_02057_),
    .Q_N(_12039_),
    .Q(\scanline[33][0] ));
 sg13g2_dfrbp_1 _29730_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net717),
    .D(_02058_),
    .Q_N(_12038_),
    .Q(\scanline[33][1] ));
 sg13g2_dfrbp_1 _29731_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net716),
    .D(_02059_),
    .Q_N(_12037_),
    .Q(\scanline[33][2] ));
 sg13g2_dfrbp_1 _29732_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net715),
    .D(_02060_),
    .Q_N(_12036_),
    .Q(\scanline[33][3] ));
 sg13g2_dfrbp_1 _29733_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net714),
    .D(_02061_),
    .Q_N(_12035_),
    .Q(\scanline[33][4] ));
 sg13g2_dfrbp_1 _29734_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net713),
    .D(_02062_),
    .Q_N(_12034_),
    .Q(\scanline[33][5] ));
 sg13g2_dfrbp_1 _29735_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net712),
    .D(_02063_),
    .Q_N(_12033_),
    .Q(\scanline[33][6] ));
 sg13g2_dfrbp_1 _29736_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net711),
    .D(_02064_),
    .Q_N(_12032_),
    .Q(\scanline[34][0] ));
 sg13g2_dfrbp_1 _29737_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net710),
    .D(_02065_),
    .Q_N(_12031_),
    .Q(\scanline[34][1] ));
 sg13g2_dfrbp_1 _29738_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net709),
    .D(_02066_),
    .Q_N(_12030_),
    .Q(\scanline[34][2] ));
 sg13g2_dfrbp_1 _29739_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net708),
    .D(_02067_),
    .Q_N(_12029_),
    .Q(\scanline[34][3] ));
 sg13g2_dfrbp_1 _29740_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net707),
    .D(_02068_),
    .Q_N(_12028_),
    .Q(\scanline[34][4] ));
 sg13g2_dfrbp_1 _29741_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net706),
    .D(_02069_),
    .Q_N(_12027_),
    .Q(\scanline[34][5] ));
 sg13g2_dfrbp_1 _29742_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net705),
    .D(_02070_),
    .Q_N(_12026_),
    .Q(\scanline[34][6] ));
 sg13g2_dfrbp_1 _29743_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net704),
    .D(_02071_),
    .Q_N(_12025_),
    .Q(\scanline[35][0] ));
 sg13g2_dfrbp_1 _29744_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net703),
    .D(_02072_),
    .Q_N(_12024_),
    .Q(\scanline[35][1] ));
 sg13g2_dfrbp_1 _29745_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net702),
    .D(_02073_),
    .Q_N(_12023_),
    .Q(\scanline[35][2] ));
 sg13g2_dfrbp_1 _29746_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net701),
    .D(_02074_),
    .Q_N(_12022_),
    .Q(\scanline[35][3] ));
 sg13g2_dfrbp_1 _29747_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net700),
    .D(_02075_),
    .Q_N(_12021_),
    .Q(\scanline[35][4] ));
 sg13g2_dfrbp_1 _29748_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net699),
    .D(_02076_),
    .Q_N(_12020_),
    .Q(\scanline[35][5] ));
 sg13g2_dfrbp_1 _29749_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net698),
    .D(_02077_),
    .Q_N(_12019_),
    .Q(\scanline[35][6] ));
 sg13g2_dfrbp_1 _29750_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net697),
    .D(_02078_),
    .Q_N(_12018_),
    .Q(\scanline[36][0] ));
 sg13g2_dfrbp_1 _29751_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net696),
    .D(_02079_),
    .Q_N(_12017_),
    .Q(\scanline[36][1] ));
 sg13g2_dfrbp_1 _29752_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net695),
    .D(_02080_),
    .Q_N(_12016_),
    .Q(\scanline[36][2] ));
 sg13g2_dfrbp_1 _29753_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net694),
    .D(_02081_),
    .Q_N(_12015_),
    .Q(\scanline[36][3] ));
 sg13g2_dfrbp_1 _29754_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net693),
    .D(_02082_),
    .Q_N(_12014_),
    .Q(\scanline[36][4] ));
 sg13g2_dfrbp_1 _29755_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net692),
    .D(_02083_),
    .Q_N(_12013_),
    .Q(\scanline[36][5] ));
 sg13g2_dfrbp_1 _29756_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net691),
    .D(_02084_),
    .Q_N(_12012_),
    .Q(\scanline[36][6] ));
 sg13g2_dfrbp_1 _29757_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net690),
    .D(_02085_),
    .Q_N(_12011_),
    .Q(\scanline[37][0] ));
 sg13g2_dfrbp_1 _29758_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net689),
    .D(_02086_),
    .Q_N(_12010_),
    .Q(\scanline[37][1] ));
 sg13g2_dfrbp_1 _29759_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net688),
    .D(_02087_),
    .Q_N(_12009_),
    .Q(\scanline[37][2] ));
 sg13g2_dfrbp_1 _29760_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net687),
    .D(_02088_),
    .Q_N(_12008_),
    .Q(\scanline[37][3] ));
 sg13g2_dfrbp_1 _29761_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net686),
    .D(_02089_),
    .Q_N(_12007_),
    .Q(\scanline[37][4] ));
 sg13g2_dfrbp_1 _29762_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net685),
    .D(_02090_),
    .Q_N(_12006_),
    .Q(\scanline[37][5] ));
 sg13g2_dfrbp_1 _29763_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net684),
    .D(_02091_),
    .Q_N(_12005_),
    .Q(\scanline[37][6] ));
 sg13g2_dfrbp_1 _29764_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net683),
    .D(_02092_),
    .Q_N(_12004_),
    .Q(\scanline[38][0] ));
 sg13g2_dfrbp_1 _29765_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net682),
    .D(_02093_),
    .Q_N(_12003_),
    .Q(\scanline[38][1] ));
 sg13g2_dfrbp_1 _29766_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net681),
    .D(_02094_),
    .Q_N(_12002_),
    .Q(\scanline[38][2] ));
 sg13g2_dfrbp_1 _29767_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net680),
    .D(_02095_),
    .Q_N(_12001_),
    .Q(\scanline[38][3] ));
 sg13g2_dfrbp_1 _29768_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net679),
    .D(_02096_),
    .Q_N(_12000_),
    .Q(\scanline[38][4] ));
 sg13g2_dfrbp_1 _29769_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net678),
    .D(_02097_),
    .Q_N(_11999_),
    .Q(\scanline[38][5] ));
 sg13g2_dfrbp_1 _29770_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net677),
    .D(_02098_),
    .Q_N(_11998_),
    .Q(\scanline[38][6] ));
 sg13g2_dfrbp_1 _29771_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net676),
    .D(_02099_),
    .Q_N(_11997_),
    .Q(\scanline[3][0] ));
 sg13g2_dfrbp_1 _29772_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net675),
    .D(_02100_),
    .Q_N(_11996_),
    .Q(\scanline[3][1] ));
 sg13g2_dfrbp_1 _29773_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net674),
    .D(_02101_),
    .Q_N(_11995_),
    .Q(\scanline[3][2] ));
 sg13g2_dfrbp_1 _29774_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net673),
    .D(_02102_),
    .Q_N(_11994_),
    .Q(\scanline[3][3] ));
 sg13g2_dfrbp_1 _29775_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net672),
    .D(_02103_),
    .Q_N(_11993_),
    .Q(\scanline[3][4] ));
 sg13g2_dfrbp_1 _29776_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net671),
    .D(_02104_),
    .Q_N(_11992_),
    .Q(\scanline[3][5] ));
 sg13g2_dfrbp_1 _29777_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net670),
    .D(_02105_),
    .Q_N(_11991_),
    .Q(\scanline[3][6] ));
 sg13g2_dfrbp_1 _29778_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net669),
    .D(_02106_),
    .Q_N(_11990_),
    .Q(\scanline[40][0] ));
 sg13g2_dfrbp_1 _29779_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net668),
    .D(_02107_),
    .Q_N(_11989_),
    .Q(\scanline[40][1] ));
 sg13g2_dfrbp_1 _29780_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net667),
    .D(_02108_),
    .Q_N(_11988_),
    .Q(\scanline[40][2] ));
 sg13g2_dfrbp_1 _29781_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net666),
    .D(_02109_),
    .Q_N(_11987_),
    .Q(\scanline[40][3] ));
 sg13g2_dfrbp_1 _29782_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net665),
    .D(_02110_),
    .Q_N(_11986_),
    .Q(\scanline[40][4] ));
 sg13g2_dfrbp_1 _29783_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net664),
    .D(_02111_),
    .Q_N(_11985_),
    .Q(\scanline[40][5] ));
 sg13g2_dfrbp_1 _29784_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net663),
    .D(_02112_),
    .Q_N(_11984_),
    .Q(\scanline[40][6] ));
 sg13g2_dfrbp_1 _29785_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net662),
    .D(_02113_),
    .Q_N(_11983_),
    .Q(\scanline[41][0] ));
 sg13g2_dfrbp_1 _29786_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net661),
    .D(_02114_),
    .Q_N(_11982_),
    .Q(\scanline[41][1] ));
 sg13g2_dfrbp_1 _29787_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net660),
    .D(_02115_),
    .Q_N(_11981_),
    .Q(\scanline[41][2] ));
 sg13g2_dfrbp_1 _29788_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net659),
    .D(_02116_),
    .Q_N(_11980_),
    .Q(\scanline[41][3] ));
 sg13g2_dfrbp_1 _29789_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net658),
    .D(_02117_),
    .Q_N(_11979_),
    .Q(\scanline[41][4] ));
 sg13g2_dfrbp_1 _29790_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net657),
    .D(_02118_),
    .Q_N(_11978_),
    .Q(\scanline[41][5] ));
 sg13g2_dfrbp_1 _29791_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net656),
    .D(_02119_),
    .Q_N(_11977_),
    .Q(\scanline[41][6] ));
 sg13g2_dfrbp_1 _29792_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net655),
    .D(_02120_),
    .Q_N(_11976_),
    .Q(\scanline[42][0] ));
 sg13g2_dfrbp_1 _29793_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net654),
    .D(_02121_),
    .Q_N(_11975_),
    .Q(\scanline[42][1] ));
 sg13g2_dfrbp_1 _29794_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net653),
    .D(_02122_),
    .Q_N(_11974_),
    .Q(\scanline[42][2] ));
 sg13g2_dfrbp_1 _29795_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net652),
    .D(_02123_),
    .Q_N(_11973_),
    .Q(\scanline[42][3] ));
 sg13g2_dfrbp_1 _29796_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net651),
    .D(_02124_),
    .Q_N(_11972_),
    .Q(\scanline[42][4] ));
 sg13g2_dfrbp_1 _29797_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net650),
    .D(_02125_),
    .Q_N(_11971_),
    .Q(\scanline[42][5] ));
 sg13g2_dfrbp_1 _29798_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net649),
    .D(_02126_),
    .Q_N(_11970_),
    .Q(\scanline[42][6] ));
 sg13g2_dfrbp_1 _29799_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net648),
    .D(_02127_),
    .Q_N(_11969_),
    .Q(\scanline[43][0] ));
 sg13g2_dfrbp_1 _29800_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net647),
    .D(_02128_),
    .Q_N(_11968_),
    .Q(\scanline[43][1] ));
 sg13g2_dfrbp_1 _29801_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net646),
    .D(_02129_),
    .Q_N(_11967_),
    .Q(\scanline[43][2] ));
 sg13g2_dfrbp_1 _29802_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net645),
    .D(_02130_),
    .Q_N(_11966_),
    .Q(\scanline[43][3] ));
 sg13g2_dfrbp_1 _29803_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net644),
    .D(_02131_),
    .Q_N(_11965_),
    .Q(\scanline[43][4] ));
 sg13g2_dfrbp_1 _29804_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net643),
    .D(_02132_),
    .Q_N(_11964_),
    .Q(\scanline[43][5] ));
 sg13g2_dfrbp_1 _29805_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net642),
    .D(_02133_),
    .Q_N(_11963_),
    .Q(\scanline[43][6] ));
 sg13g2_dfrbp_1 _29806_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net641),
    .D(_02134_),
    .Q_N(_11962_),
    .Q(\scanline[44][0] ));
 sg13g2_dfrbp_1 _29807_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net640),
    .D(_02135_),
    .Q_N(_11961_),
    .Q(\scanline[44][1] ));
 sg13g2_dfrbp_1 _29808_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net639),
    .D(_02136_),
    .Q_N(_11960_),
    .Q(\scanline[44][2] ));
 sg13g2_dfrbp_1 _29809_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net638),
    .D(_02137_),
    .Q_N(_11959_),
    .Q(\scanline[44][3] ));
 sg13g2_dfrbp_1 _29810_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net637),
    .D(_02138_),
    .Q_N(_11958_),
    .Q(\scanline[44][4] ));
 sg13g2_dfrbp_1 _29811_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net636),
    .D(_02139_),
    .Q_N(_11957_),
    .Q(\scanline[44][5] ));
 sg13g2_dfrbp_1 _29812_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net635),
    .D(_02140_),
    .Q_N(_11956_),
    .Q(\scanline[44][6] ));
 sg13g2_dfrbp_1 _29813_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net634),
    .D(_02141_),
    .Q_N(_11955_),
    .Q(\scanline[45][0] ));
 sg13g2_dfrbp_1 _29814_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net633),
    .D(_02142_),
    .Q_N(_11954_),
    .Q(\scanline[45][1] ));
 sg13g2_dfrbp_1 _29815_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net632),
    .D(_02143_),
    .Q_N(_11953_),
    .Q(\scanline[45][2] ));
 sg13g2_dfrbp_1 _29816_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net631),
    .D(_02144_),
    .Q_N(_11952_),
    .Q(\scanline[45][3] ));
 sg13g2_dfrbp_1 _29817_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net630),
    .D(_02145_),
    .Q_N(_11951_),
    .Q(\scanline[45][4] ));
 sg13g2_dfrbp_1 _29818_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net629),
    .D(_02146_),
    .Q_N(_11950_),
    .Q(\scanline[45][5] ));
 sg13g2_dfrbp_1 _29819_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net628),
    .D(_02147_),
    .Q_N(_11949_),
    .Q(\scanline[45][6] ));
 sg13g2_dfrbp_1 _29820_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net627),
    .D(_02148_),
    .Q_N(_11948_),
    .Q(\scanline[46][0] ));
 sg13g2_dfrbp_1 _29821_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net626),
    .D(_02149_),
    .Q_N(_11947_),
    .Q(\scanline[46][1] ));
 sg13g2_dfrbp_1 _29822_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net625),
    .D(_02150_),
    .Q_N(_11946_),
    .Q(\scanline[46][2] ));
 sg13g2_dfrbp_1 _29823_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net624),
    .D(_02151_),
    .Q_N(_11945_),
    .Q(\scanline[46][3] ));
 sg13g2_dfrbp_1 _29824_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net623),
    .D(_02152_),
    .Q_N(_11944_),
    .Q(\scanline[46][4] ));
 sg13g2_dfrbp_1 _29825_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net622),
    .D(_02153_),
    .Q_N(_11943_),
    .Q(\scanline[46][5] ));
 sg13g2_dfrbp_1 _29826_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net621),
    .D(_02154_),
    .Q_N(_11942_),
    .Q(\scanline[46][6] ));
 sg13g2_dfrbp_1 _29827_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net620),
    .D(_02155_),
    .Q_N(_11941_),
    .Q(\scanline[47][0] ));
 sg13g2_dfrbp_1 _29828_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net619),
    .D(_02156_),
    .Q_N(_11940_),
    .Q(\scanline[47][1] ));
 sg13g2_dfrbp_1 _29829_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net618),
    .D(_02157_),
    .Q_N(_11939_),
    .Q(\scanline[47][2] ));
 sg13g2_dfrbp_1 _29830_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net617),
    .D(_02158_),
    .Q_N(_11938_),
    .Q(\scanline[47][3] ));
 sg13g2_dfrbp_1 _29831_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net616),
    .D(_02159_),
    .Q_N(_11937_),
    .Q(\scanline[47][4] ));
 sg13g2_dfrbp_1 _29832_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net615),
    .D(_02160_),
    .Q_N(_11936_),
    .Q(\scanline[47][5] ));
 sg13g2_dfrbp_1 _29833_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net614),
    .D(_02161_),
    .Q_N(_11935_),
    .Q(\scanline[47][6] ));
 sg13g2_dfrbp_1 _29834_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net613),
    .D(_02162_),
    .Q_N(_11934_),
    .Q(\scanline[48][0] ));
 sg13g2_dfrbp_1 _29835_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net612),
    .D(_02163_),
    .Q_N(_11933_),
    .Q(\scanline[48][1] ));
 sg13g2_dfrbp_1 _29836_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net611),
    .D(_02164_),
    .Q_N(_11932_),
    .Q(\scanline[48][2] ));
 sg13g2_dfrbp_1 _29837_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net610),
    .D(_02165_),
    .Q_N(_11931_),
    .Q(\scanline[48][3] ));
 sg13g2_dfrbp_1 _29838_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net609),
    .D(_02166_),
    .Q_N(_11930_),
    .Q(\scanline[48][4] ));
 sg13g2_dfrbp_1 _29839_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net608),
    .D(_02167_),
    .Q_N(_11929_),
    .Q(\scanline[48][5] ));
 sg13g2_dfrbp_1 _29840_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net607),
    .D(_02168_),
    .Q_N(_11928_),
    .Q(\scanline[48][6] ));
 sg13g2_dfrbp_1 _29841_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net606),
    .D(_02169_),
    .Q_N(_11927_),
    .Q(\scanline[4][0] ));
 sg13g2_dfrbp_1 _29842_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net605),
    .D(_02170_),
    .Q_N(_11926_),
    .Q(\scanline[4][1] ));
 sg13g2_dfrbp_1 _29843_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net604),
    .D(_02171_),
    .Q_N(_11925_),
    .Q(\scanline[4][2] ));
 sg13g2_dfrbp_1 _29844_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net603),
    .D(_02172_),
    .Q_N(_11924_),
    .Q(\scanline[4][3] ));
 sg13g2_dfrbp_1 _29845_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net602),
    .D(_02173_),
    .Q_N(_11923_),
    .Q(\scanline[4][4] ));
 sg13g2_dfrbp_1 _29846_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net601),
    .D(_02174_),
    .Q_N(_11922_),
    .Q(\scanline[4][5] ));
 sg13g2_dfrbp_1 _29847_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net600),
    .D(_02175_),
    .Q_N(_11921_),
    .Q(\scanline[4][6] ));
 sg13g2_dfrbp_1 _29848_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net599),
    .D(_02176_),
    .Q_N(_11920_),
    .Q(\scanline[50][0] ));
 sg13g2_dfrbp_1 _29849_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net598),
    .D(_02177_),
    .Q_N(_11919_),
    .Q(\scanline[50][1] ));
 sg13g2_dfrbp_1 _29850_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net597),
    .D(_02178_),
    .Q_N(_11918_),
    .Q(\scanline[50][2] ));
 sg13g2_dfrbp_1 _29851_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net596),
    .D(_02179_),
    .Q_N(_11917_),
    .Q(\scanline[50][3] ));
 sg13g2_dfrbp_1 _29852_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net595),
    .D(_02180_),
    .Q_N(_11916_),
    .Q(\scanline[50][4] ));
 sg13g2_dfrbp_1 _29853_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net594),
    .D(_02181_),
    .Q_N(_11915_),
    .Q(\scanline[50][5] ));
 sg13g2_dfrbp_1 _29854_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net593),
    .D(_02182_),
    .Q_N(_11914_),
    .Q(\scanline[50][6] ));
 sg13g2_dfrbp_1 _29855_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net592),
    .D(_02183_),
    .Q_N(_11913_),
    .Q(\scanline[51][0] ));
 sg13g2_dfrbp_1 _29856_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net591),
    .D(_02184_),
    .Q_N(_11912_),
    .Q(\scanline[51][1] ));
 sg13g2_dfrbp_1 _29857_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net590),
    .D(_02185_),
    .Q_N(_11911_),
    .Q(\scanline[51][2] ));
 sg13g2_dfrbp_1 _29858_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net589),
    .D(_02186_),
    .Q_N(_11910_),
    .Q(\scanline[51][3] ));
 sg13g2_dfrbp_1 _29859_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net588),
    .D(_02187_),
    .Q_N(_11909_),
    .Q(\scanline[51][4] ));
 sg13g2_dfrbp_1 _29860_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net587),
    .D(_02188_),
    .Q_N(_11908_),
    .Q(\scanline[51][5] ));
 sg13g2_dfrbp_1 _29861_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net586),
    .D(_02189_),
    .Q_N(_11907_),
    .Q(\scanline[51][6] ));
 sg13g2_dfrbp_1 _29862_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net585),
    .D(_02190_),
    .Q_N(_11906_),
    .Q(\scanline[52][0] ));
 sg13g2_dfrbp_1 _29863_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net584),
    .D(_02191_),
    .Q_N(_11905_),
    .Q(\scanline[52][1] ));
 sg13g2_dfrbp_1 _29864_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net583),
    .D(_02192_),
    .Q_N(_11904_),
    .Q(\scanline[52][2] ));
 sg13g2_dfrbp_1 _29865_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net582),
    .D(_02193_),
    .Q_N(_11903_),
    .Q(\scanline[52][3] ));
 sg13g2_dfrbp_1 _29866_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net581),
    .D(_02194_),
    .Q_N(_11902_),
    .Q(\scanline[52][4] ));
 sg13g2_dfrbp_1 _29867_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net580),
    .D(_02195_),
    .Q_N(_11901_),
    .Q(\scanline[52][5] ));
 sg13g2_dfrbp_1 _29868_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net579),
    .D(_02196_),
    .Q_N(_11900_),
    .Q(\scanline[52][6] ));
 sg13g2_dfrbp_1 _29869_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net578),
    .D(_02197_),
    .Q_N(_11899_),
    .Q(\scanline[53][0] ));
 sg13g2_dfrbp_1 _29870_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net577),
    .D(_02198_),
    .Q_N(_11898_),
    .Q(\scanline[53][1] ));
 sg13g2_dfrbp_1 _29871_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net576),
    .D(_02199_),
    .Q_N(_11897_),
    .Q(\scanline[53][2] ));
 sg13g2_dfrbp_1 _29872_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net575),
    .D(_02200_),
    .Q_N(_11896_),
    .Q(\scanline[53][3] ));
 sg13g2_dfrbp_1 _29873_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net574),
    .D(_02201_),
    .Q_N(_11895_),
    .Q(\scanline[53][4] ));
 sg13g2_dfrbp_1 _29874_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net573),
    .D(_02202_),
    .Q_N(_11894_),
    .Q(\scanline[53][5] ));
 sg13g2_dfrbp_1 _29875_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net572),
    .D(_02203_),
    .Q_N(_11893_),
    .Q(\scanline[53][6] ));
 sg13g2_dfrbp_1 _29876_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net571),
    .D(_02204_),
    .Q_N(_11892_),
    .Q(\scanline[54][0] ));
 sg13g2_dfrbp_1 _29877_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net570),
    .D(_02205_),
    .Q_N(_11891_),
    .Q(\scanline[54][1] ));
 sg13g2_dfrbp_1 _29878_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net569),
    .D(_02206_),
    .Q_N(_11890_),
    .Q(\scanline[54][2] ));
 sg13g2_dfrbp_1 _29879_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net568),
    .D(_02207_),
    .Q_N(_11889_),
    .Q(\scanline[54][3] ));
 sg13g2_dfrbp_1 _29880_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net567),
    .D(_02208_),
    .Q_N(_11888_),
    .Q(\scanline[54][4] ));
 sg13g2_dfrbp_1 _29881_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net566),
    .D(_02209_),
    .Q_N(_11887_),
    .Q(\scanline[54][5] ));
 sg13g2_dfrbp_1 _29882_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net565),
    .D(_02210_),
    .Q_N(_11886_),
    .Q(\scanline[54][6] ));
 sg13g2_dfrbp_1 _29883_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net564),
    .D(_02211_),
    .Q_N(_11885_),
    .Q(\scanline[55][0] ));
 sg13g2_dfrbp_1 _29884_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net563),
    .D(_02212_),
    .Q_N(_11884_),
    .Q(\scanline[55][1] ));
 sg13g2_dfrbp_1 _29885_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net562),
    .D(_02213_),
    .Q_N(_11883_),
    .Q(\scanline[55][2] ));
 sg13g2_dfrbp_1 _29886_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net561),
    .D(_02214_),
    .Q_N(_11882_),
    .Q(\scanline[55][3] ));
 sg13g2_dfrbp_1 _29887_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net560),
    .D(_02215_),
    .Q_N(_11881_),
    .Q(\scanline[55][4] ));
 sg13g2_dfrbp_1 _29888_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net559),
    .D(_02216_),
    .Q_N(_11880_),
    .Q(\scanline[55][5] ));
 sg13g2_dfrbp_1 _29889_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net558),
    .D(_02217_),
    .Q_N(_11879_),
    .Q(\scanline[55][6] ));
 sg13g2_dfrbp_1 _29890_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net557),
    .D(_02218_),
    .Q_N(_11878_),
    .Q(\scanline[56][0] ));
 sg13g2_dfrbp_1 _29891_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net556),
    .D(_02219_),
    .Q_N(_11877_),
    .Q(\scanline[56][1] ));
 sg13g2_dfrbp_1 _29892_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net555),
    .D(_02220_),
    .Q_N(_11876_),
    .Q(\scanline[56][2] ));
 sg13g2_dfrbp_1 _29893_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net554),
    .D(_02221_),
    .Q_N(_11875_),
    .Q(\scanline[56][3] ));
 sg13g2_dfrbp_1 _29894_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net553),
    .D(_02222_),
    .Q_N(_11874_),
    .Q(\scanline[56][4] ));
 sg13g2_dfrbp_1 _29895_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net552),
    .D(_02223_),
    .Q_N(_11873_),
    .Q(\scanline[56][5] ));
 sg13g2_dfrbp_1 _29896_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net551),
    .D(_02224_),
    .Q_N(_11872_),
    .Q(\scanline[56][6] ));
 sg13g2_dfrbp_1 _29897_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net550),
    .D(_02225_),
    .Q_N(_11871_),
    .Q(\scanline[57][0] ));
 sg13g2_dfrbp_1 _29898_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net549),
    .D(_02226_),
    .Q_N(_11870_),
    .Q(\scanline[57][1] ));
 sg13g2_dfrbp_1 _29899_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net548),
    .D(_02227_),
    .Q_N(_11869_),
    .Q(\scanline[57][2] ));
 sg13g2_dfrbp_1 _29900_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net547),
    .D(_02228_),
    .Q_N(_11868_),
    .Q(\scanline[57][3] ));
 sg13g2_dfrbp_1 _29901_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net546),
    .D(_02229_),
    .Q_N(_11867_),
    .Q(\scanline[57][4] ));
 sg13g2_dfrbp_1 _29902_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net545),
    .D(_02230_),
    .Q_N(_11866_),
    .Q(\scanline[57][5] ));
 sg13g2_dfrbp_1 _29903_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net544),
    .D(_02231_),
    .Q_N(_11865_),
    .Q(\scanline[57][6] ));
 sg13g2_dfrbp_1 _29904_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net543),
    .D(_02232_),
    .Q_N(_11864_),
    .Q(\scanline[58][0] ));
 sg13g2_dfrbp_1 _29905_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net542),
    .D(_02233_),
    .Q_N(_11863_),
    .Q(\scanline[58][1] ));
 sg13g2_dfrbp_1 _29906_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net541),
    .D(_02234_),
    .Q_N(_11862_),
    .Q(\scanline[58][2] ));
 sg13g2_dfrbp_1 _29907_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net540),
    .D(_02235_),
    .Q_N(_11861_),
    .Q(\scanline[58][3] ));
 sg13g2_dfrbp_1 _29908_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net539),
    .D(_02236_),
    .Q_N(_11860_),
    .Q(\scanline[58][4] ));
 sg13g2_dfrbp_1 _29909_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net538),
    .D(_02237_),
    .Q_N(_11859_),
    .Q(\scanline[58][5] ));
 sg13g2_dfrbp_1 _29910_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net537),
    .D(_02238_),
    .Q_N(_11858_),
    .Q(\scanline[58][6] ));
 sg13g2_dfrbp_1 _29911_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net536),
    .D(_02239_),
    .Q_N(_11857_),
    .Q(\scanline[5][0] ));
 sg13g2_dfrbp_1 _29912_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net535),
    .D(_02240_),
    .Q_N(_11856_),
    .Q(\scanline[5][1] ));
 sg13g2_dfrbp_1 _29913_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net534),
    .D(_02241_),
    .Q_N(_11855_),
    .Q(\scanline[5][2] ));
 sg13g2_dfrbp_1 _29914_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net533),
    .D(_02242_),
    .Q_N(_11854_),
    .Q(\scanline[5][3] ));
 sg13g2_dfrbp_1 _29915_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net532),
    .D(_02243_),
    .Q_N(_11853_),
    .Q(\scanline[5][4] ));
 sg13g2_dfrbp_1 _29916_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net531),
    .D(_02244_),
    .Q_N(_11852_),
    .Q(\scanline[5][5] ));
 sg13g2_dfrbp_1 _29917_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net530),
    .D(_02245_),
    .Q_N(_11851_),
    .Q(\scanline[5][6] ));
 sg13g2_dfrbp_1 _29918_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net529),
    .D(_02246_),
    .Q_N(_11850_),
    .Q(\scanline[60][0] ));
 sg13g2_dfrbp_1 _29919_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net528),
    .D(_02247_),
    .Q_N(_11849_),
    .Q(\scanline[60][1] ));
 sg13g2_dfrbp_1 _29920_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net527),
    .D(_02248_),
    .Q_N(_11848_),
    .Q(\scanline[60][2] ));
 sg13g2_dfrbp_1 _29921_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net526),
    .D(_02249_),
    .Q_N(_11847_),
    .Q(\scanline[60][3] ));
 sg13g2_dfrbp_1 _29922_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net525),
    .D(_02250_),
    .Q_N(_11846_),
    .Q(\scanline[60][4] ));
 sg13g2_dfrbp_1 _29923_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net524),
    .D(_02251_),
    .Q_N(_11845_),
    .Q(\scanline[60][5] ));
 sg13g2_dfrbp_1 _29924_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net523),
    .D(_02252_),
    .Q_N(_11844_),
    .Q(\scanline[60][6] ));
 sg13g2_dfrbp_1 _29925_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net522),
    .D(_02253_),
    .Q_N(_11843_),
    .Q(\scanline[61][0] ));
 sg13g2_dfrbp_1 _29926_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net521),
    .D(_02254_),
    .Q_N(_11842_),
    .Q(\scanline[61][1] ));
 sg13g2_dfrbp_1 _29927_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net520),
    .D(_02255_),
    .Q_N(_11841_),
    .Q(\scanline[61][2] ));
 sg13g2_dfrbp_1 _29928_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net519),
    .D(_02256_),
    .Q_N(_11840_),
    .Q(\scanline[61][3] ));
 sg13g2_dfrbp_1 _29929_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net518),
    .D(_02257_),
    .Q_N(_11839_),
    .Q(\scanline[61][4] ));
 sg13g2_dfrbp_1 _29930_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net517),
    .D(_02258_),
    .Q_N(_11838_),
    .Q(\scanline[61][5] ));
 sg13g2_dfrbp_1 _29931_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net516),
    .D(_02259_),
    .Q_N(_11837_),
    .Q(\scanline[61][6] ));
 sg13g2_dfrbp_1 _29932_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net515),
    .D(_02260_),
    .Q_N(_11836_),
    .Q(\scanline[62][0] ));
 sg13g2_dfrbp_1 _29933_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net514),
    .D(_02261_),
    .Q_N(_11835_),
    .Q(\scanline[62][1] ));
 sg13g2_dfrbp_1 _29934_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net513),
    .D(_02262_),
    .Q_N(_11834_),
    .Q(\scanline[62][2] ));
 sg13g2_dfrbp_1 _29935_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net512),
    .D(_02263_),
    .Q_N(_11833_),
    .Q(\scanline[62][3] ));
 sg13g2_dfrbp_1 _29936_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net511),
    .D(_02264_),
    .Q_N(_11832_),
    .Q(\scanline[62][4] ));
 sg13g2_dfrbp_1 _29937_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net510),
    .D(_02265_),
    .Q_N(_11831_),
    .Q(\scanline[62][5] ));
 sg13g2_dfrbp_1 _29938_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net509),
    .D(_02266_),
    .Q_N(_11830_),
    .Q(\scanline[62][6] ));
 sg13g2_dfrbp_1 _29939_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net508),
    .D(_02267_),
    .Q_N(_11829_),
    .Q(\scanline[63][0] ));
 sg13g2_dfrbp_1 _29940_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net507),
    .D(_02268_),
    .Q_N(_11828_),
    .Q(\scanline[63][1] ));
 sg13g2_dfrbp_1 _29941_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net506),
    .D(_02269_),
    .Q_N(_11827_),
    .Q(\scanline[63][2] ));
 sg13g2_dfrbp_1 _29942_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net505),
    .D(_02270_),
    .Q_N(_11826_),
    .Q(\scanline[63][3] ));
 sg13g2_dfrbp_1 _29943_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net504),
    .D(_02271_),
    .Q_N(_11825_),
    .Q(\scanline[63][4] ));
 sg13g2_dfrbp_1 _29944_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net503),
    .D(_02272_),
    .Q_N(_11824_),
    .Q(\scanline[63][5] ));
 sg13g2_dfrbp_1 _29945_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net502),
    .D(_02273_),
    .Q_N(_11823_),
    .Q(\scanline[63][6] ));
 sg13g2_dfrbp_1 _29946_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net501),
    .D(_02274_),
    .Q_N(_11822_),
    .Q(\scanline[64][0] ));
 sg13g2_dfrbp_1 _29947_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net500),
    .D(_02275_),
    .Q_N(_11821_),
    .Q(\scanline[64][1] ));
 sg13g2_dfrbp_1 _29948_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net499),
    .D(_02276_),
    .Q_N(_11820_),
    .Q(\scanline[64][2] ));
 sg13g2_dfrbp_1 _29949_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net498),
    .D(_02277_),
    .Q_N(_11819_),
    .Q(\scanline[64][3] ));
 sg13g2_dfrbp_1 _29950_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net497),
    .D(_02278_),
    .Q_N(_11818_),
    .Q(\scanline[64][4] ));
 sg13g2_dfrbp_1 _29951_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net496),
    .D(_02279_),
    .Q_N(_11817_),
    .Q(\scanline[64][5] ));
 sg13g2_dfrbp_1 _29952_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net495),
    .D(_02280_),
    .Q_N(_11816_),
    .Q(\scanline[64][6] ));
 sg13g2_dfrbp_1 _29953_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net494),
    .D(_02281_),
    .Q_N(_11815_),
    .Q(\scanline[65][0] ));
 sg13g2_dfrbp_1 _29954_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net493),
    .D(_02282_),
    .Q_N(_11814_),
    .Q(\scanline[65][1] ));
 sg13g2_dfrbp_1 _29955_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net492),
    .D(_02283_),
    .Q_N(_11813_),
    .Q(\scanline[65][2] ));
 sg13g2_dfrbp_1 _29956_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net491),
    .D(_02284_),
    .Q_N(_11812_),
    .Q(\scanline[65][3] ));
 sg13g2_dfrbp_1 _29957_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net490),
    .D(_02285_),
    .Q_N(_11811_),
    .Q(\scanline[65][4] ));
 sg13g2_dfrbp_1 _29958_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net489),
    .D(_02286_),
    .Q_N(_11810_),
    .Q(\scanline[65][5] ));
 sg13g2_dfrbp_1 _29959_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net488),
    .D(_02287_),
    .Q_N(_11809_),
    .Q(\scanline[65][6] ));
 sg13g2_dfrbp_1 _29960_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net487),
    .D(_02288_),
    .Q_N(_11808_),
    .Q(\scanline[66][0] ));
 sg13g2_dfrbp_1 _29961_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net486),
    .D(_02289_),
    .Q_N(_11807_),
    .Q(\scanline[66][1] ));
 sg13g2_dfrbp_1 _29962_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net485),
    .D(_02290_),
    .Q_N(_11806_),
    .Q(\scanline[66][2] ));
 sg13g2_dfrbp_1 _29963_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net484),
    .D(_02291_),
    .Q_N(_11805_),
    .Q(\scanline[66][3] ));
 sg13g2_dfrbp_1 _29964_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net483),
    .D(_02292_),
    .Q_N(_11804_),
    .Q(\scanline[66][4] ));
 sg13g2_dfrbp_1 _29965_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net482),
    .D(_02293_),
    .Q_N(_11803_),
    .Q(\scanline[66][5] ));
 sg13g2_dfrbp_1 _29966_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net481),
    .D(_02294_),
    .Q_N(_11802_),
    .Q(\scanline[66][6] ));
 sg13g2_dfrbp_1 _29967_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net480),
    .D(_02295_),
    .Q_N(_11801_),
    .Q(\scanline[67][0] ));
 sg13g2_dfrbp_1 _29968_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net479),
    .D(_02296_),
    .Q_N(_11800_),
    .Q(\scanline[67][1] ));
 sg13g2_dfrbp_1 _29969_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net478),
    .D(_02297_),
    .Q_N(_11799_),
    .Q(\scanline[67][2] ));
 sg13g2_dfrbp_1 _29970_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net477),
    .D(_02298_),
    .Q_N(_11798_),
    .Q(\scanline[67][3] ));
 sg13g2_dfrbp_1 _29971_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net476),
    .D(_02299_),
    .Q_N(_11797_),
    .Q(\scanline[67][4] ));
 sg13g2_dfrbp_1 _29972_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net475),
    .D(_02300_),
    .Q_N(_11796_),
    .Q(\scanline[67][5] ));
 sg13g2_dfrbp_1 _29973_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net474),
    .D(_02301_),
    .Q_N(_11795_),
    .Q(\scanline[67][6] ));
 sg13g2_dfrbp_1 _29974_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net473),
    .D(_02302_),
    .Q_N(_11794_),
    .Q(\scanline[68][0] ));
 sg13g2_dfrbp_1 _29975_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net472),
    .D(_02303_),
    .Q_N(_11793_),
    .Q(\scanline[68][1] ));
 sg13g2_dfrbp_1 _29976_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net471),
    .D(_02304_),
    .Q_N(_11792_),
    .Q(\scanline[68][2] ));
 sg13g2_dfrbp_1 _29977_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net470),
    .D(_02305_),
    .Q_N(_11791_),
    .Q(\scanline[68][3] ));
 sg13g2_dfrbp_1 _29978_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net469),
    .D(_02306_),
    .Q_N(_11790_),
    .Q(\scanline[68][4] ));
 sg13g2_dfrbp_1 _29979_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net468),
    .D(_02307_),
    .Q_N(_11789_),
    .Q(\scanline[68][5] ));
 sg13g2_dfrbp_1 _29980_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net467),
    .D(_02308_),
    .Q_N(_11788_),
    .Q(\scanline[68][6] ));
 sg13g2_dfrbp_1 _29981_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net466),
    .D(_02309_),
    .Q_N(_11787_),
    .Q(\scanline[6][0] ));
 sg13g2_dfrbp_1 _29982_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net465),
    .D(_02310_),
    .Q_N(_11786_),
    .Q(\scanline[6][1] ));
 sg13g2_dfrbp_1 _29983_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net464),
    .D(_02311_),
    .Q_N(_11785_),
    .Q(\scanline[6][2] ));
 sg13g2_dfrbp_1 _29984_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net463),
    .D(_02312_),
    .Q_N(_11784_),
    .Q(\scanline[6][3] ));
 sg13g2_dfrbp_1 _29985_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net462),
    .D(_02313_),
    .Q_N(_11783_),
    .Q(\scanline[6][4] ));
 sg13g2_dfrbp_1 _29986_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net461),
    .D(_02314_),
    .Q_N(_11782_),
    .Q(\scanline[6][5] ));
 sg13g2_dfrbp_1 _29987_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net460),
    .D(_02315_),
    .Q_N(_11781_),
    .Q(\scanline[6][6] ));
 sg13g2_dfrbp_1 _29988_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net459),
    .D(_02316_),
    .Q_N(_11780_),
    .Q(\scanline[70][0] ));
 sg13g2_dfrbp_1 _29989_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net458),
    .D(_02317_),
    .Q_N(_11779_),
    .Q(\scanline[70][1] ));
 sg13g2_dfrbp_1 _29990_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net457),
    .D(_02318_),
    .Q_N(_11778_),
    .Q(\scanline[70][2] ));
 sg13g2_dfrbp_1 _29991_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net456),
    .D(_02319_),
    .Q_N(_11777_),
    .Q(\scanline[70][3] ));
 sg13g2_dfrbp_1 _29992_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net455),
    .D(_02320_),
    .Q_N(_11776_),
    .Q(\scanline[70][4] ));
 sg13g2_dfrbp_1 _29993_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net454),
    .D(_02321_),
    .Q_N(_11775_),
    .Q(\scanline[70][5] ));
 sg13g2_dfrbp_1 _29994_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net453),
    .D(_02322_),
    .Q_N(_11774_),
    .Q(\scanline[70][6] ));
 sg13g2_dfrbp_1 _29995_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net452),
    .D(_02323_),
    .Q_N(_11773_),
    .Q(\scanline[71][0] ));
 sg13g2_dfrbp_1 _29996_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net451),
    .D(_02324_),
    .Q_N(_11772_),
    .Q(\scanline[71][1] ));
 sg13g2_dfrbp_1 _29997_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net450),
    .D(_02325_),
    .Q_N(_11771_),
    .Q(\scanline[71][2] ));
 sg13g2_dfrbp_1 _29998_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net449),
    .D(_02326_),
    .Q_N(_11770_),
    .Q(\scanline[71][3] ));
 sg13g2_dfrbp_1 _29999_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net448),
    .D(_02327_),
    .Q_N(_11769_),
    .Q(\scanline[71][4] ));
 sg13g2_dfrbp_1 _30000_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net447),
    .D(_02328_),
    .Q_N(_11768_),
    .Q(\scanline[71][5] ));
 sg13g2_dfrbp_1 _30001_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net446),
    .D(_02329_),
    .Q_N(_11767_),
    .Q(\scanline[71][6] ));
 sg13g2_dfrbp_1 _30002_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net445),
    .D(_02330_),
    .Q_N(_11766_),
    .Q(\scanline[72][0] ));
 sg13g2_dfrbp_1 _30003_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net444),
    .D(_02331_),
    .Q_N(_11765_),
    .Q(\scanline[72][1] ));
 sg13g2_dfrbp_1 _30004_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net443),
    .D(_02332_),
    .Q_N(_11764_),
    .Q(\scanline[72][2] ));
 sg13g2_dfrbp_1 _30005_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net442),
    .D(_02333_),
    .Q_N(_11763_),
    .Q(\scanline[72][3] ));
 sg13g2_dfrbp_1 _30006_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net441),
    .D(_02334_),
    .Q_N(_11762_),
    .Q(\scanline[72][4] ));
 sg13g2_dfrbp_1 _30007_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net440),
    .D(_02335_),
    .Q_N(_11761_),
    .Q(\scanline[72][5] ));
 sg13g2_dfrbp_1 _30008_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net439),
    .D(_02336_),
    .Q_N(_11760_),
    .Q(\scanline[72][6] ));
 sg13g2_dfrbp_1 _30009_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net438),
    .D(_02337_),
    .Q_N(_11759_),
    .Q(\scanline[73][0] ));
 sg13g2_dfrbp_1 _30010_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net437),
    .D(_02338_),
    .Q_N(_11758_),
    .Q(\scanline[73][1] ));
 sg13g2_dfrbp_1 _30011_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net436),
    .D(_02339_),
    .Q_N(_11757_),
    .Q(\scanline[73][2] ));
 sg13g2_dfrbp_1 _30012_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net435),
    .D(_02340_),
    .Q_N(_11756_),
    .Q(\scanline[73][3] ));
 sg13g2_dfrbp_1 _30013_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net434),
    .D(_02341_),
    .Q_N(_11755_),
    .Q(\scanline[73][4] ));
 sg13g2_dfrbp_1 _30014_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net433),
    .D(_02342_),
    .Q_N(_11754_),
    .Q(\scanline[73][5] ));
 sg13g2_dfrbp_1 _30015_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net432),
    .D(_02343_),
    .Q_N(_11753_),
    .Q(\scanline[73][6] ));
 sg13g2_dfrbp_1 _30016_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net431),
    .D(_02344_),
    .Q_N(_11752_),
    .Q(\scanline[74][0] ));
 sg13g2_dfrbp_1 _30017_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net430),
    .D(_02345_),
    .Q_N(_11751_),
    .Q(\scanline[74][1] ));
 sg13g2_dfrbp_1 _30018_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net429),
    .D(_02346_),
    .Q_N(_11750_),
    .Q(\scanline[74][2] ));
 sg13g2_dfrbp_1 _30019_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net428),
    .D(_02347_),
    .Q_N(_11749_),
    .Q(\scanline[74][3] ));
 sg13g2_dfrbp_1 _30020_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net427),
    .D(_02348_),
    .Q_N(_11748_),
    .Q(\scanline[74][4] ));
 sg13g2_dfrbp_1 _30021_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net426),
    .D(_02349_),
    .Q_N(_11747_),
    .Q(\scanline[74][5] ));
 sg13g2_dfrbp_1 _30022_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net425),
    .D(_02350_),
    .Q_N(_11746_),
    .Q(\scanline[74][6] ));
 sg13g2_dfrbp_1 _30023_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net424),
    .D(_02351_),
    .Q_N(_11745_),
    .Q(\scanline[75][0] ));
 sg13g2_dfrbp_1 _30024_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net423),
    .D(_02352_),
    .Q_N(_11744_),
    .Q(\scanline[75][1] ));
 sg13g2_dfrbp_1 _30025_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net422),
    .D(_02353_),
    .Q_N(_11743_),
    .Q(\scanline[75][2] ));
 sg13g2_dfrbp_1 _30026_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net421),
    .D(_02354_),
    .Q_N(_11742_),
    .Q(\scanline[75][3] ));
 sg13g2_dfrbp_1 _30027_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net420),
    .D(_02355_),
    .Q_N(_11741_),
    .Q(\scanline[75][4] ));
 sg13g2_dfrbp_1 _30028_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net419),
    .D(_02356_),
    .Q_N(_11740_),
    .Q(\scanline[75][5] ));
 sg13g2_dfrbp_1 _30029_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net418),
    .D(_02357_),
    .Q_N(_11739_),
    .Q(\scanline[75][6] ));
 sg13g2_dfrbp_1 _30030_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net417),
    .D(_02358_),
    .Q_N(_11738_),
    .Q(\scanline[76][0] ));
 sg13g2_dfrbp_1 _30031_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net416),
    .D(_02359_),
    .Q_N(_11737_),
    .Q(\scanline[76][1] ));
 sg13g2_dfrbp_1 _30032_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net415),
    .D(_02360_),
    .Q_N(_11736_),
    .Q(\scanline[76][2] ));
 sg13g2_dfrbp_1 _30033_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net414),
    .D(_02361_),
    .Q_N(_11735_),
    .Q(\scanline[76][3] ));
 sg13g2_dfrbp_1 _30034_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net413),
    .D(_02362_),
    .Q_N(_11734_),
    .Q(\scanline[76][4] ));
 sg13g2_dfrbp_1 _30035_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net412),
    .D(_02363_),
    .Q_N(_11733_),
    .Q(\scanline[76][5] ));
 sg13g2_dfrbp_1 _30036_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net411),
    .D(_02364_),
    .Q_N(_11732_),
    .Q(\scanline[76][6] ));
 sg13g2_dfrbp_1 _30037_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net410),
    .D(_02365_),
    .Q_N(_11731_),
    .Q(\scanline[77][0] ));
 sg13g2_dfrbp_1 _30038_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net409),
    .D(_02366_),
    .Q_N(_11730_),
    .Q(\scanline[77][1] ));
 sg13g2_dfrbp_1 _30039_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net408),
    .D(_02367_),
    .Q_N(_11729_),
    .Q(\scanline[77][2] ));
 sg13g2_dfrbp_1 _30040_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net407),
    .D(_02368_),
    .Q_N(_11728_),
    .Q(\scanline[77][3] ));
 sg13g2_dfrbp_1 _30041_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net406),
    .D(_02369_),
    .Q_N(_11727_),
    .Q(\scanline[77][4] ));
 sg13g2_dfrbp_1 _30042_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net405),
    .D(_02370_),
    .Q_N(_11726_),
    .Q(\scanline[77][5] ));
 sg13g2_dfrbp_1 _30043_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net404),
    .D(_02371_),
    .Q_N(_11725_),
    .Q(\scanline[77][6] ));
 sg13g2_dfrbp_1 _30044_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net403),
    .D(_02372_),
    .Q_N(_11724_),
    .Q(\scanline[78][0] ));
 sg13g2_dfrbp_1 _30045_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net402),
    .D(_02373_),
    .Q_N(_11723_),
    .Q(\scanline[78][1] ));
 sg13g2_dfrbp_1 _30046_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net401),
    .D(_02374_),
    .Q_N(_11722_),
    .Q(\scanline[78][2] ));
 sg13g2_dfrbp_1 _30047_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net400),
    .D(_02375_),
    .Q_N(_11721_),
    .Q(\scanline[78][3] ));
 sg13g2_dfrbp_1 _30048_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net399),
    .D(_02376_),
    .Q_N(_11720_),
    .Q(\scanline[78][4] ));
 sg13g2_dfrbp_1 _30049_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net398),
    .D(_02377_),
    .Q_N(_11719_),
    .Q(\scanline[78][5] ));
 sg13g2_dfrbp_1 _30050_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net397),
    .D(_02378_),
    .Q_N(_11718_),
    .Q(\scanline[78][6] ));
 sg13g2_dfrbp_1 _30051_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net396),
    .D(_02379_),
    .Q_N(_11717_),
    .Q(\scanline[7][0] ));
 sg13g2_dfrbp_1 _30052_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net395),
    .D(_02380_),
    .Q_N(_11716_),
    .Q(\scanline[7][1] ));
 sg13g2_dfrbp_1 _30053_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net394),
    .D(_02381_),
    .Q_N(_11715_),
    .Q(\scanline[7][2] ));
 sg13g2_dfrbp_1 _30054_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net393),
    .D(_02382_),
    .Q_N(_11714_),
    .Q(\scanline[7][3] ));
 sg13g2_dfrbp_1 _30055_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net392),
    .D(_02383_),
    .Q_N(_11713_),
    .Q(\scanline[7][4] ));
 sg13g2_dfrbp_1 _30056_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net391),
    .D(_02384_),
    .Q_N(_11712_),
    .Q(\scanline[7][5] ));
 sg13g2_dfrbp_1 _30057_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net390),
    .D(_02385_),
    .Q_N(_11711_),
    .Q(\scanline[7][6] ));
 sg13g2_dfrbp_1 _30058_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net389),
    .D(_02386_),
    .Q_N(_11710_),
    .Q(\scanline[80][0] ));
 sg13g2_dfrbp_1 _30059_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net388),
    .D(_02387_),
    .Q_N(_11709_),
    .Q(\scanline[80][1] ));
 sg13g2_dfrbp_1 _30060_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net387),
    .D(_02388_),
    .Q_N(_11708_),
    .Q(\scanline[80][2] ));
 sg13g2_dfrbp_1 _30061_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net386),
    .D(_02389_),
    .Q_N(_11707_),
    .Q(\scanline[80][3] ));
 sg13g2_dfrbp_1 _30062_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net385),
    .D(_02390_),
    .Q_N(_11706_),
    .Q(\scanline[80][4] ));
 sg13g2_dfrbp_1 _30063_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net384),
    .D(_02391_),
    .Q_N(_11705_),
    .Q(\scanline[80][5] ));
 sg13g2_dfrbp_1 _30064_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net383),
    .D(_02392_),
    .Q_N(_11704_),
    .Q(\scanline[80][6] ));
 sg13g2_dfrbp_1 _30065_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net382),
    .D(_02393_),
    .Q_N(_11703_),
    .Q(\scanline[81][0] ));
 sg13g2_dfrbp_1 _30066_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net381),
    .D(_02394_),
    .Q_N(_11702_),
    .Q(\scanline[81][1] ));
 sg13g2_dfrbp_1 _30067_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net380),
    .D(_02395_),
    .Q_N(_11701_),
    .Q(\scanline[81][2] ));
 sg13g2_dfrbp_1 _30068_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net379),
    .D(_02396_),
    .Q_N(_11700_),
    .Q(\scanline[81][3] ));
 sg13g2_dfrbp_1 _30069_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net378),
    .D(_02397_),
    .Q_N(_11699_),
    .Q(\scanline[81][4] ));
 sg13g2_dfrbp_1 _30070_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net377),
    .D(_02398_),
    .Q_N(_11698_),
    .Q(\scanline[81][5] ));
 sg13g2_dfrbp_1 _30071_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net376),
    .D(_02399_),
    .Q_N(_11697_),
    .Q(\scanline[81][6] ));
 sg13g2_dfrbp_1 _30072_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net375),
    .D(_02400_),
    .Q_N(_11696_),
    .Q(\scanline[82][0] ));
 sg13g2_dfrbp_1 _30073_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net374),
    .D(_02401_),
    .Q_N(_11695_),
    .Q(\scanline[82][1] ));
 sg13g2_dfrbp_1 _30074_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net373),
    .D(_02402_),
    .Q_N(_11694_),
    .Q(\scanline[82][2] ));
 sg13g2_dfrbp_1 _30075_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net372),
    .D(_02403_),
    .Q_N(_11693_),
    .Q(\scanline[82][3] ));
 sg13g2_dfrbp_1 _30076_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net371),
    .D(_02404_),
    .Q_N(_11692_),
    .Q(\scanline[82][4] ));
 sg13g2_dfrbp_1 _30077_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net370),
    .D(_02405_),
    .Q_N(_11691_),
    .Q(\scanline[82][5] ));
 sg13g2_dfrbp_1 _30078_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net369),
    .D(_02406_),
    .Q_N(_11690_),
    .Q(\scanline[82][6] ));
 sg13g2_dfrbp_1 _30079_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net368),
    .D(_02407_),
    .Q_N(_11689_),
    .Q(\scanline[83][0] ));
 sg13g2_dfrbp_1 _30080_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net367),
    .D(_02408_),
    .Q_N(_11688_),
    .Q(\scanline[83][1] ));
 sg13g2_dfrbp_1 _30081_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net366),
    .D(_02409_),
    .Q_N(_11687_),
    .Q(\scanline[83][2] ));
 sg13g2_dfrbp_1 _30082_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net365),
    .D(_02410_),
    .Q_N(_11686_),
    .Q(\scanline[83][3] ));
 sg13g2_dfrbp_1 _30083_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net364),
    .D(_02411_),
    .Q_N(_11685_),
    .Q(\scanline[83][4] ));
 sg13g2_dfrbp_1 _30084_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net363),
    .D(_02412_),
    .Q_N(_11684_),
    .Q(\scanline[83][5] ));
 sg13g2_dfrbp_1 _30085_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net362),
    .D(_02413_),
    .Q_N(_11683_),
    .Q(\scanline[83][6] ));
 sg13g2_dfrbp_1 _30086_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net361),
    .D(_02414_),
    .Q_N(_11682_),
    .Q(\scanline[84][0] ));
 sg13g2_dfrbp_1 _30087_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net360),
    .D(_02415_),
    .Q_N(_11681_),
    .Q(\scanline[84][1] ));
 sg13g2_dfrbp_1 _30088_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net359),
    .D(_02416_),
    .Q_N(_11680_),
    .Q(\scanline[84][2] ));
 sg13g2_dfrbp_1 _30089_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net358),
    .D(_02417_),
    .Q_N(_11679_),
    .Q(\scanline[84][3] ));
 sg13g2_dfrbp_1 _30090_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net357),
    .D(_02418_),
    .Q_N(_11678_),
    .Q(\scanline[84][4] ));
 sg13g2_dfrbp_1 _30091_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net356),
    .D(_02419_),
    .Q_N(_11677_),
    .Q(\scanline[84][5] ));
 sg13g2_dfrbp_1 _30092_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net355),
    .D(_02420_),
    .Q_N(_11676_),
    .Q(\scanline[84][6] ));
 sg13g2_dfrbp_1 _30093_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net354),
    .D(_02421_),
    .Q_N(_11675_),
    .Q(\scanline[85][0] ));
 sg13g2_dfrbp_1 _30094_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net353),
    .D(_02422_),
    .Q_N(_11674_),
    .Q(\scanline[85][1] ));
 sg13g2_dfrbp_1 _30095_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net352),
    .D(_02423_),
    .Q_N(_11673_),
    .Q(\scanline[85][2] ));
 sg13g2_dfrbp_1 _30096_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net351),
    .D(_02424_),
    .Q_N(_11672_),
    .Q(\scanline[85][3] ));
 sg13g2_dfrbp_1 _30097_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net350),
    .D(_02425_),
    .Q_N(_11671_),
    .Q(\scanline[85][4] ));
 sg13g2_dfrbp_1 _30098_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net349),
    .D(_02426_),
    .Q_N(_11670_),
    .Q(\scanline[85][5] ));
 sg13g2_dfrbp_1 _30099_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net348),
    .D(_02427_),
    .Q_N(_11669_),
    .Q(\scanline[85][6] ));
 sg13g2_dfrbp_1 _30100_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net347),
    .D(_02428_),
    .Q_N(_11668_),
    .Q(\scanline[86][0] ));
 sg13g2_dfrbp_1 _30101_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net346),
    .D(_02429_),
    .Q_N(_11667_),
    .Q(\scanline[86][1] ));
 sg13g2_dfrbp_1 _30102_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net345),
    .D(_02430_),
    .Q_N(_11666_),
    .Q(\scanline[86][2] ));
 sg13g2_dfrbp_1 _30103_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net344),
    .D(_02431_),
    .Q_N(_11665_),
    .Q(\scanline[86][3] ));
 sg13g2_dfrbp_1 _30104_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net343),
    .D(_02432_),
    .Q_N(_11664_),
    .Q(\scanline[86][4] ));
 sg13g2_dfrbp_1 _30105_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net342),
    .D(_02433_),
    .Q_N(_11663_),
    .Q(\scanline[86][5] ));
 sg13g2_dfrbp_1 _30106_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net341),
    .D(_02434_),
    .Q_N(_11662_),
    .Q(\scanline[86][6] ));
 sg13g2_dfrbp_1 _30107_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net340),
    .D(_02435_),
    .Q_N(_11661_),
    .Q(\scanline[87][0] ));
 sg13g2_dfrbp_1 _30108_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net339),
    .D(_02436_),
    .Q_N(_11660_),
    .Q(\scanline[87][1] ));
 sg13g2_dfrbp_1 _30109_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net338),
    .D(_02437_),
    .Q_N(_11659_),
    .Q(\scanline[87][2] ));
 sg13g2_dfrbp_1 _30110_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net337),
    .D(_02438_),
    .Q_N(_11658_),
    .Q(\scanline[87][3] ));
 sg13g2_dfrbp_1 _30111_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net336),
    .D(_02439_),
    .Q_N(_11657_),
    .Q(\scanline[87][4] ));
 sg13g2_dfrbp_1 _30112_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net335),
    .D(_02440_),
    .Q_N(_11656_),
    .Q(\scanline[87][5] ));
 sg13g2_dfrbp_1 _30113_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net334),
    .D(_02441_),
    .Q_N(_11655_),
    .Q(\scanline[87][6] ));
 sg13g2_dfrbp_1 _30114_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net333),
    .D(_02442_),
    .Q_N(_11654_),
    .Q(\scanline[88][0] ));
 sg13g2_dfrbp_1 _30115_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net332),
    .D(_02443_),
    .Q_N(_11653_),
    .Q(\scanline[88][1] ));
 sg13g2_dfrbp_1 _30116_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net331),
    .D(_02444_),
    .Q_N(_11652_),
    .Q(\scanline[88][2] ));
 sg13g2_dfrbp_1 _30117_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net330),
    .D(_02445_),
    .Q_N(_11651_),
    .Q(\scanline[88][3] ));
 sg13g2_dfrbp_1 _30118_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net329),
    .D(_02446_),
    .Q_N(_11650_),
    .Q(\scanline[88][4] ));
 sg13g2_dfrbp_1 _30119_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net328),
    .D(_02447_),
    .Q_N(_11649_),
    .Q(\scanline[88][5] ));
 sg13g2_dfrbp_1 _30120_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net327),
    .D(_02448_),
    .Q_N(_11648_),
    .Q(\scanline[88][6] ));
 sg13g2_dfrbp_1 _30121_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net326),
    .D(_02449_),
    .Q_N(_11647_),
    .Q(\scanline[8][0] ));
 sg13g2_dfrbp_1 _30122_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net325),
    .D(_02450_),
    .Q_N(_11646_),
    .Q(\scanline[8][1] ));
 sg13g2_dfrbp_1 _30123_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net324),
    .D(_02451_),
    .Q_N(_11645_),
    .Q(\scanline[8][2] ));
 sg13g2_dfrbp_1 _30124_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net323),
    .D(_02452_),
    .Q_N(_11644_),
    .Q(\scanline[8][3] ));
 sg13g2_dfrbp_1 _30125_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net322),
    .D(_02453_),
    .Q_N(_11643_),
    .Q(\scanline[8][4] ));
 sg13g2_dfrbp_1 _30126_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net321),
    .D(_02454_),
    .Q_N(_11642_),
    .Q(\scanline[8][5] ));
 sg13g2_dfrbp_1 _30127_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net320),
    .D(_02455_),
    .Q_N(_11641_),
    .Q(\scanline[8][6] ));
 sg13g2_dfrbp_1 _30128_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net319),
    .D(_02456_),
    .Q_N(_11640_),
    .Q(\scanline[90][0] ));
 sg13g2_dfrbp_1 _30129_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net318),
    .D(_02457_),
    .Q_N(_11639_),
    .Q(\scanline[90][1] ));
 sg13g2_dfrbp_1 _30130_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net317),
    .D(_02458_),
    .Q_N(_11638_),
    .Q(\scanline[90][2] ));
 sg13g2_dfrbp_1 _30131_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net316),
    .D(_02459_),
    .Q_N(_11637_),
    .Q(\scanline[90][3] ));
 sg13g2_dfrbp_1 _30132_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net315),
    .D(_02460_),
    .Q_N(_11636_),
    .Q(\scanline[90][4] ));
 sg13g2_dfrbp_1 _30133_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net314),
    .D(_02461_),
    .Q_N(_11635_),
    .Q(\scanline[90][5] ));
 sg13g2_dfrbp_1 _30134_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net313),
    .D(_02462_),
    .Q_N(_11634_),
    .Q(\scanline[90][6] ));
 sg13g2_dfrbp_1 _30135_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net312),
    .D(_02463_),
    .Q_N(_11633_),
    .Q(\scanline[91][0] ));
 sg13g2_dfrbp_1 _30136_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net311),
    .D(_02464_),
    .Q_N(_11632_),
    .Q(\scanline[91][1] ));
 sg13g2_dfrbp_1 _30137_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net310),
    .D(_02465_),
    .Q_N(_11631_),
    .Q(\scanline[91][2] ));
 sg13g2_dfrbp_1 _30138_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net309),
    .D(_02466_),
    .Q_N(_11630_),
    .Q(\scanline[91][3] ));
 sg13g2_dfrbp_1 _30139_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net308),
    .D(_02467_),
    .Q_N(_11629_),
    .Q(\scanline[91][4] ));
 sg13g2_dfrbp_1 _30140_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net300),
    .D(_02468_),
    .Q_N(_11628_),
    .Q(\scanline[91][5] ));
 sg13g2_dfrbp_1 _30141_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net299),
    .D(_02469_),
    .Q_N(_11627_),
    .Q(\scanline[91][6] ));
 sg13g2_dfrbp_1 _30142_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net298),
    .D(_02470_),
    .Q_N(_11626_),
    .Q(\scanline[92][0] ));
 sg13g2_dfrbp_1 _30143_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net297),
    .D(_02471_),
    .Q_N(_11625_),
    .Q(\scanline[92][1] ));
 sg13g2_dfrbp_1 _30144_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net296),
    .D(_02472_),
    .Q_N(_11624_),
    .Q(\scanline[92][2] ));
 sg13g2_dfrbp_1 _30145_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net295),
    .D(_02473_),
    .Q_N(_11623_),
    .Q(\scanline[92][3] ));
 sg13g2_dfrbp_1 _30146_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net294),
    .D(_02474_),
    .Q_N(_11622_),
    .Q(\scanline[92][4] ));
 sg13g2_dfrbp_1 _30147_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net293),
    .D(_02475_),
    .Q_N(_11621_),
    .Q(\scanline[92][5] ));
 sg13g2_dfrbp_1 _30148_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net292),
    .D(_02476_),
    .Q_N(_11620_),
    .Q(\scanline[92][6] ));
 sg13g2_dfrbp_1 _30149_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net291),
    .D(_02477_),
    .Q_N(_11619_),
    .Q(\scanline[93][0] ));
 sg13g2_dfrbp_1 _30150_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net290),
    .D(_02478_),
    .Q_N(_11618_),
    .Q(\scanline[93][1] ));
 sg13g2_dfrbp_1 _30151_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net289),
    .D(_02479_),
    .Q_N(_11617_),
    .Q(\scanline[93][2] ));
 sg13g2_dfrbp_1 _30152_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net288),
    .D(_02480_),
    .Q_N(_11616_),
    .Q(\scanline[93][3] ));
 sg13g2_dfrbp_1 _30153_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net287),
    .D(_02481_),
    .Q_N(_11615_),
    .Q(\scanline[93][4] ));
 sg13g2_dfrbp_1 _30154_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net286),
    .D(_02482_),
    .Q_N(_11614_),
    .Q(\scanline[93][5] ));
 sg13g2_dfrbp_1 _30155_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net285),
    .D(_02483_),
    .Q_N(_11613_),
    .Q(\scanline[93][6] ));
 sg13g2_dfrbp_1 _30156_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net284),
    .D(_02484_),
    .Q_N(_11612_),
    .Q(\scanline[94][0] ));
 sg13g2_dfrbp_1 _30157_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net283),
    .D(_02485_),
    .Q_N(_11611_),
    .Q(\scanline[94][1] ));
 sg13g2_dfrbp_1 _30158_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net282),
    .D(_02486_),
    .Q_N(_11610_),
    .Q(\scanline[94][2] ));
 sg13g2_dfrbp_1 _30159_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net281),
    .D(_02487_),
    .Q_N(_11609_),
    .Q(\scanline[94][3] ));
 sg13g2_dfrbp_1 _30160_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net280),
    .D(_02488_),
    .Q_N(_11608_),
    .Q(\scanline[94][4] ));
 sg13g2_dfrbp_1 _30161_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net279),
    .D(_02489_),
    .Q_N(_11607_),
    .Q(\scanline[94][5] ));
 sg13g2_dfrbp_1 _30162_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net278),
    .D(_02490_),
    .Q_N(_11606_),
    .Q(\scanline[94][6] ));
 sg13g2_dfrbp_1 _30163_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net277),
    .D(_02491_),
    .Q_N(_11605_),
    .Q(\scanline[95][0] ));
 sg13g2_dfrbp_1 _30164_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net276),
    .D(_02492_),
    .Q_N(_11604_),
    .Q(\scanline[95][1] ));
 sg13g2_dfrbp_1 _30165_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net275),
    .D(_02493_),
    .Q_N(_11603_),
    .Q(\scanline[95][2] ));
 sg13g2_dfrbp_1 _30166_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net274),
    .D(_02494_),
    .Q_N(_11602_),
    .Q(\scanline[95][3] ));
 sg13g2_dfrbp_1 _30167_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net273),
    .D(_02495_),
    .Q_N(_11601_),
    .Q(\scanline[95][4] ));
 sg13g2_dfrbp_1 _30168_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net272),
    .D(_02496_),
    .Q_N(_11600_),
    .Q(\scanline[95][5] ));
 sg13g2_dfrbp_1 _30169_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net271),
    .D(_02497_),
    .Q_N(_11599_),
    .Q(\scanline[95][6] ));
 sg13g2_dfrbp_1 _30170_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net270),
    .D(_02498_),
    .Q_N(_11598_),
    .Q(\scanline[96][0] ));
 sg13g2_dfrbp_1 _30171_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net269),
    .D(_02499_),
    .Q_N(_11597_),
    .Q(\scanline[96][1] ));
 sg13g2_dfrbp_1 _30172_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net268),
    .D(_02500_),
    .Q_N(_11596_),
    .Q(\scanline[96][2] ));
 sg13g2_dfrbp_1 _30173_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net267),
    .D(_02501_),
    .Q_N(_11595_),
    .Q(\scanline[96][3] ));
 sg13g2_dfrbp_1 _30174_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net266),
    .D(_02502_),
    .Q_N(_11594_),
    .Q(\scanline[96][4] ));
 sg13g2_dfrbp_1 _30175_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net265),
    .D(_02503_),
    .Q_N(_11593_),
    .Q(\scanline[96][5] ));
 sg13g2_dfrbp_1 _30176_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net264),
    .D(_02504_),
    .Q_N(_11592_),
    .Q(\scanline[96][6] ));
 sg13g2_dfrbp_1 _30177_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net263),
    .D(_02505_),
    .Q_N(_11591_),
    .Q(\scanline[97][0] ));
 sg13g2_dfrbp_1 _30178_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net262),
    .D(_02506_),
    .Q_N(_11590_),
    .Q(\scanline[97][1] ));
 sg13g2_dfrbp_1 _30179_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net261),
    .D(_02507_),
    .Q_N(_11589_),
    .Q(\scanline[97][2] ));
 sg13g2_dfrbp_1 _30180_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net260),
    .D(_02508_),
    .Q_N(_11588_),
    .Q(\scanline[97][3] ));
 sg13g2_dfrbp_1 _30181_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net259),
    .D(_02509_),
    .Q_N(_11587_),
    .Q(\scanline[97][4] ));
 sg13g2_dfrbp_1 _30182_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net258),
    .D(_02510_),
    .Q_N(_11586_),
    .Q(\scanline[97][5] ));
 sg13g2_dfrbp_1 _30183_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net257),
    .D(_02511_),
    .Q_N(_11585_),
    .Q(\scanline[97][6] ));
 sg13g2_dfrbp_1 _30184_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net256),
    .D(_02512_),
    .Q_N(_11584_),
    .Q(\scanline[98][0] ));
 sg13g2_dfrbp_1 _30185_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net255),
    .D(_02513_),
    .Q_N(_11583_),
    .Q(\scanline[98][1] ));
 sg13g2_dfrbp_1 _30186_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net254),
    .D(_02514_),
    .Q_N(_11582_),
    .Q(\scanline[98][2] ));
 sg13g2_dfrbp_1 _30187_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net253),
    .D(_02515_),
    .Q_N(_11581_),
    .Q(\scanline[98][3] ));
 sg13g2_dfrbp_1 _30188_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net252),
    .D(_02516_),
    .Q_N(_11580_),
    .Q(\scanline[98][4] ));
 sg13g2_dfrbp_1 _30189_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net251),
    .D(_02517_),
    .Q_N(_11579_),
    .Q(\scanline[98][5] ));
 sg13g2_dfrbp_1 _30190_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net250),
    .D(_02518_),
    .Q_N(_11578_),
    .Q(\scanline[98][6] ));
 sg13g2_dfrbp_1 _30191_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net249),
    .D(_02519_),
    .Q_N(_11577_),
    .Q(\scanline[0][0] ));
 sg13g2_dfrbp_1 _30192_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net248),
    .D(_02520_),
    .Q_N(_11576_),
    .Q(\scanline[0][1] ));
 sg13g2_dfrbp_1 _30193_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net247),
    .D(_02521_),
    .Q_N(_11575_),
    .Q(\scanline[0][2] ));
 sg13g2_dfrbp_1 _30194_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net246),
    .D(_02522_),
    .Q_N(_11574_),
    .Q(\scanline[0][3] ));
 sg13g2_dfrbp_1 _30195_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net245),
    .D(_02523_),
    .Q_N(_11573_),
    .Q(\scanline[0][4] ));
 sg13g2_dfrbp_1 _30196_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net244),
    .D(_02524_),
    .Q_N(_11572_),
    .Q(\scanline[0][5] ));
 sg13g2_dfrbp_1 _30197_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net243),
    .D(_02525_),
    .Q_N(_11571_),
    .Q(\scanline[0][6] ));
 sg13g2_dfrbp_1 _30198_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net242),
    .D(_02526_),
    .Q_N(_11570_),
    .Q(\scanline[100][0] ));
 sg13g2_dfrbp_1 _30199_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net241),
    .D(_02527_),
    .Q_N(_11569_),
    .Q(\scanline[100][1] ));
 sg13g2_dfrbp_1 _30200_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net240),
    .D(_02528_),
    .Q_N(_11568_),
    .Q(\scanline[100][2] ));
 sg13g2_dfrbp_1 _30201_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net239),
    .D(_02529_),
    .Q_N(_11567_),
    .Q(\scanline[100][3] ));
 sg13g2_dfrbp_1 _30202_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net238),
    .D(_02530_),
    .Q_N(_11566_),
    .Q(\scanline[100][4] ));
 sg13g2_dfrbp_1 _30203_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net237),
    .D(_02531_),
    .Q_N(_11565_),
    .Q(\scanline[100][5] ));
 sg13g2_dfrbp_1 _30204_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net236),
    .D(_02532_),
    .Q_N(_11564_),
    .Q(\scanline[100][6] ));
 sg13g2_dfrbp_1 _30205_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net235),
    .D(_02533_),
    .Q_N(_11563_),
    .Q(\scanline[101][0] ));
 sg13g2_dfrbp_1 _30206_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net234),
    .D(_02534_),
    .Q_N(_11562_),
    .Q(\scanline[101][1] ));
 sg13g2_dfrbp_1 _30207_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net233),
    .D(_02535_),
    .Q_N(_11561_),
    .Q(\scanline[101][2] ));
 sg13g2_dfrbp_1 _30208_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net232),
    .D(_02536_),
    .Q_N(_11560_),
    .Q(\scanline[101][3] ));
 sg13g2_dfrbp_1 _30209_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net231),
    .D(_02537_),
    .Q_N(_11559_),
    .Q(\scanline[101][4] ));
 sg13g2_dfrbp_1 _30210_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net230),
    .D(_02538_),
    .Q_N(_11558_),
    .Q(\scanline[101][5] ));
 sg13g2_dfrbp_1 _30211_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net229),
    .D(_02539_),
    .Q_N(_11557_),
    .Q(\scanline[101][6] ));
 sg13g2_dfrbp_1 _30212_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net228),
    .D(_02540_),
    .Q_N(_11556_),
    .Q(\scanline[102][0] ));
 sg13g2_dfrbp_1 _30213_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net227),
    .D(_02541_),
    .Q_N(_11555_),
    .Q(\scanline[102][1] ));
 sg13g2_dfrbp_1 _30214_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net226),
    .D(_02542_),
    .Q_N(_11554_),
    .Q(\scanline[102][2] ));
 sg13g2_dfrbp_1 _30215_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net225),
    .D(_02543_),
    .Q_N(_11553_),
    .Q(\scanline[102][3] ));
 sg13g2_dfrbp_1 _30216_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net224),
    .D(_02544_),
    .Q_N(_11552_),
    .Q(\scanline[102][4] ));
 sg13g2_dfrbp_1 _30217_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net223),
    .D(_02545_),
    .Q_N(_11551_),
    .Q(\scanline[102][5] ));
 sg13g2_dfrbp_1 _30218_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net222),
    .D(_02546_),
    .Q_N(_11550_),
    .Q(\scanline[102][6] ));
 sg13g2_dfrbp_1 _30219_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net221),
    .D(_02547_),
    .Q_N(_11549_),
    .Q(\scanline[103][0] ));
 sg13g2_dfrbp_1 _30220_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net220),
    .D(_02548_),
    .Q_N(_11548_),
    .Q(\scanline[103][1] ));
 sg13g2_dfrbp_1 _30221_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net217),
    .D(_02549_),
    .Q_N(_11547_),
    .Q(\scanline[103][2] ));
 sg13g2_dfrbp_1 _30222_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net216),
    .D(_02550_),
    .Q_N(_11546_),
    .Q(\scanline[103][3] ));
 sg13g2_dfrbp_1 _30223_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net215),
    .D(_02551_),
    .Q_N(_11545_),
    .Q(\scanline[103][4] ));
 sg13g2_dfrbp_1 _30224_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net214),
    .D(_02552_),
    .Q_N(_11544_),
    .Q(\scanline[103][5] ));
 sg13g2_dfrbp_1 _30225_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net213),
    .D(_02553_),
    .Q_N(_11543_),
    .Q(\scanline[103][6] ));
 sg13g2_dfrbp_1 _30226_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net212),
    .D(_02554_),
    .Q_N(_11542_),
    .Q(\scanline[104][0] ));
 sg13g2_dfrbp_1 _30227_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net211),
    .D(_02555_),
    .Q_N(_11541_),
    .Q(\scanline[104][1] ));
 sg13g2_dfrbp_1 _30228_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net210),
    .D(_02556_),
    .Q_N(_11540_),
    .Q(\scanline[104][2] ));
 sg13g2_dfrbp_1 _30229_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net209),
    .D(_02557_),
    .Q_N(_11539_),
    .Q(\scanline[104][3] ));
 sg13g2_dfrbp_1 _30230_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net208),
    .D(_02558_),
    .Q_N(_11538_),
    .Q(\scanline[104][4] ));
 sg13g2_dfrbp_1 _30231_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net207),
    .D(_02559_),
    .Q_N(_11537_),
    .Q(\scanline[104][5] ));
 sg13g2_dfrbp_1 _30232_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net206),
    .D(_02560_),
    .Q_N(_11536_),
    .Q(\scanline[104][6] ));
 sg13g2_dfrbp_1 _30233_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net205),
    .D(_02561_),
    .Q_N(_11535_),
    .Q(\scanline[105][0] ));
 sg13g2_dfrbp_1 _30234_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net204),
    .D(_02562_),
    .Q_N(_11534_),
    .Q(\scanline[105][1] ));
 sg13g2_dfrbp_1 _30235_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net203),
    .D(_02563_),
    .Q_N(_11533_),
    .Q(\scanline[105][2] ));
 sg13g2_dfrbp_1 _30236_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net202),
    .D(_02564_),
    .Q_N(_11532_),
    .Q(\scanline[105][3] ));
 sg13g2_dfrbp_1 _30237_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net201),
    .D(_02565_),
    .Q_N(_11531_),
    .Q(\scanline[105][4] ));
 sg13g2_dfrbp_1 _30238_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net200),
    .D(_02566_),
    .Q_N(_11530_),
    .Q(\scanline[105][5] ));
 sg13g2_dfrbp_1 _30239_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net199),
    .D(_02567_),
    .Q_N(_11529_),
    .Q(\scanline[105][6] ));
 sg13g2_dfrbp_1 _30240_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net198),
    .D(_02568_),
    .Q_N(_11528_),
    .Q(\scanline[106][0] ));
 sg13g2_dfrbp_1 _30241_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net197),
    .D(_02569_),
    .Q_N(_11527_),
    .Q(\scanline[106][1] ));
 sg13g2_dfrbp_1 _30242_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net196),
    .D(_02570_),
    .Q_N(_11526_),
    .Q(\scanline[106][2] ));
 sg13g2_dfrbp_1 _30243_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net195),
    .D(_02571_),
    .Q_N(_11525_),
    .Q(\scanline[106][3] ));
 sg13g2_dfrbp_1 _30244_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net194),
    .D(_02572_),
    .Q_N(_11524_),
    .Q(\scanline[106][4] ));
 sg13g2_dfrbp_1 _30245_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net193),
    .D(_02573_),
    .Q_N(_11523_),
    .Q(\scanline[106][5] ));
 sg13g2_dfrbp_1 _30246_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net192),
    .D(_02574_),
    .Q_N(_11522_),
    .Q(\scanline[106][6] ));
 sg13g2_dfrbp_1 _30247_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net191),
    .D(_02575_),
    .Q_N(_11521_),
    .Q(\scanline[107][0] ));
 sg13g2_dfrbp_1 _30248_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net190),
    .D(_02576_),
    .Q_N(_11520_),
    .Q(\scanline[107][1] ));
 sg13g2_dfrbp_1 _30249_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net189),
    .D(_02577_),
    .Q_N(_11519_),
    .Q(\scanline[107][2] ));
 sg13g2_dfrbp_1 _30250_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net187),
    .D(_02578_),
    .Q_N(_11518_),
    .Q(\scanline[107][3] ));
 sg13g2_dfrbp_1 _30251_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net186),
    .D(_02579_),
    .Q_N(_11517_),
    .Q(\scanline[107][4] ));
 sg13g2_dfrbp_1 _30252_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net185),
    .D(_02580_),
    .Q_N(_11516_),
    .Q(\scanline[107][5] ));
 sg13g2_dfrbp_1 _30253_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net184),
    .D(_02581_),
    .Q_N(_11515_),
    .Q(\scanline[107][6] ));
 sg13g2_dfrbp_1 _30254_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net183),
    .D(_02582_),
    .Q_N(_11514_),
    .Q(\scanline[108][0] ));
 sg13g2_dfrbp_1 _30255_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net182),
    .D(_02583_),
    .Q_N(_11513_),
    .Q(\scanline[108][1] ));
 sg13g2_dfrbp_1 _30256_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net181),
    .D(_02584_),
    .Q_N(_11512_),
    .Q(\scanline[108][2] ));
 sg13g2_dfrbp_1 _30257_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net180),
    .D(_02585_),
    .Q_N(_11511_),
    .Q(\scanline[108][3] ));
 sg13g2_dfrbp_1 _30258_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net179),
    .D(_02586_),
    .Q_N(_11510_),
    .Q(\scanline[108][4] ));
 sg13g2_dfrbp_1 _30259_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net178),
    .D(_02587_),
    .Q_N(_11509_),
    .Q(\scanline[108][5] ));
 sg13g2_dfrbp_1 _30260_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net177),
    .D(_02588_),
    .Q_N(_11508_),
    .Q(\scanline[108][6] ));
 sg13g2_dfrbp_1 _30261_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net176),
    .D(_02589_),
    .Q_N(_11507_),
    .Q(\scanline[10][0] ));
 sg13g2_dfrbp_1 _30262_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net175),
    .D(_02590_),
    .Q_N(_11506_),
    .Q(\scanline[10][1] ));
 sg13g2_dfrbp_1 _30263_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net174),
    .D(_02591_),
    .Q_N(_11505_),
    .Q(\scanline[10][2] ));
 sg13g2_dfrbp_1 _30264_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net173),
    .D(_02592_),
    .Q_N(_11504_),
    .Q(\scanline[10][3] ));
 sg13g2_dfrbp_1 _30265_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net172),
    .D(_02593_),
    .Q_N(_11503_),
    .Q(\scanline[10][4] ));
 sg13g2_dfrbp_1 _30266_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net171),
    .D(_02594_),
    .Q_N(_11502_),
    .Q(\scanline[10][5] ));
 sg13g2_dfrbp_1 _30267_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net170),
    .D(_02595_),
    .Q_N(_11501_),
    .Q(\scanline[10][6] ));
 sg13g2_dfrbp_1 _30268_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net169),
    .D(_02596_),
    .Q_N(_11500_),
    .Q(\scanline[110][0] ));
 sg13g2_dfrbp_1 _30269_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net168),
    .D(_02597_),
    .Q_N(_11499_),
    .Q(\scanline[110][1] ));
 sg13g2_dfrbp_1 _30270_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net167),
    .D(_02598_),
    .Q_N(_11498_),
    .Q(\scanline[110][2] ));
 sg13g2_dfrbp_1 _30271_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net166),
    .D(_02599_),
    .Q_N(_11497_),
    .Q(\scanline[110][3] ));
 sg13g2_dfrbp_1 _30272_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net165),
    .D(_02600_),
    .Q_N(_11496_),
    .Q(\scanline[110][4] ));
 sg13g2_dfrbp_1 _30273_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net164),
    .D(_02601_),
    .Q_N(_11495_),
    .Q(\scanline[110][5] ));
 sg13g2_dfrbp_1 _30274_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net163),
    .D(_02602_),
    .Q_N(_11494_),
    .Q(\scanline[110][6] ));
 sg13g2_dfrbp_1 _30275_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net162),
    .D(_02603_),
    .Q_N(_11493_),
    .Q(\scanline[111][0] ));
 sg13g2_dfrbp_1 _30276_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net161),
    .D(_02604_),
    .Q_N(_11492_),
    .Q(\scanline[111][1] ));
 sg13g2_dfrbp_1 _30277_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net160),
    .D(_02605_),
    .Q_N(_11491_),
    .Q(\scanline[111][2] ));
 sg13g2_dfrbp_1 _30278_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net159),
    .D(_02606_),
    .Q_N(_11490_),
    .Q(\scanline[111][3] ));
 sg13g2_dfrbp_1 _30279_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net158),
    .D(_02607_),
    .Q_N(_11489_),
    .Q(\scanline[111][4] ));
 sg13g2_dfrbp_1 _30280_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net157),
    .D(_02608_),
    .Q_N(_11488_),
    .Q(\scanline[111][5] ));
 sg13g2_dfrbp_1 _30281_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net156),
    .D(_02609_),
    .Q_N(_11487_),
    .Q(\scanline[111][6] ));
 sg13g2_dfrbp_1 _30282_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net155),
    .D(_02610_),
    .Q_N(_11486_),
    .Q(\scanline[112][0] ));
 sg13g2_dfrbp_1 _30283_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net154),
    .D(_02611_),
    .Q_N(_11485_),
    .Q(\scanline[112][1] ));
 sg13g2_dfrbp_1 _30284_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net153),
    .D(_02612_),
    .Q_N(_11484_),
    .Q(\scanline[112][2] ));
 sg13g2_dfrbp_1 _30285_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net152),
    .D(_02613_),
    .Q_N(_11483_),
    .Q(\scanline[112][3] ));
 sg13g2_dfrbp_1 _30286_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net151),
    .D(_02614_),
    .Q_N(_11482_),
    .Q(\scanline[112][4] ));
 sg13g2_dfrbp_1 _30287_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net150),
    .D(_02615_),
    .Q_N(_11481_),
    .Q(\scanline[112][5] ));
 sg13g2_dfrbp_1 _30288_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net149),
    .D(_02616_),
    .Q_N(_11480_),
    .Q(\scanline[112][6] ));
 sg13g2_dfrbp_1 _30289_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net148),
    .D(_02617_),
    .Q_N(_11479_),
    .Q(\scanline[113][0] ));
 sg13g2_dfrbp_1 _30290_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net147),
    .D(_02618_),
    .Q_N(_11478_),
    .Q(\scanline[113][1] ));
 sg13g2_dfrbp_1 _30291_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net146),
    .D(_02619_),
    .Q_N(_11477_),
    .Q(\scanline[113][2] ));
 sg13g2_dfrbp_1 _30292_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net145),
    .D(_02620_),
    .Q_N(_11476_),
    .Q(\scanline[113][3] ));
 sg13g2_dfrbp_1 _30293_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net144),
    .D(_02621_),
    .Q_N(_11475_),
    .Q(\scanline[113][4] ));
 sg13g2_dfrbp_1 _30294_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net143),
    .D(_02622_),
    .Q_N(_11474_),
    .Q(\scanline[113][5] ));
 sg13g2_dfrbp_1 _30295_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net142),
    .D(_02623_),
    .Q_N(_11473_),
    .Q(\scanline[113][6] ));
 sg13g2_dfrbp_1 _30296_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net141),
    .D(_02624_),
    .Q_N(_11472_),
    .Q(\scanline[114][0] ));
 sg13g2_dfrbp_1 _30297_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net140),
    .D(_02625_),
    .Q_N(_11471_),
    .Q(\scanline[114][1] ));
 sg13g2_dfrbp_1 _30298_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net139),
    .D(_02626_),
    .Q_N(_11470_),
    .Q(\scanline[114][2] ));
 sg13g2_dfrbp_1 _30299_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net138),
    .D(_02627_),
    .Q_N(_11469_),
    .Q(\scanline[114][3] ));
 sg13g2_dfrbp_1 _30300_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net137),
    .D(_02628_),
    .Q_N(_11468_),
    .Q(\scanline[114][4] ));
 sg13g2_dfrbp_1 _30301_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net136),
    .D(_02629_),
    .Q_N(_11467_),
    .Q(\scanline[114][5] ));
 sg13g2_dfrbp_1 _30302_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net135),
    .D(_02630_),
    .Q_N(_11466_),
    .Q(\scanline[114][6] ));
 sg13g2_dfrbp_1 _30303_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net134),
    .D(_02631_),
    .Q_N(_11465_),
    .Q(\scanline[115][0] ));
 sg13g2_dfrbp_1 _30304_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net133),
    .D(_02632_),
    .Q_N(_11464_),
    .Q(\scanline[115][1] ));
 sg13g2_dfrbp_1 _30305_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net132),
    .D(_02633_),
    .Q_N(_11463_),
    .Q(\scanline[115][2] ));
 sg13g2_dfrbp_1 _30306_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net131),
    .D(_02634_),
    .Q_N(_11462_),
    .Q(\scanline[115][3] ));
 sg13g2_dfrbp_1 _30307_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net130),
    .D(_02635_),
    .Q_N(_11461_),
    .Q(\scanline[115][4] ));
 sg13g2_dfrbp_1 _30308_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net129),
    .D(_02636_),
    .Q_N(_11460_),
    .Q(\scanline[115][5] ));
 sg13g2_dfrbp_1 _30309_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net128),
    .D(_02637_),
    .Q_N(_11459_),
    .Q(\scanline[115][6] ));
 sg13g2_dfrbp_1 _30310_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net127),
    .D(_02638_),
    .Q_N(_11458_),
    .Q(\scanline[116][0] ));
 sg13g2_dfrbp_1 _30311_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net126),
    .D(_02639_),
    .Q_N(_11457_),
    .Q(\scanline[116][1] ));
 sg13g2_dfrbp_1 _30312_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net125),
    .D(_02640_),
    .Q_N(_11456_),
    .Q(\scanline[116][2] ));
 sg13g2_dfrbp_1 _30313_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net124),
    .D(_02641_),
    .Q_N(_11455_),
    .Q(\scanline[116][3] ));
 sg13g2_dfrbp_1 _30314_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net123),
    .D(_02642_),
    .Q_N(_11454_),
    .Q(\scanline[116][4] ));
 sg13g2_dfrbp_1 _30315_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net122),
    .D(_02643_),
    .Q_N(_11453_),
    .Q(\scanline[116][5] ));
 sg13g2_dfrbp_1 _30316_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net121),
    .D(_02644_),
    .Q_N(_11452_),
    .Q(\scanline[116][6] ));
 sg13g2_dfrbp_1 _30317_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net120),
    .D(_02645_),
    .Q_N(_11451_),
    .Q(\scanline[117][0] ));
 sg13g2_dfrbp_1 _30318_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net119),
    .D(_02646_),
    .Q_N(_11450_),
    .Q(\scanline[117][1] ));
 sg13g2_dfrbp_1 _30319_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net118),
    .D(_02647_),
    .Q_N(_11449_),
    .Q(\scanline[117][2] ));
 sg13g2_dfrbp_1 _30320_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net117),
    .D(_02648_),
    .Q_N(_11448_),
    .Q(\scanline[117][3] ));
 sg13g2_dfrbp_1 _30321_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net116),
    .D(_02649_),
    .Q_N(_11447_),
    .Q(\scanline[117][4] ));
 sg13g2_dfrbp_1 _30322_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net115),
    .D(_02650_),
    .Q_N(_11446_),
    .Q(\scanline[117][5] ));
 sg13g2_dfrbp_1 _30323_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net114),
    .D(_02651_),
    .Q_N(_11445_),
    .Q(\scanline[117][6] ));
 sg13g2_dfrbp_1 _30324_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net113),
    .D(_02652_),
    .Q_N(_11444_),
    .Q(\scanline[118][0] ));
 sg13g2_dfrbp_1 _30325_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net112),
    .D(_02653_),
    .Q_N(_11443_),
    .Q(\scanline[118][1] ));
 sg13g2_dfrbp_1 _30326_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net111),
    .D(_02654_),
    .Q_N(_11442_),
    .Q(\scanline[118][2] ));
 sg13g2_dfrbp_1 _30327_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net110),
    .D(_02655_),
    .Q_N(_11441_),
    .Q(\scanline[118][3] ));
 sg13g2_dfrbp_1 _30328_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net109),
    .D(_02656_),
    .Q_N(_11440_),
    .Q(\scanline[118][4] ));
 sg13g2_dfrbp_1 _30329_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net108),
    .D(_02657_),
    .Q_N(_11439_),
    .Q(\scanline[118][5] ));
 sg13g2_dfrbp_1 _30330_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net107),
    .D(_02658_),
    .Q_N(_11438_),
    .Q(\scanline[118][6] ));
 sg13g2_dfrbp_1 _30331_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net106),
    .D(_02659_),
    .Q_N(_11437_),
    .Q(\scanline[11][0] ));
 sg13g2_dfrbp_1 _30332_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net105),
    .D(_02660_),
    .Q_N(_11436_),
    .Q(\scanline[11][1] ));
 sg13g2_dfrbp_1 _30333_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net104),
    .D(_02661_),
    .Q_N(_11435_),
    .Q(\scanline[11][2] ));
 sg13g2_dfrbp_1 _30334_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net103),
    .D(_02662_),
    .Q_N(_11434_),
    .Q(\scanline[11][3] ));
 sg13g2_dfrbp_1 _30335_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net102),
    .D(_02663_),
    .Q_N(_11433_),
    .Q(\scanline[11][4] ));
 sg13g2_dfrbp_1 _30336_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net101),
    .D(_02664_),
    .Q_N(_11432_),
    .Q(\scanline[11][5] ));
 sg13g2_dfrbp_1 _30337_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net100),
    .D(_02665_),
    .Q_N(_11431_),
    .Q(\scanline[11][6] ));
 sg13g2_dfrbp_1 _30338_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net97),
    .D(_02666_),
    .Q_N(_11430_),
    .Q(\scanline[120][0] ));
 sg13g2_dfrbp_1 _30339_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net96),
    .D(_02667_),
    .Q_N(_11429_),
    .Q(\scanline[120][1] ));
 sg13g2_dfrbp_1 _30340_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net95),
    .D(_02668_),
    .Q_N(_11428_),
    .Q(\scanline[120][2] ));
 sg13g2_dfrbp_1 _30341_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net94),
    .D(_02669_),
    .Q_N(_11427_),
    .Q(\scanline[120][3] ));
 sg13g2_dfrbp_1 _30342_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net93),
    .D(_02670_),
    .Q_N(_11426_),
    .Q(\scanline[120][4] ));
 sg13g2_dfrbp_1 _30343_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net92),
    .D(_02671_),
    .Q_N(_11425_),
    .Q(\scanline[120][5] ));
 sg13g2_dfrbp_1 _30344_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net91),
    .D(_02672_),
    .Q_N(_11424_),
    .Q(\scanline[120][6] ));
 sg13g2_dfrbp_1 _30345_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net90),
    .D(_02673_),
    .Q_N(_11423_),
    .Q(\scanline[121][0] ));
 sg13g2_dfrbp_1 _30346_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net89),
    .D(_02674_),
    .Q_N(_11422_),
    .Q(\scanline[121][1] ));
 sg13g2_dfrbp_1 _30347_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net88),
    .D(_02675_),
    .Q_N(_11421_),
    .Q(\scanline[121][2] ));
 sg13g2_dfrbp_1 _30348_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net87),
    .D(_02676_),
    .Q_N(_11420_),
    .Q(\scanline[121][3] ));
 sg13g2_dfrbp_1 _30349_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net86),
    .D(_02677_),
    .Q_N(_11419_),
    .Q(\scanline[121][4] ));
 sg13g2_dfrbp_1 _30350_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net85),
    .D(_02678_),
    .Q_N(_11418_),
    .Q(\scanline[121][5] ));
 sg13g2_dfrbp_1 _30351_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net84),
    .D(_02679_),
    .Q_N(_11417_),
    .Q(\scanline[121][6] ));
 sg13g2_dfrbp_1 _30352_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net83),
    .D(_02680_),
    .Q_N(_11416_),
    .Q(\scanline[122][0] ));
 sg13g2_dfrbp_1 _30353_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net82),
    .D(_02681_),
    .Q_N(_11415_),
    .Q(\scanline[122][1] ));
 sg13g2_dfrbp_1 _30354_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net81),
    .D(_02682_),
    .Q_N(_11414_),
    .Q(\scanline[122][2] ));
 sg13g2_dfrbp_1 _30355_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net80),
    .D(_02683_),
    .Q_N(_11413_),
    .Q(\scanline[122][3] ));
 sg13g2_dfrbp_1 _30356_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net79),
    .D(_02684_),
    .Q_N(_11412_),
    .Q(\scanline[122][4] ));
 sg13g2_dfrbp_1 _30357_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net78),
    .D(_02685_),
    .Q_N(_11411_),
    .Q(\scanline[122][5] ));
 sg13g2_dfrbp_1 _30358_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net77),
    .D(_02686_),
    .Q_N(_11410_),
    .Q(\scanline[122][6] ));
 sg13g2_dfrbp_1 _30359_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net76),
    .D(_02687_),
    .Q_N(_11409_),
    .Q(\scanline[123][0] ));
 sg13g2_dfrbp_1 _30360_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net75),
    .D(_02688_),
    .Q_N(_11408_),
    .Q(\scanline[123][1] ));
 sg13g2_dfrbp_1 _30361_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net74),
    .D(_02689_),
    .Q_N(_11407_),
    .Q(\scanline[123][2] ));
 sg13g2_dfrbp_1 _30362_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net73),
    .D(_02690_),
    .Q_N(_11406_),
    .Q(\scanline[123][3] ));
 sg13g2_dfrbp_1 _30363_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net72),
    .D(_02691_),
    .Q_N(_11405_),
    .Q(\scanline[123][4] ));
 sg13g2_dfrbp_1 _30364_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net71),
    .D(_02692_),
    .Q_N(_11404_),
    .Q(\scanline[123][5] ));
 sg13g2_dfrbp_1 _30365_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net70),
    .D(_02693_),
    .Q_N(_11403_),
    .Q(\scanline[123][6] ));
 sg13g2_dfrbp_1 _30366_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net69),
    .D(_02694_),
    .Q_N(_11402_),
    .Q(\scanline[124][0] ));
 sg13g2_dfrbp_1 _30367_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net68),
    .D(_02695_),
    .Q_N(_11401_),
    .Q(\scanline[124][1] ));
 sg13g2_dfrbp_1 _30368_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net67),
    .D(_02696_),
    .Q_N(_11400_),
    .Q(\scanline[124][2] ));
 sg13g2_dfrbp_1 _30369_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net66),
    .D(_02697_),
    .Q_N(_11399_),
    .Q(\scanline[124][3] ));
 sg13g2_dfrbp_1 _30370_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net65),
    .D(_02698_),
    .Q_N(_11398_),
    .Q(\scanline[124][4] ));
 sg13g2_dfrbp_1 _30371_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net64),
    .D(_02699_),
    .Q_N(_11397_),
    .Q(\scanline[124][5] ));
 sg13g2_dfrbp_1 _30372_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net63),
    .D(_02700_),
    .Q_N(_11396_),
    .Q(\scanline[124][6] ));
 sg13g2_dfrbp_1 _30373_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net62),
    .D(_02701_),
    .Q_N(_11395_),
    .Q(\scanline[125][0] ));
 sg13g2_dfrbp_1 _30374_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net61),
    .D(_02702_),
    .Q_N(_11394_),
    .Q(\scanline[125][1] ));
 sg13g2_dfrbp_1 _30375_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net60),
    .D(_02703_),
    .Q_N(_11393_),
    .Q(\scanline[125][2] ));
 sg13g2_dfrbp_1 _30376_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net59),
    .D(_02704_),
    .Q_N(_11392_),
    .Q(\scanline[125][3] ));
 sg13g2_dfrbp_1 _30377_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net58),
    .D(_02705_),
    .Q_N(_11391_),
    .Q(\scanline[125][4] ));
 sg13g2_dfrbp_1 _30378_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net57),
    .D(_02706_),
    .Q_N(_11390_),
    .Q(\scanline[125][5] ));
 sg13g2_dfrbp_1 _30379_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net56),
    .D(_02707_),
    .Q_N(_11389_),
    .Q(\scanline[125][6] ));
 sg13g2_dfrbp_1 _30380_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net55),
    .D(_02708_),
    .Q_N(_11388_),
    .Q(\scanline[126][0] ));
 sg13g2_dfrbp_1 _30381_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net54),
    .D(_02709_),
    .Q_N(_11387_),
    .Q(\scanline[126][1] ));
 sg13g2_dfrbp_1 _30382_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net53),
    .D(_02710_),
    .Q_N(_11386_),
    .Q(\scanline[126][2] ));
 sg13g2_dfrbp_1 _30383_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net52),
    .D(_02711_),
    .Q_N(_11385_),
    .Q(\scanline[126][3] ));
 sg13g2_dfrbp_1 _30384_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net51),
    .D(_02712_),
    .Q_N(_11384_),
    .Q(\scanline[126][4] ));
 sg13g2_dfrbp_1 _30385_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net50),
    .D(_02713_),
    .Q_N(_11383_),
    .Q(\scanline[126][5] ));
 sg13g2_dfrbp_1 _30386_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net49),
    .D(_02714_),
    .Q_N(_11382_),
    .Q(\scanline[126][6] ));
 sg13g2_dfrbp_1 _30387_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net48),
    .D(_02715_),
    .Q_N(_11381_),
    .Q(\scanline[127][0] ));
 sg13g2_dfrbp_1 _30388_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net47),
    .D(_02716_),
    .Q_N(_11380_),
    .Q(\scanline[127][1] ));
 sg13g2_dfrbp_1 _30389_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net46),
    .D(_02717_),
    .Q_N(_11379_),
    .Q(\scanline[127][2] ));
 sg13g2_dfrbp_1 _30390_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net45),
    .D(_02718_),
    .Q_N(_11378_),
    .Q(\scanline[127][3] ));
 sg13g2_dfrbp_1 _30391_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net44),
    .D(_02719_),
    .Q_N(_11377_),
    .Q(\scanline[127][4] ));
 sg13g2_dfrbp_1 _30392_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net43),
    .D(_02720_),
    .Q_N(_11376_),
    .Q(\scanline[127][5] ));
 sg13g2_dfrbp_1 _30393_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net42),
    .D(_02721_),
    .Q_N(_11375_),
    .Q(\scanline[127][6] ));
 sg13g2_dfrbp_1 _30394_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net41),
    .D(_02722_),
    .Q_N(_11374_),
    .Q(\scanline[128][0] ));
 sg13g2_dfrbp_1 _30395_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net40),
    .D(_02723_),
    .Q_N(_11373_),
    .Q(\scanline[128][1] ));
 sg13g2_dfrbp_1 _30396_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net39),
    .D(_02724_),
    .Q_N(_11372_),
    .Q(\scanline[128][2] ));
 sg13g2_dfrbp_1 _30397_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net38),
    .D(_02725_),
    .Q_N(_11371_),
    .Q(\scanline[128][3] ));
 sg13g2_dfrbp_1 _30398_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net37),
    .D(_02726_),
    .Q_N(_11370_),
    .Q(\scanline[128][4] ));
 sg13g2_dfrbp_1 _30399_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net36),
    .D(_02727_),
    .Q_N(_11369_),
    .Q(\scanline[128][5] ));
 sg13g2_dfrbp_1 _30400_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net35),
    .D(_02728_),
    .Q_N(_11368_),
    .Q(\scanline[128][6] ));
 sg13g2_dfrbp_1 _30401_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net34),
    .D(_02729_),
    .Q_N(_11367_),
    .Q(\scanline[12][0] ));
 sg13g2_dfrbp_1 _30402_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net33),
    .D(_02730_),
    .Q_N(_11366_),
    .Q(\scanline[12][1] ));
 sg13g2_dfrbp_1 _30403_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net32),
    .D(_02731_),
    .Q_N(_11365_),
    .Q(\scanline[12][2] ));
 sg13g2_dfrbp_1 _30404_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net31),
    .D(_02732_),
    .Q_N(_11364_),
    .Q(\scanline[12][3] ));
 sg13g2_dfrbp_1 _30405_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net30),
    .D(_02733_),
    .Q_N(_11363_),
    .Q(\scanline[12][4] ));
 sg13g2_dfrbp_1 _30406_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net29),
    .D(_02734_),
    .Q_N(_11362_),
    .Q(\scanline[12][5] ));
 sg13g2_dfrbp_1 _30407_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net28),
    .D(_02735_),
    .Q_N(_11361_),
    .Q(\scanline[12][6] ));
 sg13g2_dfrbp_1 _30408_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net27),
    .D(_02736_),
    .Q_N(_11360_),
    .Q(\scanline[130][0] ));
 sg13g2_dfrbp_1 _30409_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net26),
    .D(_02737_),
    .Q_N(_11359_),
    .Q(\scanline[130][1] ));
 sg13g2_dfrbp_1 _30410_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net25),
    .D(_02738_),
    .Q_N(_11358_),
    .Q(\scanline[130][2] ));
 sg13g2_dfrbp_1 _30411_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net24),
    .D(_02739_),
    .Q_N(_11357_),
    .Q(\scanline[130][3] ));
 sg13g2_dfrbp_1 _30412_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net23),
    .D(_02740_),
    .Q_N(_11356_),
    .Q(\scanline[130][4] ));
 sg13g2_dfrbp_1 _30413_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net22),
    .D(_02741_),
    .Q_N(_11355_),
    .Q(\scanline[130][5] ));
 sg13g2_dfrbp_1 _30414_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net21),
    .D(_02742_),
    .Q_N(_11354_),
    .Q(\scanline[130][6] ));
 sg13g2_dfrbp_1 _30415_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net20),
    .D(_02743_),
    .Q_N(_11353_),
    .Q(\scanline[131][0] ));
 sg13g2_dfrbp_1 _30416_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net19),
    .D(_02744_),
    .Q_N(_11352_),
    .Q(\scanline[131][1] ));
 sg13g2_dfrbp_1 _30417_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net18),
    .D(_02745_),
    .Q_N(_11351_),
    .Q(\scanline[131][2] ));
 sg13g2_dfrbp_1 _30418_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net17),
    .D(_02746_),
    .Q_N(_11350_),
    .Q(\scanline[131][3] ));
 sg13g2_dfrbp_1 _30419_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net16),
    .D(_02747_),
    .Q_N(_11349_),
    .Q(\scanline[131][4] ));
 sg13g2_dfrbp_1 _30420_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net15),
    .D(_02748_),
    .Q_N(_11348_),
    .Q(\scanline[131][5] ));
 sg13g2_dfrbp_1 _30421_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net14),
    .D(_02749_),
    .Q_N(_11347_),
    .Q(\scanline[131][6] ));
 sg13g2_dfrbp_1 _30422_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net13),
    .D(_02750_),
    .Q_N(_11346_),
    .Q(\scanline[132][0] ));
 sg13g2_dfrbp_1 _30423_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2922),
    .D(_02751_),
    .Q_N(_11345_),
    .Q(\scanline[132][1] ));
 sg13g2_dfrbp_1 _30424_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2921),
    .D(_02752_),
    .Q_N(_11344_),
    .Q(\scanline[132][2] ));
 sg13g2_dfrbp_1 _30425_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2920),
    .D(_02753_),
    .Q_N(_11343_),
    .Q(\scanline[132][3] ));
 sg13g2_dfrbp_1 _30426_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2919),
    .D(_02754_),
    .Q_N(_11342_),
    .Q(\scanline[132][4] ));
 sg13g2_dfrbp_1 _30427_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2918),
    .D(_02755_),
    .Q_N(_11341_),
    .Q(\scanline[132][5] ));
 sg13g2_dfrbp_1 _30428_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2917),
    .D(_02756_),
    .Q_N(_11340_),
    .Q(\scanline[132][6] ));
 sg13g2_dfrbp_1 _30429_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2916),
    .D(_02757_),
    .Q_N(_11339_),
    .Q(\scanline[133][0] ));
 sg13g2_dfrbp_1 _30430_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2915),
    .D(_02758_),
    .Q_N(_11338_),
    .Q(\scanline[133][1] ));
 sg13g2_dfrbp_1 _30431_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2914),
    .D(_02759_),
    .Q_N(_11337_),
    .Q(\scanline[133][2] ));
 sg13g2_dfrbp_1 _30432_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2913),
    .D(_02760_),
    .Q_N(_11336_),
    .Q(\scanline[133][3] ));
 sg13g2_dfrbp_1 _30433_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2912),
    .D(_02761_),
    .Q_N(_11335_),
    .Q(\scanline[133][4] ));
 sg13g2_dfrbp_1 _30434_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2911),
    .D(_02762_),
    .Q_N(_11334_),
    .Q(\scanline[133][5] ));
 sg13g2_dfrbp_1 _30435_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2910),
    .D(_02763_),
    .Q_N(_11333_),
    .Q(\scanline[133][6] ));
 sg13g2_dfrbp_1 _30436_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2909),
    .D(_02764_),
    .Q_N(_11332_),
    .Q(\scanline[134][0] ));
 sg13g2_dfrbp_1 _30437_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2908),
    .D(_02765_),
    .Q_N(_11331_),
    .Q(\scanline[134][1] ));
 sg13g2_dfrbp_1 _30438_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2907),
    .D(_02766_),
    .Q_N(_11330_),
    .Q(\scanline[134][2] ));
 sg13g2_dfrbp_1 _30439_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2906),
    .D(_02767_),
    .Q_N(_11329_),
    .Q(\scanline[134][3] ));
 sg13g2_dfrbp_1 _30440_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2905),
    .D(_02768_),
    .Q_N(_11328_),
    .Q(\scanline[134][4] ));
 sg13g2_dfrbp_1 _30441_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2904),
    .D(_02769_),
    .Q_N(_11327_),
    .Q(\scanline[134][5] ));
 sg13g2_dfrbp_1 _30442_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2903),
    .D(_02770_),
    .Q_N(_11326_),
    .Q(\scanline[134][6] ));
 sg13g2_dfrbp_1 _30443_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2902),
    .D(_02771_),
    .Q_N(_11325_),
    .Q(\scanline[135][0] ));
 sg13g2_dfrbp_1 _30444_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2901),
    .D(_02772_),
    .Q_N(_11324_),
    .Q(\scanline[135][1] ));
 sg13g2_dfrbp_1 _30445_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2900),
    .D(_02773_),
    .Q_N(_11323_),
    .Q(\scanline[135][2] ));
 sg13g2_dfrbp_1 _30446_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2899),
    .D(_02774_),
    .Q_N(_11322_),
    .Q(\scanline[135][3] ));
 sg13g2_dfrbp_1 _30447_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2898),
    .D(_02775_),
    .Q_N(_11321_),
    .Q(\scanline[135][4] ));
 sg13g2_dfrbp_1 _30448_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2897),
    .D(_02776_),
    .Q_N(_11320_),
    .Q(\scanline[135][5] ));
 sg13g2_dfrbp_1 _30449_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2896),
    .D(_02777_),
    .Q_N(_11319_),
    .Q(\scanline[135][6] ));
 sg13g2_dfrbp_1 _30450_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2895),
    .D(_02778_),
    .Q_N(_11318_),
    .Q(\scanline[136][0] ));
 sg13g2_dfrbp_1 _30451_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net2894),
    .D(_02779_),
    .Q_N(_11317_),
    .Q(\scanline[136][1] ));
 sg13g2_dfrbp_1 _30452_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2893),
    .D(_02780_),
    .Q_N(_11316_),
    .Q(\scanline[136][2] ));
 sg13g2_dfrbp_1 _30453_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2892),
    .D(_02781_),
    .Q_N(_11315_),
    .Q(\scanline[136][3] ));
 sg13g2_dfrbp_1 _30454_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2891),
    .D(_02782_),
    .Q_N(_11314_),
    .Q(\scanline[136][4] ));
 sg13g2_dfrbp_1 _30455_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2890),
    .D(_02783_),
    .Q_N(_11313_),
    .Q(\scanline[136][5] ));
 sg13g2_dfrbp_1 _30456_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2889),
    .D(_02784_),
    .Q_N(_11312_),
    .Q(\scanline[136][6] ));
 sg13g2_dfrbp_1 _30457_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2888),
    .D(_02785_),
    .Q_N(_11311_),
    .Q(\scanline[137][0] ));
 sg13g2_dfrbp_1 _30458_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2887),
    .D(_02786_),
    .Q_N(_11310_),
    .Q(\scanline[137][1] ));
 sg13g2_dfrbp_1 _30459_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2886),
    .D(_02787_),
    .Q_N(_11309_),
    .Q(\scanline[137][2] ));
 sg13g2_dfrbp_1 _30460_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2885),
    .D(_02788_),
    .Q_N(_11308_),
    .Q(\scanline[137][3] ));
 sg13g2_dfrbp_1 _30461_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2884),
    .D(_02789_),
    .Q_N(_11307_),
    .Q(\scanline[137][4] ));
 sg13g2_dfrbp_1 _30462_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2883),
    .D(_02790_),
    .Q_N(_11306_),
    .Q(\scanline[137][5] ));
 sg13g2_dfrbp_1 _30463_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2882),
    .D(_02791_),
    .Q_N(_11305_),
    .Q(\scanline[137][6] ));
 sg13g2_dfrbp_1 _30464_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2881),
    .D(_02792_),
    .Q_N(_11304_),
    .Q(\scanline[138][0] ));
 sg13g2_dfrbp_1 _30465_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net2880),
    .D(_02793_),
    .Q_N(_11303_),
    .Q(\scanline[138][1] ));
 sg13g2_dfrbp_1 _30466_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2879),
    .D(_02794_),
    .Q_N(_11302_),
    .Q(\scanline[138][2] ));
 sg13g2_dfrbp_1 _30467_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2878),
    .D(_02795_),
    .Q_N(_11301_),
    .Q(\scanline[138][3] ));
 sg13g2_dfrbp_1 _30468_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2877),
    .D(_02796_),
    .Q_N(_11300_),
    .Q(\scanline[138][4] ));
 sg13g2_dfrbp_1 _30469_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2876),
    .D(_02797_),
    .Q_N(_11299_),
    .Q(\scanline[138][5] ));
 sg13g2_dfrbp_1 _30470_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2875),
    .D(_02798_),
    .Q_N(_11298_),
    .Q(\scanline[138][6] ));
 sg13g2_dfrbp_1 _30471_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2874),
    .D(_02799_),
    .Q_N(_11297_),
    .Q(\scanline[13][0] ));
 sg13g2_dfrbp_1 _30472_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2873),
    .D(_02800_),
    .Q_N(_11296_),
    .Q(\scanline[13][1] ));
 sg13g2_dfrbp_1 _30473_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2872),
    .D(_02801_),
    .Q_N(_11295_),
    .Q(\scanline[13][2] ));
 sg13g2_dfrbp_1 _30474_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2871),
    .D(_02802_),
    .Q_N(_11294_),
    .Q(\scanline[13][3] ));
 sg13g2_dfrbp_1 _30475_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2870),
    .D(_02803_),
    .Q_N(_11293_),
    .Q(\scanline[13][4] ));
 sg13g2_dfrbp_1 _30476_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2869),
    .D(_02804_),
    .Q_N(_11292_),
    .Q(\scanline[13][5] ));
 sg13g2_dfrbp_1 _30477_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2868),
    .D(_02805_),
    .Q_N(_11291_),
    .Q(\scanline[13][6] ));
 sg13g2_dfrbp_1 _30478_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2867),
    .D(_02806_),
    .Q_N(_11290_),
    .Q(\scanline[140][0] ));
 sg13g2_dfrbp_1 _30479_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2866),
    .D(_02807_),
    .Q_N(_11289_),
    .Q(\scanline[140][1] ));
 sg13g2_dfrbp_1 _30480_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2865),
    .D(_02808_),
    .Q_N(_11288_),
    .Q(\scanline[140][2] ));
 sg13g2_dfrbp_1 _30481_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2864),
    .D(_02809_),
    .Q_N(_11287_),
    .Q(\scanline[140][3] ));
 sg13g2_dfrbp_1 _30482_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2863),
    .D(_02810_),
    .Q_N(_11286_),
    .Q(\scanline[140][4] ));
 sg13g2_dfrbp_1 _30483_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2862),
    .D(_02811_),
    .Q_N(_11285_),
    .Q(\scanline[140][5] ));
 sg13g2_dfrbp_1 _30484_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2861),
    .D(_02812_),
    .Q_N(_11284_),
    .Q(\scanline[140][6] ));
 sg13g2_dfrbp_1 _30485_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2860),
    .D(_02813_),
    .Q_N(_11283_),
    .Q(\scanline[141][0] ));
 sg13g2_dfrbp_1 _30486_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2859),
    .D(_02814_),
    .Q_N(_11282_),
    .Q(\scanline[141][1] ));
 sg13g2_dfrbp_1 _30487_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2858),
    .D(_02815_),
    .Q_N(_11281_),
    .Q(\scanline[141][2] ));
 sg13g2_dfrbp_1 _30488_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2857),
    .D(_02816_),
    .Q_N(_11280_),
    .Q(\scanline[141][3] ));
 sg13g2_dfrbp_1 _30489_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2856),
    .D(_02817_),
    .Q_N(_11279_),
    .Q(\scanline[141][4] ));
 sg13g2_dfrbp_1 _30490_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2855),
    .D(_02818_),
    .Q_N(_11278_),
    .Q(\scanline[141][5] ));
 sg13g2_dfrbp_1 _30491_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2854),
    .D(_02819_),
    .Q_N(_11277_),
    .Q(\scanline[141][6] ));
 sg13g2_dfrbp_1 _30492_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2853),
    .D(_02820_),
    .Q_N(_11276_),
    .Q(\scanline[142][0] ));
 sg13g2_dfrbp_1 _30493_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2852),
    .D(_02821_),
    .Q_N(_11275_),
    .Q(\scanline[142][1] ));
 sg13g2_dfrbp_1 _30494_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2851),
    .D(_02822_),
    .Q_N(_11274_),
    .Q(\scanline[142][2] ));
 sg13g2_dfrbp_1 _30495_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2850),
    .D(_02823_),
    .Q_N(_11273_),
    .Q(\scanline[142][3] ));
 sg13g2_dfrbp_1 _30496_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2849),
    .D(_02824_),
    .Q_N(_11272_),
    .Q(\scanline[142][4] ));
 sg13g2_dfrbp_1 _30497_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2848),
    .D(_02825_),
    .Q_N(_11271_),
    .Q(\scanline[142][5] ));
 sg13g2_dfrbp_1 _30498_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2847),
    .D(_02826_),
    .Q_N(_11270_),
    .Q(\scanline[142][6] ));
 sg13g2_dfrbp_1 _30499_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2846),
    .D(_02827_),
    .Q_N(_11269_),
    .Q(\scanline[143][0] ));
 sg13g2_dfrbp_1 _30500_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2845),
    .D(_02828_),
    .Q_N(_11268_),
    .Q(\scanline[143][1] ));
 sg13g2_dfrbp_1 _30501_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2844),
    .D(_02829_),
    .Q_N(_11267_),
    .Q(\scanline[143][2] ));
 sg13g2_dfrbp_1 _30502_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2843),
    .D(_02830_),
    .Q_N(_11266_),
    .Q(\scanline[143][3] ));
 sg13g2_dfrbp_1 _30503_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2842),
    .D(_02831_),
    .Q_N(_11265_),
    .Q(\scanline[143][4] ));
 sg13g2_dfrbp_1 _30504_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2841),
    .D(_02832_),
    .Q_N(_11264_),
    .Q(\scanline[143][5] ));
 sg13g2_dfrbp_1 _30505_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2840),
    .D(_02833_),
    .Q_N(_11263_),
    .Q(\scanline[143][6] ));
 sg13g2_dfrbp_1 _30506_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2839),
    .D(_02834_),
    .Q_N(_11262_),
    .Q(\scanline[144][0] ));
 sg13g2_dfrbp_1 _30507_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2838),
    .D(_02835_),
    .Q_N(_11261_),
    .Q(\scanline[144][1] ));
 sg13g2_dfrbp_1 _30508_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2837),
    .D(_02836_),
    .Q_N(_11260_),
    .Q(\scanline[144][2] ));
 sg13g2_dfrbp_1 _30509_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2836),
    .D(_02837_),
    .Q_N(_11259_),
    .Q(\scanline[144][3] ));
 sg13g2_dfrbp_1 _30510_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2835),
    .D(_02838_),
    .Q_N(_11258_),
    .Q(\scanline[144][4] ));
 sg13g2_dfrbp_1 _30511_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2834),
    .D(_02839_),
    .Q_N(_11257_),
    .Q(\scanline[144][5] ));
 sg13g2_dfrbp_1 _30512_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2833),
    .D(_02840_),
    .Q_N(_11256_),
    .Q(\scanline[144][6] ));
 sg13g2_dfrbp_1 _30513_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2832),
    .D(_02841_),
    .Q_N(_11255_),
    .Q(\scanline[145][0] ));
 sg13g2_dfrbp_1 _30514_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2831),
    .D(_02842_),
    .Q_N(_11254_),
    .Q(\scanline[145][1] ));
 sg13g2_dfrbp_1 _30515_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2830),
    .D(_02843_),
    .Q_N(_11253_),
    .Q(\scanline[145][2] ));
 sg13g2_dfrbp_1 _30516_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2829),
    .D(_02844_),
    .Q_N(_11252_),
    .Q(\scanline[145][3] ));
 sg13g2_dfrbp_1 _30517_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2828),
    .D(_02845_),
    .Q_N(_11251_),
    .Q(\scanline[145][4] ));
 sg13g2_dfrbp_1 _30518_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2827),
    .D(_02846_),
    .Q_N(_11250_),
    .Q(\scanline[145][5] ));
 sg13g2_dfrbp_1 _30519_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2826),
    .D(_02847_),
    .Q_N(_11249_),
    .Q(\scanline[145][6] ));
 sg13g2_dfrbp_1 _30520_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2825),
    .D(_02848_),
    .Q_N(_11248_),
    .Q(\scanline[146][0] ));
 sg13g2_dfrbp_1 _30521_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2824),
    .D(_02849_),
    .Q_N(_11247_),
    .Q(\scanline[146][1] ));
 sg13g2_dfrbp_1 _30522_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2823),
    .D(_02850_),
    .Q_N(_11246_),
    .Q(\scanline[146][2] ));
 sg13g2_dfrbp_1 _30523_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2822),
    .D(_02851_),
    .Q_N(_11245_),
    .Q(\scanline[146][3] ));
 sg13g2_dfrbp_1 _30524_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2821),
    .D(_02852_),
    .Q_N(_11244_),
    .Q(\scanline[146][4] ));
 sg13g2_dfrbp_1 _30525_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2820),
    .D(_02853_),
    .Q_N(_11243_),
    .Q(\scanline[146][5] ));
 sg13g2_dfrbp_1 _30526_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2819),
    .D(_02854_),
    .Q_N(_11242_),
    .Q(\scanline[146][6] ));
 sg13g2_dfrbp_1 _30527_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2818),
    .D(_02855_),
    .Q_N(_11241_),
    .Q(\scanline[147][0] ));
 sg13g2_dfrbp_1 _30528_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2817),
    .D(_02856_),
    .Q_N(_11240_),
    .Q(\scanline[147][1] ));
 sg13g2_dfrbp_1 _30529_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2816),
    .D(_02857_),
    .Q_N(_11239_),
    .Q(\scanline[147][2] ));
 sg13g2_dfrbp_1 _30530_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2815),
    .D(_02858_),
    .Q_N(_11238_),
    .Q(\scanline[147][3] ));
 sg13g2_dfrbp_1 _30531_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2814),
    .D(_02859_),
    .Q_N(_11237_),
    .Q(\scanline[147][4] ));
 sg13g2_dfrbp_1 _30532_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2813),
    .D(_02860_),
    .Q_N(_11236_),
    .Q(\scanline[147][5] ));
 sg13g2_dfrbp_1 _30533_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2812),
    .D(_02861_),
    .Q_N(_11235_),
    .Q(\scanline[147][6] ));
 sg13g2_dfrbp_1 _30534_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2811),
    .D(_02862_),
    .Q_N(_11234_),
    .Q(\scanline[148][0] ));
 sg13g2_dfrbp_1 _30535_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2810),
    .D(_02863_),
    .Q_N(_11233_),
    .Q(\scanline[148][1] ));
 sg13g2_dfrbp_1 _30536_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2809),
    .D(_02864_),
    .Q_N(_11232_),
    .Q(\scanline[148][2] ));
 sg13g2_dfrbp_1 _30537_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2808),
    .D(_02865_),
    .Q_N(_11231_),
    .Q(\scanline[148][3] ));
 sg13g2_dfrbp_1 _30538_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2807),
    .D(_02866_),
    .Q_N(_11230_),
    .Q(\scanline[148][4] ));
 sg13g2_dfrbp_1 _30539_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2806),
    .D(_02867_),
    .Q_N(_11229_),
    .Q(\scanline[148][5] ));
 sg13g2_dfrbp_1 _30540_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2805),
    .D(_02868_),
    .Q_N(_11228_),
    .Q(\scanline[148][6] ));
 sg13g2_dfrbp_1 _30541_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2804),
    .D(_02869_),
    .Q_N(_11227_),
    .Q(\scanline[14][0] ));
 sg13g2_dfrbp_1 _30542_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2803),
    .D(_02870_),
    .Q_N(_11226_),
    .Q(\scanline[14][1] ));
 sg13g2_dfrbp_1 _30543_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2802),
    .D(_02871_),
    .Q_N(_11225_),
    .Q(\scanline[14][2] ));
 sg13g2_dfrbp_1 _30544_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2801),
    .D(_02872_),
    .Q_N(_11224_),
    .Q(\scanline[14][3] ));
 sg13g2_dfrbp_1 _30545_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2800),
    .D(_02873_),
    .Q_N(_11223_),
    .Q(\scanline[14][4] ));
 sg13g2_dfrbp_1 _30546_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2799),
    .D(_02874_),
    .Q_N(_11222_),
    .Q(\scanline[14][5] ));
 sg13g2_dfrbp_1 _30547_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2798),
    .D(_02875_),
    .Q_N(_11221_),
    .Q(\scanline[14][6] ));
 sg13g2_dfrbp_1 _30548_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2797),
    .D(_02876_),
    .Q_N(_11220_),
    .Q(\scanline[150][0] ));
 sg13g2_dfrbp_1 _30549_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2796),
    .D(_02877_),
    .Q_N(_11219_),
    .Q(\scanline[150][1] ));
 sg13g2_dfrbp_1 _30550_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2795),
    .D(_02878_),
    .Q_N(_11218_),
    .Q(\scanline[150][2] ));
 sg13g2_dfrbp_1 _30551_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2794),
    .D(_02879_),
    .Q_N(_11217_),
    .Q(\scanline[150][3] ));
 sg13g2_dfrbp_1 _30552_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2793),
    .D(_02880_),
    .Q_N(_11216_),
    .Q(\scanline[150][4] ));
 sg13g2_dfrbp_1 _30553_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2792),
    .D(_02881_),
    .Q_N(_11215_),
    .Q(\scanline[150][5] ));
 sg13g2_dfrbp_1 _30554_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2791),
    .D(_02882_),
    .Q_N(_11214_),
    .Q(\scanline[150][6] ));
 sg13g2_dfrbp_1 _30555_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2790),
    .D(_02883_),
    .Q_N(_11213_),
    .Q(\scanline[151][0] ));
 sg13g2_dfrbp_1 _30556_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2789),
    .D(_02884_),
    .Q_N(_11212_),
    .Q(\scanline[151][1] ));
 sg13g2_dfrbp_1 _30557_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2788),
    .D(_02885_),
    .Q_N(_11211_),
    .Q(\scanline[151][2] ));
 sg13g2_dfrbp_1 _30558_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2787),
    .D(_02886_),
    .Q_N(_11210_),
    .Q(\scanline[151][3] ));
 sg13g2_dfrbp_1 _30559_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2786),
    .D(_02887_),
    .Q_N(_11209_),
    .Q(\scanline[151][4] ));
 sg13g2_dfrbp_1 _30560_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2785),
    .D(_02888_),
    .Q_N(_11208_),
    .Q(\scanline[151][5] ));
 sg13g2_dfrbp_1 _30561_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2784),
    .D(_02889_),
    .Q_N(_11207_),
    .Q(\scanline[151][6] ));
 sg13g2_dfrbp_1 _30562_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2783),
    .D(_02890_),
    .Q_N(_11206_),
    .Q(\scanline[152][0] ));
 sg13g2_dfrbp_1 _30563_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2782),
    .D(_02891_),
    .Q_N(_11205_),
    .Q(\scanline[152][1] ));
 sg13g2_dfrbp_1 _30564_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2781),
    .D(_02892_),
    .Q_N(_11204_),
    .Q(\scanline[152][2] ));
 sg13g2_dfrbp_1 _30565_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2780),
    .D(_02893_),
    .Q_N(_11203_),
    .Q(\scanline[152][3] ));
 sg13g2_dfrbp_1 _30566_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2779),
    .D(_02894_),
    .Q_N(_11202_),
    .Q(\scanline[152][4] ));
 sg13g2_dfrbp_1 _30567_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2778),
    .D(_02895_),
    .Q_N(_11201_),
    .Q(\scanline[152][5] ));
 sg13g2_dfrbp_1 _30568_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2777),
    .D(_02896_),
    .Q_N(_11200_),
    .Q(\scanline[152][6] ));
 sg13g2_dfrbp_1 _30569_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2776),
    .D(_02897_),
    .Q_N(_11199_),
    .Q(\scanline[153][0] ));
 sg13g2_dfrbp_1 _30570_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2775),
    .D(_02898_),
    .Q_N(_11198_),
    .Q(\scanline[153][1] ));
 sg13g2_dfrbp_1 _30571_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2774),
    .D(_02899_),
    .Q_N(_11197_),
    .Q(\scanline[153][2] ));
 sg13g2_dfrbp_1 _30572_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2773),
    .D(_02900_),
    .Q_N(_11196_),
    .Q(\scanline[153][3] ));
 sg13g2_dfrbp_1 _30573_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2772),
    .D(_02901_),
    .Q_N(_11195_),
    .Q(\scanline[153][4] ));
 sg13g2_dfrbp_1 _30574_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2771),
    .D(_02902_),
    .Q_N(_11194_),
    .Q(\scanline[153][5] ));
 sg13g2_dfrbp_1 _30575_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2770),
    .D(_02903_),
    .Q_N(_11193_),
    .Q(\scanline[153][6] ));
 sg13g2_dfrbp_1 _30576_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2769),
    .D(_02904_),
    .Q_N(_11192_),
    .Q(\scanline[154][0] ));
 sg13g2_dfrbp_1 _30577_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2768),
    .D(_02905_),
    .Q_N(_11191_),
    .Q(\scanline[154][1] ));
 sg13g2_dfrbp_1 _30578_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2767),
    .D(_02906_),
    .Q_N(_11190_),
    .Q(\scanline[154][2] ));
 sg13g2_dfrbp_1 _30579_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2766),
    .D(_02907_),
    .Q_N(_11189_),
    .Q(\scanline[154][3] ));
 sg13g2_dfrbp_1 _30580_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2765),
    .D(_02908_),
    .Q_N(_11188_),
    .Q(\scanline[154][4] ));
 sg13g2_dfrbp_1 _30581_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2764),
    .D(_02909_),
    .Q_N(_11187_),
    .Q(\scanline[154][5] ));
 sg13g2_dfrbp_1 _30582_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2763),
    .D(_02910_),
    .Q_N(_11186_),
    .Q(\scanline[154][6] ));
 sg13g2_dfrbp_1 _30583_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2762),
    .D(_02911_),
    .Q_N(_11185_),
    .Q(\scanline[155][0] ));
 sg13g2_dfrbp_1 _30584_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2761),
    .D(_02912_),
    .Q_N(_11184_),
    .Q(\scanline[155][1] ));
 sg13g2_dfrbp_1 _30585_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2760),
    .D(_02913_),
    .Q_N(_11183_),
    .Q(\scanline[155][2] ));
 sg13g2_dfrbp_1 _30586_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2759),
    .D(_02914_),
    .Q_N(_11182_),
    .Q(\scanline[155][3] ));
 sg13g2_dfrbp_1 _30587_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2758),
    .D(_02915_),
    .Q_N(_11181_),
    .Q(\scanline[155][4] ));
 sg13g2_dfrbp_1 _30588_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2757),
    .D(_02916_),
    .Q_N(_11180_),
    .Q(\scanline[155][5] ));
 sg13g2_dfrbp_1 _30589_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2756),
    .D(_02917_),
    .Q_N(_11179_),
    .Q(\scanline[155][6] ));
 sg13g2_dfrbp_1 _30590_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2755),
    .D(_02918_),
    .Q_N(_11178_),
    .Q(\scanline[156][0] ));
 sg13g2_dfrbp_1 _30591_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2754),
    .D(_02919_),
    .Q_N(_11177_),
    .Q(\scanline[156][1] ));
 sg13g2_dfrbp_1 _30592_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2753),
    .D(_02920_),
    .Q_N(_11176_),
    .Q(\scanline[156][2] ));
 sg13g2_dfrbp_1 _30593_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2752),
    .D(_02921_),
    .Q_N(_11175_),
    .Q(\scanline[156][3] ));
 sg13g2_dfrbp_1 _30594_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2751),
    .D(_02922_),
    .Q_N(_11174_),
    .Q(\scanline[156][4] ));
 sg13g2_dfrbp_1 _30595_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2750),
    .D(_02923_),
    .Q_N(_11173_),
    .Q(\scanline[156][5] ));
 sg13g2_dfrbp_1 _30596_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2749),
    .D(_02924_),
    .Q_N(_11172_),
    .Q(\scanline[156][6] ));
 sg13g2_dfrbp_1 _30597_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2748),
    .D(_02925_),
    .Q_N(_11171_),
    .Q(\scanline[157][0] ));
 sg13g2_dfrbp_1 _30598_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2747),
    .D(_02926_),
    .Q_N(_11170_),
    .Q(\scanline[157][1] ));
 sg13g2_dfrbp_1 _30599_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2746),
    .D(_02927_),
    .Q_N(_11169_),
    .Q(\scanline[157][2] ));
 sg13g2_dfrbp_1 _30600_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2745),
    .D(_02928_),
    .Q_N(_11168_),
    .Q(\scanline[157][3] ));
 sg13g2_dfrbp_1 _30601_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2744),
    .D(_02929_),
    .Q_N(_11167_),
    .Q(\scanline[157][4] ));
 sg13g2_dfrbp_1 _30602_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2743),
    .D(_02930_),
    .Q_N(_11166_),
    .Q(\scanline[157][5] ));
 sg13g2_dfrbp_1 _30603_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2742),
    .D(_02931_),
    .Q_N(_11165_),
    .Q(\scanline[157][6] ));
 sg13g2_dfrbp_1 _30604_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2741),
    .D(_02932_),
    .Q_N(_11164_),
    .Q(\scanline[158][0] ));
 sg13g2_dfrbp_1 _30605_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2740),
    .D(_02933_),
    .Q_N(_11163_),
    .Q(\scanline[158][1] ));
 sg13g2_dfrbp_1 _30606_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2739),
    .D(_02934_),
    .Q_N(_11162_),
    .Q(\scanline[158][2] ));
 sg13g2_dfrbp_1 _30607_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2738),
    .D(_02935_),
    .Q_N(_11161_),
    .Q(\scanline[158][3] ));
 sg13g2_dfrbp_1 _30608_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2737),
    .D(_02936_),
    .Q_N(_11160_),
    .Q(\scanline[158][4] ));
 sg13g2_dfrbp_1 _30609_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2736),
    .D(_02937_),
    .Q_N(_11159_),
    .Q(\scanline[158][5] ));
 sg13g2_dfrbp_1 _30610_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2735),
    .D(_02938_),
    .Q_N(_11158_),
    .Q(\scanline[158][6] ));
 sg13g2_dfrbp_1 _30611_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2734),
    .D(_02939_),
    .Q_N(_11157_),
    .Q(\scanline[15][0] ));
 sg13g2_dfrbp_1 _30612_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2733),
    .D(_02940_),
    .Q_N(_11156_),
    .Q(\scanline[15][1] ));
 sg13g2_dfrbp_1 _30613_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2732),
    .D(_02941_),
    .Q_N(_11155_),
    .Q(\scanline[15][2] ));
 sg13g2_dfrbp_1 _30614_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2731),
    .D(_02942_),
    .Q_N(_11154_),
    .Q(\scanline[15][3] ));
 sg13g2_dfrbp_1 _30615_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2730),
    .D(_02943_),
    .Q_N(_11153_),
    .Q(\scanline[15][4] ));
 sg13g2_dfrbp_1 _30616_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2729),
    .D(_02944_),
    .Q_N(_11152_),
    .Q(\scanline[15][5] ));
 sg13g2_dfrbp_1 _30617_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2728),
    .D(_02945_),
    .Q_N(_11151_),
    .Q(\scanline[15][6] ));
 sg13g2_dfrbp_1 _30618_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2727),
    .D(_02946_),
    .Q_N(_11150_),
    .Q(\scanline[16][0] ));
 sg13g2_dfrbp_1 _30619_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2726),
    .D(_02947_),
    .Q_N(_11149_),
    .Q(\scanline[16][1] ));
 sg13g2_dfrbp_1 _30620_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2725),
    .D(_02948_),
    .Q_N(_11148_),
    .Q(\scanline[16][2] ));
 sg13g2_dfrbp_1 _30621_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2724),
    .D(_02949_),
    .Q_N(_11147_),
    .Q(\scanline[16][3] ));
 sg13g2_dfrbp_1 _30622_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2723),
    .D(_02950_),
    .Q_N(_11146_),
    .Q(\scanline[16][4] ));
 sg13g2_dfrbp_1 _30623_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2722),
    .D(_02951_),
    .Q_N(_11145_),
    .Q(\scanline[16][5] ));
 sg13g2_dfrbp_1 _30624_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2721),
    .D(_02952_),
    .Q_N(_11144_),
    .Q(\scanline[16][6] ));
 sg13g2_dfrbp_1 _30625_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2720),
    .D(_02953_),
    .Q_N(_11143_),
    .Q(\scanline[17][0] ));
 sg13g2_dfrbp_1 _30626_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2719),
    .D(_02954_),
    .Q_N(_11142_),
    .Q(\scanline[17][1] ));
 sg13g2_dfrbp_1 _30627_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2718),
    .D(_02955_),
    .Q_N(_11141_),
    .Q(\scanline[17][2] ));
 sg13g2_dfrbp_1 _30628_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2717),
    .D(_02956_),
    .Q_N(_11140_),
    .Q(\scanline[17][3] ));
 sg13g2_dfrbp_1 _30629_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2716),
    .D(_02957_),
    .Q_N(_11139_),
    .Q(\scanline[17][4] ));
 sg13g2_dfrbp_1 _30630_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2715),
    .D(_02958_),
    .Q_N(_11138_),
    .Q(\scanline[17][5] ));
 sg13g2_dfrbp_1 _30631_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2714),
    .D(_02959_),
    .Q_N(_11137_),
    .Q(\scanline[17][6] ));
 sg13g2_dfrbp_1 _30632_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2713),
    .D(_02960_),
    .Q_N(_11136_),
    .Q(\scanline[18][0] ));
 sg13g2_dfrbp_1 _30633_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2712),
    .D(_02961_),
    .Q_N(_11135_),
    .Q(\scanline[18][1] ));
 sg13g2_dfrbp_1 _30634_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2711),
    .D(_02962_),
    .Q_N(_11134_),
    .Q(\scanline[18][2] ));
 sg13g2_dfrbp_1 _30635_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2710),
    .D(_02963_),
    .Q_N(_11133_),
    .Q(\scanline[18][3] ));
 sg13g2_dfrbp_1 _30636_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2709),
    .D(_02964_),
    .Q_N(_11132_),
    .Q(\scanline[18][4] ));
 sg13g2_dfrbp_1 _30637_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2708),
    .D(_02965_),
    .Q_N(_11131_),
    .Q(\scanline[18][5] ));
 sg13g2_dfrbp_1 _30638_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2707),
    .D(_02966_),
    .Q_N(_11130_),
    .Q(\scanline[18][6] ));
 sg13g2_dfrbp_1 _30639_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2706),
    .D(_02967_),
    .Q_N(_11129_),
    .Q(\scanline[1][0] ));
 sg13g2_dfrbp_1 _30640_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2705),
    .D(_02968_),
    .Q_N(_11128_),
    .Q(\scanline[1][1] ));
 sg13g2_dfrbp_1 _30641_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2704),
    .D(_02969_),
    .Q_N(_11127_),
    .Q(\scanline[1][2] ));
 sg13g2_dfrbp_1 _30642_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2703),
    .D(_02970_),
    .Q_N(_11126_),
    .Q(\scanline[1][3] ));
 sg13g2_dfrbp_1 _30643_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2702),
    .D(_02971_),
    .Q_N(_11125_),
    .Q(\scanline[1][4] ));
 sg13g2_dfrbp_1 _30644_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2701),
    .D(_02972_),
    .Q_N(_11124_),
    .Q(\scanline[1][5] ));
 sg13g2_dfrbp_1 _30645_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2700),
    .D(_02973_),
    .Q_N(_11123_),
    .Q(\scanline[1][6] ));
 sg13g2_dfrbp_1 _30646_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1982),
    .D(_02974_),
    .Q_N(_11122_),
    .Q(\scanline[20][0] ));
 sg13g2_dfrbp_1 _30647_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1980),
    .D(_02975_),
    .Q_N(_11121_),
    .Q(\scanline[20][1] ));
 sg13g2_dfrbp_1 _30648_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1978),
    .D(_02976_),
    .Q_N(_11120_),
    .Q(\scanline[20][2] ));
 sg13g2_dfrbp_1 _30649_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1951),
    .D(_02977_),
    .Q_N(_11119_),
    .Q(\scanline[20][3] ));
 sg13g2_dfrbp_1 _30650_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1949),
    .D(_02978_),
    .Q_N(_11118_),
    .Q(\scanline[20][4] ));
 sg13g2_dfrbp_1 _30651_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1947),
    .D(_02979_),
    .Q_N(_11117_),
    .Q(\scanline[20][5] ));
 sg13g2_dfrbp_1 _30652_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1945),
    .D(_02980_),
    .Q_N(_11116_),
    .Q(\scanline[20][6] ));
 sg13g2_dfrbp_1 _30653_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1848),
    .D(_02981_),
    .Q_N(_11115_),
    .Q(\scanline[21][0] ));
 sg13g2_dfrbp_1 _30654_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1846),
    .D(_02982_),
    .Q_N(_11114_),
    .Q(\scanline[21][1] ));
 sg13g2_dfrbp_1 _30655_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1844),
    .D(_02983_),
    .Q_N(_11113_),
    .Q(\scanline[21][2] ));
 sg13g2_dfrbp_1 _30656_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1842),
    .D(_02984_),
    .Q_N(_11112_),
    .Q(\scanline[21][3] ));
 sg13g2_dfrbp_1 _30657_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1840),
    .D(_02985_),
    .Q_N(_11111_),
    .Q(\scanline[21][4] ));
 sg13g2_dfrbp_1 _30658_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1838),
    .D(_02986_),
    .Q_N(_11110_),
    .Q(\scanline[21][5] ));
 sg13g2_dfrbp_1 _30659_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1833),
    .D(_02987_),
    .Q_N(_11109_),
    .Q(\scanline[21][6] ));
 sg13g2_dfrbp_1 _30660_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1753),
    .D(_02988_),
    .Q_N(_11108_),
    .Q(\scanline[22][0] ));
 sg13g2_dfrbp_1 _30661_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1751),
    .D(_02989_),
    .Q_N(_11107_),
    .Q(\scanline[22][1] ));
 sg13g2_dfrbp_1 _30662_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1749),
    .D(_02990_),
    .Q_N(_11106_),
    .Q(\scanline[22][2] ));
 sg13g2_dfrbp_1 _30663_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1747),
    .D(_02991_),
    .Q_N(_11105_),
    .Q(\scanline[22][3] ));
 sg13g2_dfrbp_1 _30664_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1745),
    .D(_02992_),
    .Q_N(_11104_),
    .Q(\scanline[22][4] ));
 sg13g2_dfrbp_1 _30665_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1743),
    .D(_02993_),
    .Q_N(_11103_),
    .Q(\scanline[22][5] ));
 sg13g2_dfrbp_1 _30666_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1741),
    .D(_02994_),
    .Q_N(_11102_),
    .Q(\scanline[22][6] ));
 sg13g2_dfrbp_1 _30667_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1676),
    .D(_02995_),
    .Q_N(_11101_),
    .Q(\scanline[23][0] ));
 sg13g2_dfrbp_1 _30668_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1674),
    .D(_02996_),
    .Q_N(_11100_),
    .Q(\scanline[23][1] ));
 sg13g2_dfrbp_1 _30669_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1672),
    .D(_02997_),
    .Q_N(_11099_),
    .Q(\scanline[23][2] ));
 sg13g2_dfrbp_1 _30670_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1670),
    .D(_02998_),
    .Q_N(_11098_),
    .Q(\scanline[23][3] ));
 sg13g2_dfrbp_1 _30671_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1668),
    .D(_02999_),
    .Q_N(_11097_),
    .Q(\scanline[23][4] ));
 sg13g2_dfrbp_1 _30672_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1666),
    .D(_03000_),
    .Q_N(_11096_),
    .Q(\scanline[23][5] ));
 sg13g2_dfrbp_1 _30673_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1664),
    .D(_03001_),
    .Q_N(_11095_),
    .Q(\scanline[23][6] ));
 sg13g2_dfrbp_1 _30674_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1397),
    .D(_03002_),
    .Q_N(_11094_),
    .Q(\scanline[24][0] ));
 sg13g2_dfrbp_1 _30675_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1395),
    .D(_03003_),
    .Q_N(_11093_),
    .Q(\scanline[24][1] ));
 sg13g2_dfrbp_1 _30676_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1393),
    .D(_03004_),
    .Q_N(_11092_),
    .Q(\scanline[24][2] ));
 sg13g2_dfrbp_1 _30677_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1391),
    .D(_03005_),
    .Q_N(_11091_),
    .Q(\scanline[24][3] ));
 sg13g2_dfrbp_1 _30678_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1389),
    .D(_03006_),
    .Q_N(_11090_),
    .Q(\scanline[24][4] ));
 sg13g2_dfrbp_1 _30679_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1387),
    .D(_03007_),
    .Q_N(_11089_),
    .Q(\scanline[24][5] ));
 sg13g2_dfrbp_1 _30680_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1385),
    .D(_03008_),
    .Q_N(_11088_),
    .Q(\scanline[24][6] ));
 sg13g2_dfrbp_1 _30681_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1007),
    .D(_03009_),
    .Q_N(_11087_),
    .Q(\atari2600.cpu.dst_reg[1] ));
 sg13g2_dfrbp_1 _30682_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1003),
    .D(_03010_),
    .Q_N(_11086_),
    .Q(\atari2600.cpu.dst_reg[0] ));
 sg13g2_dfrbp_1 _30683_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net999),
    .D(_03011_),
    .Q_N(_00072_),
    .Q(\atari2600.cpu.src_reg[1] ));
 sg13g2_dfrbp_1 _30684_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net987),
    .D(_03012_),
    .Q_N(_00071_),
    .Q(\atari2600.cpu.src_reg[0] ));
 sg13g2_dfrbp_1 _30685_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net983),
    .D(_03013_),
    .Q_N(_11085_),
    .Q(\atari2600.cpu.op[3] ));
 sg13g2_dfrbp_1 _30686_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net979),
    .D(_03014_),
    .Q_N(_11084_),
    .Q(\atari2600.cpu.op[2] ));
 sg13g2_dfrbp_1 _30687_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1001),
    .D(_03015_),
    .Q_N(_11083_),
    .Q(\atari2600.cpu.op[1] ));
 sg13g2_dfrbp_1 _30688_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net985),
    .D(_03016_),
    .Q_N(_11082_),
    .Q(\atari2600.cpu.op[0] ));
 sg13g2_dfrbp_1 _30689_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1005),
    .D(_03017_),
    .Q_N(_11081_),
    .Q(\atari2600.tia.dat_o[7] ));
 sg13g2_dfrbp_1 _30690_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net981),
    .D(_03018_),
    .Q_N(_11080_),
    .Q(\atari2600.tia.dat_o[6] ));
 sg13g2_tiehi _30421__14 (.L_HI(net14));
 sg13g2_tiehi _30420__15 (.L_HI(net15));
 sg13g2_tiehi _30419__16 (.L_HI(net16));
 sg13g2_tiehi _30418__17 (.L_HI(net17));
 sg13g2_tiehi _30417__18 (.L_HI(net18));
 sg13g2_tiehi _30416__19 (.L_HI(net19));
 sg13g2_tiehi _30415__20 (.L_HI(net20));
 sg13g2_tiehi _30414__21 (.L_HI(net21));
 sg13g2_tiehi _30413__22 (.L_HI(net22));
 sg13g2_tiehi _30412__23 (.L_HI(net23));
 sg13g2_tiehi _30411__24 (.L_HI(net24));
 sg13g2_tiehi _30410__25 (.L_HI(net25));
 sg13g2_tiehi _30409__26 (.L_HI(net26));
 sg13g2_tiehi _30408__27 (.L_HI(net27));
 sg13g2_tiehi _30407__28 (.L_HI(net28));
 sg13g2_tiehi _30406__29 (.L_HI(net29));
 sg13g2_tiehi _30405__30 (.L_HI(net30));
 sg13g2_tiehi _30404__31 (.L_HI(net31));
 sg13g2_tiehi _30403__32 (.L_HI(net32));
 sg13g2_tiehi _30402__33 (.L_HI(net33));
 sg13g2_tiehi _30401__34 (.L_HI(net34));
 sg13g2_tiehi _30400__35 (.L_HI(net35));
 sg13g2_tiehi _30399__36 (.L_HI(net36));
 sg13g2_tiehi _30398__37 (.L_HI(net37));
 sg13g2_tiehi _30397__38 (.L_HI(net38));
 sg13g2_tiehi _30396__39 (.L_HI(net39));
 sg13g2_tiehi _30395__40 (.L_HI(net40));
 sg13g2_tiehi _30394__41 (.L_HI(net41));
 sg13g2_tiehi _30393__42 (.L_HI(net42));
 sg13g2_tiehi _30392__43 (.L_HI(net43));
 sg13g2_tiehi _30391__44 (.L_HI(net44));
 sg13g2_tiehi _30390__45 (.L_HI(net45));
 sg13g2_tiehi _30389__46 (.L_HI(net46));
 sg13g2_tiehi _30388__47 (.L_HI(net47));
 sg13g2_tiehi _30387__48 (.L_HI(net48));
 sg13g2_tiehi _30386__49 (.L_HI(net49));
 sg13g2_tiehi _30385__50 (.L_HI(net50));
 sg13g2_tiehi _30384__51 (.L_HI(net51));
 sg13g2_tiehi _30383__52 (.L_HI(net52));
 sg13g2_tiehi _30382__53 (.L_HI(net53));
 sg13g2_tiehi _30381__54 (.L_HI(net54));
 sg13g2_tiehi _30380__55 (.L_HI(net55));
 sg13g2_tiehi _30379__56 (.L_HI(net56));
 sg13g2_tiehi _30378__57 (.L_HI(net57));
 sg13g2_tiehi _30377__58 (.L_HI(net58));
 sg13g2_tiehi _30376__59 (.L_HI(net59));
 sg13g2_tiehi _30375__60 (.L_HI(net60));
 sg13g2_tiehi _30374__61 (.L_HI(net61));
 sg13g2_tiehi _30373__62 (.L_HI(net62));
 sg13g2_tiehi _30372__63 (.L_HI(net63));
 sg13g2_tiehi _30371__64 (.L_HI(net64));
 sg13g2_tiehi _30370__65 (.L_HI(net65));
 sg13g2_tiehi _30369__66 (.L_HI(net66));
 sg13g2_tiehi _30368__67 (.L_HI(net67));
 sg13g2_tiehi _30367__68 (.L_HI(net68));
 sg13g2_tiehi _30366__69 (.L_HI(net69));
 sg13g2_tiehi _30365__70 (.L_HI(net70));
 sg13g2_tiehi _30364__71 (.L_HI(net71));
 sg13g2_tiehi _30363__72 (.L_HI(net72));
 sg13g2_tiehi _30362__73 (.L_HI(net73));
 sg13g2_tiehi _30361__74 (.L_HI(net74));
 sg13g2_tiehi _30360__75 (.L_HI(net75));
 sg13g2_tiehi _30359__76 (.L_HI(net76));
 sg13g2_tiehi _30358__77 (.L_HI(net77));
 sg13g2_tiehi _30357__78 (.L_HI(net78));
 sg13g2_tiehi _30356__79 (.L_HI(net79));
 sg13g2_tiehi _30355__80 (.L_HI(net80));
 sg13g2_tiehi _30354__81 (.L_HI(net81));
 sg13g2_tiehi _30353__82 (.L_HI(net82));
 sg13g2_tiehi _30352__83 (.L_HI(net83));
 sg13g2_tiehi _30351__84 (.L_HI(net84));
 sg13g2_tiehi _30350__85 (.L_HI(net85));
 sg13g2_tiehi _30349__86 (.L_HI(net86));
 sg13g2_tiehi _30348__87 (.L_HI(net87));
 sg13g2_tiehi _30347__88 (.L_HI(net88));
 sg13g2_tiehi _30346__89 (.L_HI(net89));
 sg13g2_tiehi _30345__90 (.L_HI(net90));
 sg13g2_tiehi _30344__91 (.L_HI(net91));
 sg13g2_tiehi _30343__92 (.L_HI(net92));
 sg13g2_tiehi _30342__93 (.L_HI(net93));
 sg13g2_tiehi _30341__94 (.L_HI(net94));
 sg13g2_tiehi _30340__95 (.L_HI(net95));
 sg13g2_tiehi _30339__96 (.L_HI(net96));
 sg13g2_tiehi _30338__97 (.L_HI(net97));
 sg13g2_tiehi _27775__98 (.L_HI(net98));
 sg13g2_tiehi _27859__99 (.L_HI(net99));
 sg13g2_tiehi _30337__100 (.L_HI(net100));
 sg13g2_tiehi _30336__101 (.L_HI(net101));
 sg13g2_tiehi _30335__102 (.L_HI(net102));
 sg13g2_tiehi _30334__103 (.L_HI(net103));
 sg13g2_tiehi _30333__104 (.L_HI(net104));
 sg13g2_tiehi _30332__105 (.L_HI(net105));
 sg13g2_tiehi _30331__106 (.L_HI(net106));
 sg13g2_tiehi _30330__107 (.L_HI(net107));
 sg13g2_tiehi _30329__108 (.L_HI(net108));
 sg13g2_tiehi _30328__109 (.L_HI(net109));
 sg13g2_tiehi _30327__110 (.L_HI(net110));
 sg13g2_tiehi _30326__111 (.L_HI(net111));
 sg13g2_tiehi _30325__112 (.L_HI(net112));
 sg13g2_tiehi _30324__113 (.L_HI(net113));
 sg13g2_tiehi _30323__114 (.L_HI(net114));
 sg13g2_tiehi _30322__115 (.L_HI(net115));
 sg13g2_tiehi _30321__116 (.L_HI(net116));
 sg13g2_tiehi _30320__117 (.L_HI(net117));
 sg13g2_tiehi _30319__118 (.L_HI(net118));
 sg13g2_tiehi _30318__119 (.L_HI(net119));
 sg13g2_tiehi _30317__120 (.L_HI(net120));
 sg13g2_tiehi _30316__121 (.L_HI(net121));
 sg13g2_tiehi _30315__122 (.L_HI(net122));
 sg13g2_tiehi _30314__123 (.L_HI(net123));
 sg13g2_tiehi _30313__124 (.L_HI(net124));
 sg13g2_tiehi _30312__125 (.L_HI(net125));
 sg13g2_tiehi _30311__126 (.L_HI(net126));
 sg13g2_tiehi _30310__127 (.L_HI(net127));
 sg13g2_tiehi _30309__128 (.L_HI(net128));
 sg13g2_tiehi _30308__129 (.L_HI(net129));
 sg13g2_tiehi _30307__130 (.L_HI(net130));
 sg13g2_tiehi _30306__131 (.L_HI(net131));
 sg13g2_tiehi _30305__132 (.L_HI(net132));
 sg13g2_tiehi _30304__133 (.L_HI(net133));
 sg13g2_tiehi _30303__134 (.L_HI(net134));
 sg13g2_tiehi _30302__135 (.L_HI(net135));
 sg13g2_tiehi _30301__136 (.L_HI(net136));
 sg13g2_tiehi _30300__137 (.L_HI(net137));
 sg13g2_tiehi _30299__138 (.L_HI(net138));
 sg13g2_tiehi _30298__139 (.L_HI(net139));
 sg13g2_tiehi _30297__140 (.L_HI(net140));
 sg13g2_tiehi _30296__141 (.L_HI(net141));
 sg13g2_tiehi _30295__142 (.L_HI(net142));
 sg13g2_tiehi _30294__143 (.L_HI(net143));
 sg13g2_tiehi _30293__144 (.L_HI(net144));
 sg13g2_tiehi _30292__145 (.L_HI(net145));
 sg13g2_tiehi _30291__146 (.L_HI(net146));
 sg13g2_tiehi _30290__147 (.L_HI(net147));
 sg13g2_tiehi _30289__148 (.L_HI(net148));
 sg13g2_tiehi _30288__149 (.L_HI(net149));
 sg13g2_tiehi _30287__150 (.L_HI(net150));
 sg13g2_tiehi _30286__151 (.L_HI(net151));
 sg13g2_tiehi _30285__152 (.L_HI(net152));
 sg13g2_tiehi _30284__153 (.L_HI(net153));
 sg13g2_tiehi _30283__154 (.L_HI(net154));
 sg13g2_tiehi _30282__155 (.L_HI(net155));
 sg13g2_tiehi _30281__156 (.L_HI(net156));
 sg13g2_tiehi _30280__157 (.L_HI(net157));
 sg13g2_tiehi _30279__158 (.L_HI(net158));
 sg13g2_tiehi _30278__159 (.L_HI(net159));
 sg13g2_tiehi _30277__160 (.L_HI(net160));
 sg13g2_tiehi _30276__161 (.L_HI(net161));
 sg13g2_tiehi _30275__162 (.L_HI(net162));
 sg13g2_tiehi _30274__163 (.L_HI(net163));
 sg13g2_tiehi _30273__164 (.L_HI(net164));
 sg13g2_tiehi _30272__165 (.L_HI(net165));
 sg13g2_tiehi _30271__166 (.L_HI(net166));
 sg13g2_tiehi _30270__167 (.L_HI(net167));
 sg13g2_tiehi _30269__168 (.L_HI(net168));
 sg13g2_tiehi _30268__169 (.L_HI(net169));
 sg13g2_tiehi _30267__170 (.L_HI(net170));
 sg13g2_tiehi _30266__171 (.L_HI(net171));
 sg13g2_tiehi _30265__172 (.L_HI(net172));
 sg13g2_tiehi _30264__173 (.L_HI(net173));
 sg13g2_tiehi _30263__174 (.L_HI(net174));
 sg13g2_tiehi _30262__175 (.L_HI(net175));
 sg13g2_tiehi _30261__176 (.L_HI(net176));
 sg13g2_tiehi _30260__177 (.L_HI(net177));
 sg13g2_tiehi _30259__178 (.L_HI(net178));
 sg13g2_tiehi _30258__179 (.L_HI(net179));
 sg13g2_tiehi _30257__180 (.L_HI(net180));
 sg13g2_tiehi _30256__181 (.L_HI(net181));
 sg13g2_tiehi _30255__182 (.L_HI(net182));
 sg13g2_tiehi _30254__183 (.L_HI(net183));
 sg13g2_tiehi _30253__184 (.L_HI(net184));
 sg13g2_tiehi _30252__185 (.L_HI(net185));
 sg13g2_tiehi _30251__186 (.L_HI(net186));
 sg13g2_tiehi _30250__187 (.L_HI(net187));
 sg13g2_tiehi _27860__188 (.L_HI(net188));
 sg13g2_tiehi _30249__189 (.L_HI(net189));
 sg13g2_tiehi _30248__190 (.L_HI(net190));
 sg13g2_tiehi _30247__191 (.L_HI(net191));
 sg13g2_tiehi _30246__192 (.L_HI(net192));
 sg13g2_tiehi _30245__193 (.L_HI(net193));
 sg13g2_tiehi _30244__194 (.L_HI(net194));
 sg13g2_tiehi _30243__195 (.L_HI(net195));
 sg13g2_tiehi _30242__196 (.L_HI(net196));
 sg13g2_tiehi _30241__197 (.L_HI(net197));
 sg13g2_tiehi _30240__198 (.L_HI(net198));
 sg13g2_tiehi _30239__199 (.L_HI(net199));
 sg13g2_tiehi _30238__200 (.L_HI(net200));
 sg13g2_tiehi _30237__201 (.L_HI(net201));
 sg13g2_tiehi _30236__202 (.L_HI(net202));
 sg13g2_tiehi _30235__203 (.L_HI(net203));
 sg13g2_tiehi _30234__204 (.L_HI(net204));
 sg13g2_tiehi _30233__205 (.L_HI(net205));
 sg13g2_tiehi _30232__206 (.L_HI(net206));
 sg13g2_tiehi _30231__207 (.L_HI(net207));
 sg13g2_tiehi _30230__208 (.L_HI(net208));
 sg13g2_tiehi _30229__209 (.L_HI(net209));
 sg13g2_tiehi _30228__210 (.L_HI(net210));
 sg13g2_tiehi _30227__211 (.L_HI(net211));
 sg13g2_tiehi _30226__212 (.L_HI(net212));
 sg13g2_tiehi _30225__213 (.L_HI(net213));
 sg13g2_tiehi _30224__214 (.L_HI(net214));
 sg13g2_tiehi _30223__215 (.L_HI(net215));
 sg13g2_tiehi _30222__216 (.L_HI(net216));
 sg13g2_tiehi _30221__217 (.L_HI(net217));
 sg13g2_tiehi _27949__218 (.L_HI(net218));
 sg13g2_tiehi _27979__219 (.L_HI(net219));
 sg13g2_tiehi _30220__220 (.L_HI(net220));
 sg13g2_tiehi _30219__221 (.L_HI(net221));
 sg13g2_tiehi _30218__222 (.L_HI(net222));
 sg13g2_tiehi _30217__223 (.L_HI(net223));
 sg13g2_tiehi _30216__224 (.L_HI(net224));
 sg13g2_tiehi _30215__225 (.L_HI(net225));
 sg13g2_tiehi _30214__226 (.L_HI(net226));
 sg13g2_tiehi _30213__227 (.L_HI(net227));
 sg13g2_tiehi _30212__228 (.L_HI(net228));
 sg13g2_tiehi _30211__229 (.L_HI(net229));
 sg13g2_tiehi _30210__230 (.L_HI(net230));
 sg13g2_tiehi _30209__231 (.L_HI(net231));
 sg13g2_tiehi _30208__232 (.L_HI(net232));
 sg13g2_tiehi _30207__233 (.L_HI(net233));
 sg13g2_tiehi _30206__234 (.L_HI(net234));
 sg13g2_tiehi _30205__235 (.L_HI(net235));
 sg13g2_tiehi _30204__236 (.L_HI(net236));
 sg13g2_tiehi _30203__237 (.L_HI(net237));
 sg13g2_tiehi _30202__238 (.L_HI(net238));
 sg13g2_tiehi _30201__239 (.L_HI(net239));
 sg13g2_tiehi _30200__240 (.L_HI(net240));
 sg13g2_tiehi _30199__241 (.L_HI(net241));
 sg13g2_tiehi _30198__242 (.L_HI(net242));
 sg13g2_tiehi _30197__243 (.L_HI(net243));
 sg13g2_tiehi _30196__244 (.L_HI(net244));
 sg13g2_tiehi _30195__245 (.L_HI(net245));
 sg13g2_tiehi _30194__246 (.L_HI(net246));
 sg13g2_tiehi _30193__247 (.L_HI(net247));
 sg13g2_tiehi _30192__248 (.L_HI(net248));
 sg13g2_tiehi _30191__249 (.L_HI(net249));
 sg13g2_tiehi _30190__250 (.L_HI(net250));
 sg13g2_tiehi _30189__251 (.L_HI(net251));
 sg13g2_tiehi _30188__252 (.L_HI(net252));
 sg13g2_tiehi _30187__253 (.L_HI(net253));
 sg13g2_tiehi _30186__254 (.L_HI(net254));
 sg13g2_tiehi _30185__255 (.L_HI(net255));
 sg13g2_tiehi _30184__256 (.L_HI(net256));
 sg13g2_tiehi _30183__257 (.L_HI(net257));
 sg13g2_tiehi _30182__258 (.L_HI(net258));
 sg13g2_tiehi _30181__259 (.L_HI(net259));
 sg13g2_tiehi _30180__260 (.L_HI(net260));
 sg13g2_tiehi _30179__261 (.L_HI(net261));
 sg13g2_tiehi _30178__262 (.L_HI(net262));
 sg13g2_tiehi _30177__263 (.L_HI(net263));
 sg13g2_tiehi _30176__264 (.L_HI(net264));
 sg13g2_tiehi _30175__265 (.L_HI(net265));
 sg13g2_tiehi _30174__266 (.L_HI(net266));
 sg13g2_tiehi _30173__267 (.L_HI(net267));
 sg13g2_tiehi _30172__268 (.L_HI(net268));
 sg13g2_tiehi _30171__269 (.L_HI(net269));
 sg13g2_tiehi _30170__270 (.L_HI(net270));
 sg13g2_tiehi _30169__271 (.L_HI(net271));
 sg13g2_tiehi _30168__272 (.L_HI(net272));
 sg13g2_tiehi _30167__273 (.L_HI(net273));
 sg13g2_tiehi _30166__274 (.L_HI(net274));
 sg13g2_tiehi _30165__275 (.L_HI(net275));
 sg13g2_tiehi _30164__276 (.L_HI(net276));
 sg13g2_tiehi _30163__277 (.L_HI(net277));
 sg13g2_tiehi _30162__278 (.L_HI(net278));
 sg13g2_tiehi _30161__279 (.L_HI(net279));
 sg13g2_tiehi _30160__280 (.L_HI(net280));
 sg13g2_tiehi _30159__281 (.L_HI(net281));
 sg13g2_tiehi _30158__282 (.L_HI(net282));
 sg13g2_tiehi _30157__283 (.L_HI(net283));
 sg13g2_tiehi _30156__284 (.L_HI(net284));
 sg13g2_tiehi _30155__285 (.L_HI(net285));
 sg13g2_tiehi _30154__286 (.L_HI(net286));
 sg13g2_tiehi _30153__287 (.L_HI(net287));
 sg13g2_tiehi _30152__288 (.L_HI(net288));
 sg13g2_tiehi _30151__289 (.L_HI(net289));
 sg13g2_tiehi _30150__290 (.L_HI(net290));
 sg13g2_tiehi _30149__291 (.L_HI(net291));
 sg13g2_tiehi _30148__292 (.L_HI(net292));
 sg13g2_tiehi _30147__293 (.L_HI(net293));
 sg13g2_tiehi _30146__294 (.L_HI(net294));
 sg13g2_tiehi _30145__295 (.L_HI(net295));
 sg13g2_tiehi _30144__296 (.L_HI(net296));
 sg13g2_tiehi _30143__297 (.L_HI(net297));
 sg13g2_tiehi _30142__298 (.L_HI(net298));
 sg13g2_tiehi _30141__299 (.L_HI(net299));
 sg13g2_tiehi _30140__300 (.L_HI(net300));
 sg13g2_tiehi _28065__301 (.L_HI(net301));
 sg13g2_tiehi _28066__302 (.L_HI(net302));
 sg13g2_tiehi _28067__303 (.L_HI(net303));
 sg13g2_tiehi _28068__304 (.L_HI(net304));
 sg13g2_tiehi _28069__305 (.L_HI(net305));
 sg13g2_tiehi _28070__306 (.L_HI(net306));
 sg13g2_tiehi _28071__307 (.L_HI(net307));
 sg13g2_tiehi _30139__308 (.L_HI(net308));
 sg13g2_tiehi _30138__309 (.L_HI(net309));
 sg13g2_tiehi _30137__310 (.L_HI(net310));
 sg13g2_tiehi _30136__311 (.L_HI(net311));
 sg13g2_tiehi _30135__312 (.L_HI(net312));
 sg13g2_tiehi _30134__313 (.L_HI(net313));
 sg13g2_tiehi _30133__314 (.L_HI(net314));
 sg13g2_tiehi _30132__315 (.L_HI(net315));
 sg13g2_tiehi _30131__316 (.L_HI(net316));
 sg13g2_tiehi _30130__317 (.L_HI(net317));
 sg13g2_tiehi _30129__318 (.L_HI(net318));
 sg13g2_tiehi _30128__319 (.L_HI(net319));
 sg13g2_tiehi _30127__320 (.L_HI(net320));
 sg13g2_tiehi _30126__321 (.L_HI(net321));
 sg13g2_tiehi _30125__322 (.L_HI(net322));
 sg13g2_tiehi _30124__323 (.L_HI(net323));
 sg13g2_tiehi _30123__324 (.L_HI(net324));
 sg13g2_tiehi _30122__325 (.L_HI(net325));
 sg13g2_tiehi _30121__326 (.L_HI(net326));
 sg13g2_tiehi _30120__327 (.L_HI(net327));
 sg13g2_tiehi _30119__328 (.L_HI(net328));
 sg13g2_tiehi _30118__329 (.L_HI(net329));
 sg13g2_tiehi _30117__330 (.L_HI(net330));
 sg13g2_tiehi _30116__331 (.L_HI(net331));
 sg13g2_tiehi _30115__332 (.L_HI(net332));
 sg13g2_tiehi _30114__333 (.L_HI(net333));
 sg13g2_tiehi _30113__334 (.L_HI(net334));
 sg13g2_tiehi _30112__335 (.L_HI(net335));
 sg13g2_tiehi _30111__336 (.L_HI(net336));
 sg13g2_tiehi _30110__337 (.L_HI(net337));
 sg13g2_tiehi _30109__338 (.L_HI(net338));
 sg13g2_tiehi _30108__339 (.L_HI(net339));
 sg13g2_tiehi _30107__340 (.L_HI(net340));
 sg13g2_tiehi _30106__341 (.L_HI(net341));
 sg13g2_tiehi _30105__342 (.L_HI(net342));
 sg13g2_tiehi _30104__343 (.L_HI(net343));
 sg13g2_tiehi _30103__344 (.L_HI(net344));
 sg13g2_tiehi _30102__345 (.L_HI(net345));
 sg13g2_tiehi _30101__346 (.L_HI(net346));
 sg13g2_tiehi _30100__347 (.L_HI(net347));
 sg13g2_tiehi _30099__348 (.L_HI(net348));
 sg13g2_tiehi _30098__349 (.L_HI(net349));
 sg13g2_tiehi _30097__350 (.L_HI(net350));
 sg13g2_tiehi _30096__351 (.L_HI(net351));
 sg13g2_tiehi _30095__352 (.L_HI(net352));
 sg13g2_tiehi _30094__353 (.L_HI(net353));
 sg13g2_tiehi _30093__354 (.L_HI(net354));
 sg13g2_tiehi _30092__355 (.L_HI(net355));
 sg13g2_tiehi _30091__356 (.L_HI(net356));
 sg13g2_tiehi _30090__357 (.L_HI(net357));
 sg13g2_tiehi _30089__358 (.L_HI(net358));
 sg13g2_tiehi _30088__359 (.L_HI(net359));
 sg13g2_tiehi _30087__360 (.L_HI(net360));
 sg13g2_tiehi _30086__361 (.L_HI(net361));
 sg13g2_tiehi _30085__362 (.L_HI(net362));
 sg13g2_tiehi _30084__363 (.L_HI(net363));
 sg13g2_tiehi _30083__364 (.L_HI(net364));
 sg13g2_tiehi _30082__365 (.L_HI(net365));
 sg13g2_tiehi _30081__366 (.L_HI(net366));
 sg13g2_tiehi _30080__367 (.L_HI(net367));
 sg13g2_tiehi _30079__368 (.L_HI(net368));
 sg13g2_tiehi _30078__369 (.L_HI(net369));
 sg13g2_tiehi _30077__370 (.L_HI(net370));
 sg13g2_tiehi _30076__371 (.L_HI(net371));
 sg13g2_tiehi _30075__372 (.L_HI(net372));
 sg13g2_tiehi _30074__373 (.L_HI(net373));
 sg13g2_tiehi _30073__374 (.L_HI(net374));
 sg13g2_tiehi _30072__375 (.L_HI(net375));
 sg13g2_tiehi _30071__376 (.L_HI(net376));
 sg13g2_tiehi _30070__377 (.L_HI(net377));
 sg13g2_tiehi _30069__378 (.L_HI(net378));
 sg13g2_tiehi _30068__379 (.L_HI(net379));
 sg13g2_tiehi _30067__380 (.L_HI(net380));
 sg13g2_tiehi _30066__381 (.L_HI(net381));
 sg13g2_tiehi _30065__382 (.L_HI(net382));
 sg13g2_tiehi _30064__383 (.L_HI(net383));
 sg13g2_tiehi _30063__384 (.L_HI(net384));
 sg13g2_tiehi _30062__385 (.L_HI(net385));
 sg13g2_tiehi _30061__386 (.L_HI(net386));
 sg13g2_tiehi _30060__387 (.L_HI(net387));
 sg13g2_tiehi _30059__388 (.L_HI(net388));
 sg13g2_tiehi _30058__389 (.L_HI(net389));
 sg13g2_tiehi _30057__390 (.L_HI(net390));
 sg13g2_tiehi _30056__391 (.L_HI(net391));
 sg13g2_tiehi _30055__392 (.L_HI(net392));
 sg13g2_tiehi _30054__393 (.L_HI(net393));
 sg13g2_tiehi _30053__394 (.L_HI(net394));
 sg13g2_tiehi _30052__395 (.L_HI(net395));
 sg13g2_tiehi _30051__396 (.L_HI(net396));
 sg13g2_tiehi _30050__397 (.L_HI(net397));
 sg13g2_tiehi _30049__398 (.L_HI(net398));
 sg13g2_tiehi _30048__399 (.L_HI(net399));
 sg13g2_tiehi _30047__400 (.L_HI(net400));
 sg13g2_tiehi _30046__401 (.L_HI(net401));
 sg13g2_tiehi _30045__402 (.L_HI(net402));
 sg13g2_tiehi _30044__403 (.L_HI(net403));
 sg13g2_tiehi _30043__404 (.L_HI(net404));
 sg13g2_tiehi _30042__405 (.L_HI(net405));
 sg13g2_tiehi _30041__406 (.L_HI(net406));
 sg13g2_tiehi _30040__407 (.L_HI(net407));
 sg13g2_tiehi _30039__408 (.L_HI(net408));
 sg13g2_tiehi _30038__409 (.L_HI(net409));
 sg13g2_tiehi _30037__410 (.L_HI(net410));
 sg13g2_tiehi _30036__411 (.L_HI(net411));
 sg13g2_tiehi _30035__412 (.L_HI(net412));
 sg13g2_tiehi _30034__413 (.L_HI(net413));
 sg13g2_tiehi _30033__414 (.L_HI(net414));
 sg13g2_tiehi _30032__415 (.L_HI(net415));
 sg13g2_tiehi _30031__416 (.L_HI(net416));
 sg13g2_tiehi _30030__417 (.L_HI(net417));
 sg13g2_tiehi _30029__418 (.L_HI(net418));
 sg13g2_tiehi _30028__419 (.L_HI(net419));
 sg13g2_tiehi _30027__420 (.L_HI(net420));
 sg13g2_tiehi _30026__421 (.L_HI(net421));
 sg13g2_tiehi _30025__422 (.L_HI(net422));
 sg13g2_tiehi _30024__423 (.L_HI(net423));
 sg13g2_tiehi _30023__424 (.L_HI(net424));
 sg13g2_tiehi _30022__425 (.L_HI(net425));
 sg13g2_tiehi _30021__426 (.L_HI(net426));
 sg13g2_tiehi _30020__427 (.L_HI(net427));
 sg13g2_tiehi _30019__428 (.L_HI(net428));
 sg13g2_tiehi _30018__429 (.L_HI(net429));
 sg13g2_tiehi _30017__430 (.L_HI(net430));
 sg13g2_tiehi _30016__431 (.L_HI(net431));
 sg13g2_tiehi _30015__432 (.L_HI(net432));
 sg13g2_tiehi _30014__433 (.L_HI(net433));
 sg13g2_tiehi _30013__434 (.L_HI(net434));
 sg13g2_tiehi _30012__435 (.L_HI(net435));
 sg13g2_tiehi _30011__436 (.L_HI(net436));
 sg13g2_tiehi _30010__437 (.L_HI(net437));
 sg13g2_tiehi _30009__438 (.L_HI(net438));
 sg13g2_tiehi _30008__439 (.L_HI(net439));
 sg13g2_tiehi _30007__440 (.L_HI(net440));
 sg13g2_tiehi _30006__441 (.L_HI(net441));
 sg13g2_tiehi _30005__442 (.L_HI(net442));
 sg13g2_tiehi _30004__443 (.L_HI(net443));
 sg13g2_tiehi _30003__444 (.L_HI(net444));
 sg13g2_tiehi _30002__445 (.L_HI(net445));
 sg13g2_tiehi _30001__446 (.L_HI(net446));
 sg13g2_tiehi _30000__447 (.L_HI(net447));
 sg13g2_tiehi _29999__448 (.L_HI(net448));
 sg13g2_tiehi _29998__449 (.L_HI(net449));
 sg13g2_tiehi _29997__450 (.L_HI(net450));
 sg13g2_tiehi _29996__451 (.L_HI(net451));
 sg13g2_tiehi _29995__452 (.L_HI(net452));
 sg13g2_tiehi _29994__453 (.L_HI(net453));
 sg13g2_tiehi _29993__454 (.L_HI(net454));
 sg13g2_tiehi _29992__455 (.L_HI(net455));
 sg13g2_tiehi _29991__456 (.L_HI(net456));
 sg13g2_tiehi _29990__457 (.L_HI(net457));
 sg13g2_tiehi _29989__458 (.L_HI(net458));
 sg13g2_tiehi _29988__459 (.L_HI(net459));
 sg13g2_tiehi _29987__460 (.L_HI(net460));
 sg13g2_tiehi _29986__461 (.L_HI(net461));
 sg13g2_tiehi _29985__462 (.L_HI(net462));
 sg13g2_tiehi _29984__463 (.L_HI(net463));
 sg13g2_tiehi _29983__464 (.L_HI(net464));
 sg13g2_tiehi _29982__465 (.L_HI(net465));
 sg13g2_tiehi _29981__466 (.L_HI(net466));
 sg13g2_tiehi _29980__467 (.L_HI(net467));
 sg13g2_tiehi _29979__468 (.L_HI(net468));
 sg13g2_tiehi _29978__469 (.L_HI(net469));
 sg13g2_tiehi _29977__470 (.L_HI(net470));
 sg13g2_tiehi _29976__471 (.L_HI(net471));
 sg13g2_tiehi _29975__472 (.L_HI(net472));
 sg13g2_tiehi _29974__473 (.L_HI(net473));
 sg13g2_tiehi _29973__474 (.L_HI(net474));
 sg13g2_tiehi _29972__475 (.L_HI(net475));
 sg13g2_tiehi _29971__476 (.L_HI(net476));
 sg13g2_tiehi _29970__477 (.L_HI(net477));
 sg13g2_tiehi _29969__478 (.L_HI(net478));
 sg13g2_tiehi _29968__479 (.L_HI(net479));
 sg13g2_tiehi _29967__480 (.L_HI(net480));
 sg13g2_tiehi _29966__481 (.L_HI(net481));
 sg13g2_tiehi _29965__482 (.L_HI(net482));
 sg13g2_tiehi _29964__483 (.L_HI(net483));
 sg13g2_tiehi _29963__484 (.L_HI(net484));
 sg13g2_tiehi _29962__485 (.L_HI(net485));
 sg13g2_tiehi _29961__486 (.L_HI(net486));
 sg13g2_tiehi _29960__487 (.L_HI(net487));
 sg13g2_tiehi _29959__488 (.L_HI(net488));
 sg13g2_tiehi _29958__489 (.L_HI(net489));
 sg13g2_tiehi _29957__490 (.L_HI(net490));
 sg13g2_tiehi _29956__491 (.L_HI(net491));
 sg13g2_tiehi _29955__492 (.L_HI(net492));
 sg13g2_tiehi _29954__493 (.L_HI(net493));
 sg13g2_tiehi _29953__494 (.L_HI(net494));
 sg13g2_tiehi _29952__495 (.L_HI(net495));
 sg13g2_tiehi _29951__496 (.L_HI(net496));
 sg13g2_tiehi _29950__497 (.L_HI(net497));
 sg13g2_tiehi _29949__498 (.L_HI(net498));
 sg13g2_tiehi _29948__499 (.L_HI(net499));
 sg13g2_tiehi _29947__500 (.L_HI(net500));
 sg13g2_tiehi _29946__501 (.L_HI(net501));
 sg13g2_tiehi _29945__502 (.L_HI(net502));
 sg13g2_tiehi _29944__503 (.L_HI(net503));
 sg13g2_tiehi _29943__504 (.L_HI(net504));
 sg13g2_tiehi _29942__505 (.L_HI(net505));
 sg13g2_tiehi _29941__506 (.L_HI(net506));
 sg13g2_tiehi _29940__507 (.L_HI(net507));
 sg13g2_tiehi _29939__508 (.L_HI(net508));
 sg13g2_tiehi _29938__509 (.L_HI(net509));
 sg13g2_tiehi _29937__510 (.L_HI(net510));
 sg13g2_tiehi _29936__511 (.L_HI(net511));
 sg13g2_tiehi _29935__512 (.L_HI(net512));
 sg13g2_tiehi _29934__513 (.L_HI(net513));
 sg13g2_tiehi _29933__514 (.L_HI(net514));
 sg13g2_tiehi _29932__515 (.L_HI(net515));
 sg13g2_tiehi _29931__516 (.L_HI(net516));
 sg13g2_tiehi _29930__517 (.L_HI(net517));
 sg13g2_tiehi _29929__518 (.L_HI(net518));
 sg13g2_tiehi _29928__519 (.L_HI(net519));
 sg13g2_tiehi _29927__520 (.L_HI(net520));
 sg13g2_tiehi _29926__521 (.L_HI(net521));
 sg13g2_tiehi _29925__522 (.L_HI(net522));
 sg13g2_tiehi _29924__523 (.L_HI(net523));
 sg13g2_tiehi _29923__524 (.L_HI(net524));
 sg13g2_tiehi _29922__525 (.L_HI(net525));
 sg13g2_tiehi _29921__526 (.L_HI(net526));
 sg13g2_tiehi _29920__527 (.L_HI(net527));
 sg13g2_tiehi _29919__528 (.L_HI(net528));
 sg13g2_tiehi _29918__529 (.L_HI(net529));
 sg13g2_tiehi _29917__530 (.L_HI(net530));
 sg13g2_tiehi _29916__531 (.L_HI(net531));
 sg13g2_tiehi _29915__532 (.L_HI(net532));
 sg13g2_tiehi _29914__533 (.L_HI(net533));
 sg13g2_tiehi _29913__534 (.L_HI(net534));
 sg13g2_tiehi _29912__535 (.L_HI(net535));
 sg13g2_tiehi _29911__536 (.L_HI(net536));
 sg13g2_tiehi _29910__537 (.L_HI(net537));
 sg13g2_tiehi _29909__538 (.L_HI(net538));
 sg13g2_tiehi _29908__539 (.L_HI(net539));
 sg13g2_tiehi _29907__540 (.L_HI(net540));
 sg13g2_tiehi _29906__541 (.L_HI(net541));
 sg13g2_tiehi _29905__542 (.L_HI(net542));
 sg13g2_tiehi _29904__543 (.L_HI(net543));
 sg13g2_tiehi _29903__544 (.L_HI(net544));
 sg13g2_tiehi _29902__545 (.L_HI(net545));
 sg13g2_tiehi _29901__546 (.L_HI(net546));
 sg13g2_tiehi _29900__547 (.L_HI(net547));
 sg13g2_tiehi _29899__548 (.L_HI(net548));
 sg13g2_tiehi _29898__549 (.L_HI(net549));
 sg13g2_tiehi _29897__550 (.L_HI(net550));
 sg13g2_tiehi _29896__551 (.L_HI(net551));
 sg13g2_tiehi _29895__552 (.L_HI(net552));
 sg13g2_tiehi _29894__553 (.L_HI(net553));
 sg13g2_tiehi _29893__554 (.L_HI(net554));
 sg13g2_tiehi _29892__555 (.L_HI(net555));
 sg13g2_tiehi _29891__556 (.L_HI(net556));
 sg13g2_tiehi _29890__557 (.L_HI(net557));
 sg13g2_tiehi _29889__558 (.L_HI(net558));
 sg13g2_tiehi _29888__559 (.L_HI(net559));
 sg13g2_tiehi _29887__560 (.L_HI(net560));
 sg13g2_tiehi _29886__561 (.L_HI(net561));
 sg13g2_tiehi _29885__562 (.L_HI(net562));
 sg13g2_tiehi _29884__563 (.L_HI(net563));
 sg13g2_tiehi _29883__564 (.L_HI(net564));
 sg13g2_tiehi _29882__565 (.L_HI(net565));
 sg13g2_tiehi _29881__566 (.L_HI(net566));
 sg13g2_tiehi _29880__567 (.L_HI(net567));
 sg13g2_tiehi _29879__568 (.L_HI(net568));
 sg13g2_tiehi _29878__569 (.L_HI(net569));
 sg13g2_tiehi _29877__570 (.L_HI(net570));
 sg13g2_tiehi _29876__571 (.L_HI(net571));
 sg13g2_tiehi _29875__572 (.L_HI(net572));
 sg13g2_tiehi _29874__573 (.L_HI(net573));
 sg13g2_tiehi _29873__574 (.L_HI(net574));
 sg13g2_tiehi _29872__575 (.L_HI(net575));
 sg13g2_tiehi _29871__576 (.L_HI(net576));
 sg13g2_tiehi _29870__577 (.L_HI(net577));
 sg13g2_tiehi _29869__578 (.L_HI(net578));
 sg13g2_tiehi _29868__579 (.L_HI(net579));
 sg13g2_tiehi _29867__580 (.L_HI(net580));
 sg13g2_tiehi _29866__581 (.L_HI(net581));
 sg13g2_tiehi _29865__582 (.L_HI(net582));
 sg13g2_tiehi _29864__583 (.L_HI(net583));
 sg13g2_tiehi _29863__584 (.L_HI(net584));
 sg13g2_tiehi _29862__585 (.L_HI(net585));
 sg13g2_tiehi _29861__586 (.L_HI(net586));
 sg13g2_tiehi _29860__587 (.L_HI(net587));
 sg13g2_tiehi _29859__588 (.L_HI(net588));
 sg13g2_tiehi _29858__589 (.L_HI(net589));
 sg13g2_tiehi _29857__590 (.L_HI(net590));
 sg13g2_tiehi _29856__591 (.L_HI(net591));
 sg13g2_tiehi _29855__592 (.L_HI(net592));
 sg13g2_tiehi _29854__593 (.L_HI(net593));
 sg13g2_tiehi _29853__594 (.L_HI(net594));
 sg13g2_tiehi _29852__595 (.L_HI(net595));
 sg13g2_tiehi _29851__596 (.L_HI(net596));
 sg13g2_tiehi _29850__597 (.L_HI(net597));
 sg13g2_tiehi _29849__598 (.L_HI(net598));
 sg13g2_tiehi _29848__599 (.L_HI(net599));
 sg13g2_tiehi _29847__600 (.L_HI(net600));
 sg13g2_tiehi _29846__601 (.L_HI(net601));
 sg13g2_tiehi _29845__602 (.L_HI(net602));
 sg13g2_tiehi _29844__603 (.L_HI(net603));
 sg13g2_tiehi _29843__604 (.L_HI(net604));
 sg13g2_tiehi _29842__605 (.L_HI(net605));
 sg13g2_tiehi _29841__606 (.L_HI(net606));
 sg13g2_tiehi _29840__607 (.L_HI(net607));
 sg13g2_tiehi _29839__608 (.L_HI(net608));
 sg13g2_tiehi _29838__609 (.L_HI(net609));
 sg13g2_tiehi _29837__610 (.L_HI(net610));
 sg13g2_tiehi _29836__611 (.L_HI(net611));
 sg13g2_tiehi _29835__612 (.L_HI(net612));
 sg13g2_tiehi _29834__613 (.L_HI(net613));
 sg13g2_tiehi _29833__614 (.L_HI(net614));
 sg13g2_tiehi _29832__615 (.L_HI(net615));
 sg13g2_tiehi _29831__616 (.L_HI(net616));
 sg13g2_tiehi _29830__617 (.L_HI(net617));
 sg13g2_tiehi _29829__618 (.L_HI(net618));
 sg13g2_tiehi _29828__619 (.L_HI(net619));
 sg13g2_tiehi _29827__620 (.L_HI(net620));
 sg13g2_tiehi _29826__621 (.L_HI(net621));
 sg13g2_tiehi _29825__622 (.L_HI(net622));
 sg13g2_tiehi _29824__623 (.L_HI(net623));
 sg13g2_tiehi _29823__624 (.L_HI(net624));
 sg13g2_tiehi _29822__625 (.L_HI(net625));
 sg13g2_tiehi _29821__626 (.L_HI(net626));
 sg13g2_tiehi _29820__627 (.L_HI(net627));
 sg13g2_tiehi _29819__628 (.L_HI(net628));
 sg13g2_tiehi _29818__629 (.L_HI(net629));
 sg13g2_tiehi _29817__630 (.L_HI(net630));
 sg13g2_tiehi _29816__631 (.L_HI(net631));
 sg13g2_tiehi _29815__632 (.L_HI(net632));
 sg13g2_tiehi _29814__633 (.L_HI(net633));
 sg13g2_tiehi _29813__634 (.L_HI(net634));
 sg13g2_tiehi _29812__635 (.L_HI(net635));
 sg13g2_tiehi _29811__636 (.L_HI(net636));
 sg13g2_tiehi _29810__637 (.L_HI(net637));
 sg13g2_tiehi _29809__638 (.L_HI(net638));
 sg13g2_tiehi _29808__639 (.L_HI(net639));
 sg13g2_tiehi _29807__640 (.L_HI(net640));
 sg13g2_tiehi _29806__641 (.L_HI(net641));
 sg13g2_tiehi _29805__642 (.L_HI(net642));
 sg13g2_tiehi _29804__643 (.L_HI(net643));
 sg13g2_tiehi _29803__644 (.L_HI(net644));
 sg13g2_tiehi _29802__645 (.L_HI(net645));
 sg13g2_tiehi _29801__646 (.L_HI(net646));
 sg13g2_tiehi _29800__647 (.L_HI(net647));
 sg13g2_tiehi _29799__648 (.L_HI(net648));
 sg13g2_tiehi _29798__649 (.L_HI(net649));
 sg13g2_tiehi _29797__650 (.L_HI(net650));
 sg13g2_tiehi _29796__651 (.L_HI(net651));
 sg13g2_tiehi _29795__652 (.L_HI(net652));
 sg13g2_tiehi _29794__653 (.L_HI(net653));
 sg13g2_tiehi _29793__654 (.L_HI(net654));
 sg13g2_tiehi _29792__655 (.L_HI(net655));
 sg13g2_tiehi _29791__656 (.L_HI(net656));
 sg13g2_tiehi _29790__657 (.L_HI(net657));
 sg13g2_tiehi _29789__658 (.L_HI(net658));
 sg13g2_tiehi _29788__659 (.L_HI(net659));
 sg13g2_tiehi _29787__660 (.L_HI(net660));
 sg13g2_tiehi _29786__661 (.L_HI(net661));
 sg13g2_tiehi _29785__662 (.L_HI(net662));
 sg13g2_tiehi _29784__663 (.L_HI(net663));
 sg13g2_tiehi _29783__664 (.L_HI(net664));
 sg13g2_tiehi _29782__665 (.L_HI(net665));
 sg13g2_tiehi _29781__666 (.L_HI(net666));
 sg13g2_tiehi _29780__667 (.L_HI(net667));
 sg13g2_tiehi _29779__668 (.L_HI(net668));
 sg13g2_tiehi _29778__669 (.L_HI(net669));
 sg13g2_tiehi _29777__670 (.L_HI(net670));
 sg13g2_tiehi _29776__671 (.L_HI(net671));
 sg13g2_tiehi _29775__672 (.L_HI(net672));
 sg13g2_tiehi _29774__673 (.L_HI(net673));
 sg13g2_tiehi _29773__674 (.L_HI(net674));
 sg13g2_tiehi _29772__675 (.L_HI(net675));
 sg13g2_tiehi _29771__676 (.L_HI(net676));
 sg13g2_tiehi _29770__677 (.L_HI(net677));
 sg13g2_tiehi _29769__678 (.L_HI(net678));
 sg13g2_tiehi _29768__679 (.L_HI(net679));
 sg13g2_tiehi _29767__680 (.L_HI(net680));
 sg13g2_tiehi _29766__681 (.L_HI(net681));
 sg13g2_tiehi _29765__682 (.L_HI(net682));
 sg13g2_tiehi _29764__683 (.L_HI(net683));
 sg13g2_tiehi _29763__684 (.L_HI(net684));
 sg13g2_tiehi _29762__685 (.L_HI(net685));
 sg13g2_tiehi _29761__686 (.L_HI(net686));
 sg13g2_tiehi _29760__687 (.L_HI(net687));
 sg13g2_tiehi _29759__688 (.L_HI(net688));
 sg13g2_tiehi _29758__689 (.L_HI(net689));
 sg13g2_tiehi _29757__690 (.L_HI(net690));
 sg13g2_tiehi _29756__691 (.L_HI(net691));
 sg13g2_tiehi _29755__692 (.L_HI(net692));
 sg13g2_tiehi _29754__693 (.L_HI(net693));
 sg13g2_tiehi _29753__694 (.L_HI(net694));
 sg13g2_tiehi _29752__695 (.L_HI(net695));
 sg13g2_tiehi _29751__696 (.L_HI(net696));
 sg13g2_tiehi _29750__697 (.L_HI(net697));
 sg13g2_tiehi _29749__698 (.L_HI(net698));
 sg13g2_tiehi _29748__699 (.L_HI(net699));
 sg13g2_tiehi _29747__700 (.L_HI(net700));
 sg13g2_tiehi _29746__701 (.L_HI(net701));
 sg13g2_tiehi _29745__702 (.L_HI(net702));
 sg13g2_tiehi _29744__703 (.L_HI(net703));
 sg13g2_tiehi _29743__704 (.L_HI(net704));
 sg13g2_tiehi _29742__705 (.L_HI(net705));
 sg13g2_tiehi _29741__706 (.L_HI(net706));
 sg13g2_tiehi _29740__707 (.L_HI(net707));
 sg13g2_tiehi _29739__708 (.L_HI(net708));
 sg13g2_tiehi _29738__709 (.L_HI(net709));
 sg13g2_tiehi _29737__710 (.L_HI(net710));
 sg13g2_tiehi _29736__711 (.L_HI(net711));
 sg13g2_tiehi _29735__712 (.L_HI(net712));
 sg13g2_tiehi _29734__713 (.L_HI(net713));
 sg13g2_tiehi _29733__714 (.L_HI(net714));
 sg13g2_tiehi _29732__715 (.L_HI(net715));
 sg13g2_tiehi _29731__716 (.L_HI(net716));
 sg13g2_tiehi _29730__717 (.L_HI(net717));
 sg13g2_tiehi _29729__718 (.L_HI(net718));
 sg13g2_tiehi _29728__719 (.L_HI(net719));
 sg13g2_tiehi _29727__720 (.L_HI(net720));
 sg13g2_tiehi _29726__721 (.L_HI(net721));
 sg13g2_tiehi _29725__722 (.L_HI(net722));
 sg13g2_tiehi _29724__723 (.L_HI(net723));
 sg13g2_tiehi _29723__724 (.L_HI(net724));
 sg13g2_tiehi _29722__725 (.L_HI(net725));
 sg13g2_tiehi _29721__726 (.L_HI(net726));
 sg13g2_tiehi _29720__727 (.L_HI(net727));
 sg13g2_tiehi _29719__728 (.L_HI(net728));
 sg13g2_tiehi _29718__729 (.L_HI(net729));
 sg13g2_tiehi _29717__730 (.L_HI(net730));
 sg13g2_tiehi _29716__731 (.L_HI(net731));
 sg13g2_tiehi _29715__732 (.L_HI(net732));
 sg13g2_tiehi _29714__733 (.L_HI(net733));
 sg13g2_tiehi _29713__734 (.L_HI(net734));
 sg13g2_tiehi _29712__735 (.L_HI(net735));
 sg13g2_tiehi _29711__736 (.L_HI(net736));
 sg13g2_tiehi _29710__737 (.L_HI(net737));
 sg13g2_tiehi _29709__738 (.L_HI(net738));
 sg13g2_tiehi _29708__739 (.L_HI(net739));
 sg13g2_tiehi _29707__740 (.L_HI(net740));
 sg13g2_tiehi _29706__741 (.L_HI(net741));
 sg13g2_tiehi _29705__742 (.L_HI(net742));
 sg13g2_tiehi _29704__743 (.L_HI(net743));
 sg13g2_tiehi _29703__744 (.L_HI(net744));
 sg13g2_tiehi _29702__745 (.L_HI(net745));
 sg13g2_tiehi _29701__746 (.L_HI(net746));
 sg13g2_tiehi _29700__747 (.L_HI(net747));
 sg13g2_tiehi _29699__748 (.L_HI(net748));
 sg13g2_tiehi _29698__749 (.L_HI(net749));
 sg13g2_tiehi _29697__750 (.L_HI(net750));
 sg13g2_tiehi _29696__751 (.L_HI(net751));
 sg13g2_tiehi _29695__752 (.L_HI(net752));
 sg13g2_tiehi _29694__753 (.L_HI(net753));
 sg13g2_tiehi _29693__754 (.L_HI(net754));
 sg13g2_tiehi _29692__755 (.L_HI(net755));
 sg13g2_tiehi _29691__756 (.L_HI(net756));
 sg13g2_tiehi _29690__757 (.L_HI(net757));
 sg13g2_tiehi _29689__758 (.L_HI(net758));
 sg13g2_tiehi _29688__759 (.L_HI(net759));
 sg13g2_tiehi _29687__760 (.L_HI(net760));
 sg13g2_tiehi _29686__761 (.L_HI(net761));
 sg13g2_tiehi _29685__762 (.L_HI(net762));
 sg13g2_tiehi _29684__763 (.L_HI(net763));
 sg13g2_tiehi _29683__764 (.L_HI(net764));
 sg13g2_tiehi _29682__765 (.L_HI(net765));
 sg13g2_tiehi _29681__766 (.L_HI(net766));
 sg13g2_tiehi _29680__767 (.L_HI(net767));
 sg13g2_tiehi _29679__768 (.L_HI(net768));
 sg13g2_tiehi _29678__769 (.L_HI(net769));
 sg13g2_tiehi _29677__770 (.L_HI(net770));
 sg13g2_tiehi _29676__771 (.L_HI(net771));
 sg13g2_tiehi _29675__772 (.L_HI(net772));
 sg13g2_tiehi _29674__773 (.L_HI(net773));
 sg13g2_tiehi _29673__774 (.L_HI(net774));
 sg13g2_tiehi _29672__775 (.L_HI(net775));
 sg13g2_tiehi _29671__776 (.L_HI(net776));
 sg13g2_tiehi _29670__777 (.L_HI(net777));
 sg13g2_tiehi _29669__778 (.L_HI(net778));
 sg13g2_tiehi _29668__779 (.L_HI(net779));
 sg13g2_tiehi _29667__780 (.L_HI(net780));
 sg13g2_tiehi _29666__781 (.L_HI(net781));
 sg13g2_tiehi _29665__782 (.L_HI(net782));
 sg13g2_tiehi _29664__783 (.L_HI(net783));
 sg13g2_tiehi _29663__784 (.L_HI(net784));
 sg13g2_tiehi _29662__785 (.L_HI(net785));
 sg13g2_tiehi _29661__786 (.L_HI(net786));
 sg13g2_tiehi _29660__787 (.L_HI(net787));
 sg13g2_tiehi _29659__788 (.L_HI(net788));
 sg13g2_tiehi _29658__789 (.L_HI(net789));
 sg13g2_tiehi _29657__790 (.L_HI(net790));
 sg13g2_tiehi _29656__791 (.L_HI(net791));
 sg13g2_tiehi _29655__792 (.L_HI(net792));
 sg13g2_tiehi _29654__793 (.L_HI(net793));
 sg13g2_tiehi _29653__794 (.L_HI(net794));
 sg13g2_tiehi _29652__795 (.L_HI(net795));
 sg13g2_tiehi _29651__796 (.L_HI(net796));
 sg13g2_tiehi _29650__797 (.L_HI(net797));
 sg13g2_tiehi _29649__798 (.L_HI(net798));
 sg13g2_tiehi _29648__799 (.L_HI(net799));
 sg13g2_tiehi _29647__800 (.L_HI(net800));
 sg13g2_tiehi _29646__801 (.L_HI(net801));
 sg13g2_tiehi _29645__802 (.L_HI(net802));
 sg13g2_tiehi _29644__803 (.L_HI(net803));
 sg13g2_tiehi _29643__804 (.L_HI(net804));
 sg13g2_tiehi _28072__805 (.L_HI(net805));
 sg13g2_tiehi _28640__806 (.L_HI(net806));
 sg13g2_tiehi _28641__807 (.L_HI(net807));
 sg13g2_tiehi _28642__808 (.L_HI(net808));
 sg13g2_tiehi _28643__809 (.L_HI(net809));
 sg13g2_tiehi _28644__810 (.L_HI(net810));
 sg13g2_tiehi _28645__811 (.L_HI(net811));
 sg13g2_tiehi _28646__812 (.L_HI(net812));
 sg13g2_tiehi _28647__813 (.L_HI(net813));
 sg13g2_tiehi _28648__814 (.L_HI(net814));
 sg13g2_tiehi _28649__815 (.L_HI(net815));
 sg13g2_tiehi _28650__816 (.L_HI(net816));
 sg13g2_tiehi _28651__817 (.L_HI(net817));
 sg13g2_tiehi _28652__818 (.L_HI(net818));
 sg13g2_tiehi _28653__819 (.L_HI(net819));
 sg13g2_tiehi _28654__820 (.L_HI(net820));
 sg13g2_tiehi _28655__821 (.L_HI(net821));
 sg13g2_tiehi _29642__822 (.L_HI(net822));
 sg13g2_tiehi _29641__823 (.L_HI(net823));
 sg13g2_tiehi _29640__824 (.L_HI(net824));
 sg13g2_tiehi _29639__825 (.L_HI(net825));
 sg13g2_tiehi _29638__826 (.L_HI(net826));
 sg13g2_tiehi _29637__827 (.L_HI(net827));
 sg13g2_tiehi _29636__828 (.L_HI(net828));
 sg13g2_tiehi _29635__829 (.L_HI(net829));
 sg13g2_tiehi _29634__830 (.L_HI(net830));
 sg13g2_tiehi _29633__831 (.L_HI(net831));
 sg13g2_tiehi _29632__832 (.L_HI(net832));
 sg13g2_tiehi _29631__833 (.L_HI(net833));
 sg13g2_tiehi _29630__834 (.L_HI(net834));
 sg13g2_tiehi _29629__835 (.L_HI(net835));
 sg13g2_tiehi _29628__836 (.L_HI(net836));
 sg13g2_tiehi _29627__837 (.L_HI(net837));
 sg13g2_tiehi _29626__838 (.L_HI(net838));
 sg13g2_tiehi _29625__839 (.L_HI(net839));
 sg13g2_tiehi _29624__840 (.L_HI(net840));
 sg13g2_tiehi _29623__841 (.L_HI(net841));
 sg13g2_tiehi _29622__842 (.L_HI(net842));
 sg13g2_tiehi _29621__843 (.L_HI(net843));
 sg13g2_tiehi _29620__844 (.L_HI(net844));
 sg13g2_tiehi _29619__845 (.L_HI(net845));
 sg13g2_tiehi _29618__846 (.L_HI(net846));
 sg13g2_tiehi _29617__847 (.L_HI(net847));
 sg13g2_tiehi _29616__848 (.L_HI(net848));
 sg13g2_tiehi _29615__849 (.L_HI(net849));
 sg13g2_tiehi _29614__850 (.L_HI(net850));
 sg13g2_tiehi _29613__851 (.L_HI(net851));
 sg13g2_tiehi _29612__852 (.L_HI(net852));
 sg13g2_tiehi _29611__853 (.L_HI(net853));
 sg13g2_tiehi _29610__854 (.L_HI(net854));
 sg13g2_tiehi _29609__855 (.L_HI(net855));
 sg13g2_tiehi _29608__856 (.L_HI(net856));
 sg13g2_tiehi _29607__857 (.L_HI(net857));
 sg13g2_tiehi _29606__858 (.L_HI(net858));
 sg13g2_tiehi _29605__859 (.L_HI(net859));
 sg13g2_tiehi _29604__860 (.L_HI(net860));
 sg13g2_tiehi _29603__861 (.L_HI(net861));
 sg13g2_tiehi _29602__862 (.L_HI(net862));
 sg13g2_tiehi _29601__863 (.L_HI(net863));
 sg13g2_tiehi _29600__864 (.L_HI(net864));
 sg13g2_tiehi _29599__865 (.L_HI(net865));
 sg13g2_tiehi _29598__866 (.L_HI(net866));
 sg13g2_tiehi _29597__867 (.L_HI(net867));
 sg13g2_tiehi _29596__868 (.L_HI(net868));
 sg13g2_tiehi _29595__869 (.L_HI(net869));
 sg13g2_tiehi _29594__870 (.L_HI(net870));
 sg13g2_tiehi _29593__871 (.L_HI(net871));
 sg13g2_tiehi _29592__872 (.L_HI(net872));
 sg13g2_tiehi _29591__873 (.L_HI(net873));
 sg13g2_tiehi _29590__874 (.L_HI(net874));
 sg13g2_tiehi _29589__875 (.L_HI(net875));
 sg13g2_tiehi _29588__876 (.L_HI(net876));
 sg13g2_tiehi _29587__877 (.L_HI(net877));
 sg13g2_tiehi _29586__878 (.L_HI(net878));
 sg13g2_tiehi _29585__879 (.L_HI(net879));
 sg13g2_tiehi _29584__880 (.L_HI(net880));
 sg13g2_tiehi _29583__881 (.L_HI(net881));
 sg13g2_tiehi _29582__882 (.L_HI(net882));
 sg13g2_tiehi _29581__883 (.L_HI(net883));
 sg13g2_tiehi _29580__884 (.L_HI(net884));
 sg13g2_tiehi _29579__885 (.L_HI(net885));
 sg13g2_tiehi _29578__886 (.L_HI(net886));
 sg13g2_tiehi _29577__887 (.L_HI(net887));
 sg13g2_tiehi _29576__888 (.L_HI(net888));
 sg13g2_tiehi _29575__889 (.L_HI(net889));
 sg13g2_tiehi _29574__890 (.L_HI(net890));
 sg13g2_tiehi _29573__891 (.L_HI(net891));
 sg13g2_tiehi _29572__892 (.L_HI(net892));
 sg13g2_tiehi _29571__893 (.L_HI(net893));
 sg13g2_tiehi _29570__894 (.L_HI(net894));
 sg13g2_tiehi _29569__895 (.L_HI(net895));
 sg13g2_tiehi _29568__896 (.L_HI(net896));
 sg13g2_tiehi _29567__897 (.L_HI(net897));
 sg13g2_tiehi _29566__898 (.L_HI(net898));
 sg13g2_tiehi _29565__899 (.L_HI(net899));
 sg13g2_tiehi _29564__900 (.L_HI(net900));
 sg13g2_tiehi _29563__901 (.L_HI(net901));
 sg13g2_tiehi _29562__902 (.L_HI(net902));
 sg13g2_tiehi _29561__903 (.L_HI(net903));
 sg13g2_tiehi _29560__904 (.L_HI(net904));
 sg13g2_tiehi _29559__905 (.L_HI(net905));
 sg13g2_tiehi _29558__906 (.L_HI(net906));
 sg13g2_tiehi _29557__907 (.L_HI(net907));
 sg13g2_tiehi _29556__908 (.L_HI(net908));
 sg13g2_tiehi _29555__909 (.L_HI(net909));
 sg13g2_tiehi _29554__910 (.L_HI(net910));
 sg13g2_tiehi _29553__911 (.L_HI(net911));
 sg13g2_tiehi _29552__912 (.L_HI(net912));
 sg13g2_tiehi _29551__913 (.L_HI(net913));
 sg13g2_tiehi _29550__914 (.L_HI(net914));
 sg13g2_tiehi _29549__915 (.L_HI(net915));
 sg13g2_tiehi _29548__916 (.L_HI(net916));
 sg13g2_tiehi _29547__917 (.L_HI(net917));
 sg13g2_tiehi _29546__918 (.L_HI(net918));
 sg13g2_tiehi _29545__919 (.L_HI(net919));
 sg13g2_tiehi _29544__920 (.L_HI(net920));
 sg13g2_tiehi _29543__921 (.L_HI(net921));
 sg13g2_tiehi _29542__922 (.L_HI(net922));
 sg13g2_tiehi _29541__923 (.L_HI(net923));
 sg13g2_tiehi _29540__924 (.L_HI(net924));
 sg13g2_tiehi _29539__925 (.L_HI(net925));
 sg13g2_tiehi _29538__926 (.L_HI(net926));
 sg13g2_tiehi _29537__927 (.L_HI(net927));
 sg13g2_tiehi _29536__928 (.L_HI(net928));
 sg13g2_tiehi _29535__929 (.L_HI(net929));
 sg13g2_tiehi _29534__930 (.L_HI(net930));
 sg13g2_tiehi _29533__931 (.L_HI(net931));
 sg13g2_tiehi _29532__932 (.L_HI(net932));
 sg13g2_tiehi _29531__933 (.L_HI(net933));
 sg13g2_tiehi _29530__934 (.L_HI(net934));
 sg13g2_tiehi _29529__935 (.L_HI(net935));
 sg13g2_tiehi _29528__936 (.L_HI(net936));
 sg13g2_tiehi _29527__937 (.L_HI(net937));
 sg13g2_tiehi _29526__938 (.L_HI(net938));
 sg13g2_tiehi _29525__939 (.L_HI(net939));
 sg13g2_tiehi _29524__940 (.L_HI(net940));
 sg13g2_tiehi _29523__941 (.L_HI(net941));
 sg13g2_tiehi _29522__942 (.L_HI(net942));
 sg13g2_tiehi _29521__943 (.L_HI(net943));
 sg13g2_tiehi _29520__944 (.L_HI(net944));
 sg13g2_tiehi _29519__945 (.L_HI(net945));
 sg13g2_tiehi _29518__946 (.L_HI(net946));
 sg13g2_tiehi _29517__947 (.L_HI(net947));
 sg13g2_tiehi _29516__948 (.L_HI(net948));
 sg13g2_tiehi _29515__949 (.L_HI(net949));
 sg13g2_tiehi _29514__950 (.L_HI(net950));
 sg13g2_tiehi _29513__951 (.L_HI(net951));
 sg13g2_tiehi _29512__952 (.L_HI(net952));
 sg13g2_tiehi _29511__953 (.L_HI(net953));
 sg13g2_tiehi _29510__954 (.L_HI(net954));
 sg13g2_tiehi _29509__955 (.L_HI(net955));
 sg13g2_tiehi _29508__956 (.L_HI(net956));
 sg13g2_tiehi _29507__957 (.L_HI(net957));
 sg13g2_tiehi _29506__958 (.L_HI(net958));
 sg13g2_tiehi _29505__959 (.L_HI(net959));
 sg13g2_tiehi _29504__960 (.L_HI(net960));
 sg13g2_tiehi _29503__961 (.L_HI(net961));
 sg13g2_tiehi _29502__962 (.L_HI(net962));
 sg13g2_tiehi _29501__963 (.L_HI(net963));
 sg13g2_tiehi _28656__964 (.L_HI(net964));
 sg13g2_tiehi _28799__965 (.L_HI(net965));
 sg13g2_tiehi _28800__966 (.L_HI(net966));
 sg13g2_tiehi _28801__967 (.L_HI(net967));
 sg13g2_tiehi _28802__968 (.L_HI(net968));
 sg13g2_tiehi _28803__969 (.L_HI(net969));
 sg13g2_tiehi _28804__970 (.L_HI(net970));
 sg13g2_tiehi _28805__971 (.L_HI(net971));
 sg13g2_tiehi _28806__972 (.L_HI(net972));
 sg13g2_tiehi _28807__973 (.L_HI(net973));
 sg13g2_tiehi _28808__974 (.L_HI(net974));
 sg13g2_tiehi _28809__975 (.L_HI(net975));
 sg13g2_tiehi _28810__976 (.L_HI(net976));
 sg13g2_tiehi _28811__977 (.L_HI(net977));
 sg13g2_tiehi _28812__978 (.L_HI(net978));
 sg13g2_tiehi _30686__979 (.L_HI(net979));
 sg13g2_tiehi _29500__980 (.L_HI(net980));
 sg13g2_tiehi _30690__981 (.L_HI(net981));
 sg13g2_tiehi _29499__982 (.L_HI(net982));
 sg13g2_tiehi _30685__983 (.L_HI(net983));
 sg13g2_tiehi _29498__984 (.L_HI(net984));
 sg13g2_tiehi _30688__985 (.L_HI(net985));
 sg13g2_tiehi _29497__986 (.L_HI(net986));
 sg13g2_tiehi _30684__987 (.L_HI(net987));
 sg13g2_tiehi _29496__988 (.L_HI(net988));
 sg13g2_tiehi _29479__989 (.L_HI(net989));
 sg13g2_tiehi _29495__990 (.L_HI(net990));
 sg13g2_tiehi _29494__991 (.L_HI(net991));
 sg13g2_tiehi _29493__992 (.L_HI(net992));
 sg13g2_tiehi _29492__993 (.L_HI(net993));
 sg13g2_tiehi _29491__994 (.L_HI(net994));
 sg13g2_tiehi _29490__995 (.L_HI(net995));
 sg13g2_tiehi _29489__996 (.L_HI(net996));
 sg13g2_tiehi _29488__997 (.L_HI(net997));
 sg13g2_tiehi _29487__998 (.L_HI(net998));
 sg13g2_tiehi _30683__999 (.L_HI(net999));
 sg13g2_tiehi _29486__1000 (.L_HI(net1000));
 sg13g2_tiehi _30687__1001 (.L_HI(net1001));
 sg13g2_tiehi _29485__1002 (.L_HI(net1002));
 sg13g2_tiehi _30682__1003 (.L_HI(net1003));
 sg13g2_tiehi _29484__1004 (.L_HI(net1004));
 sg13g2_tiehi _30689__1005 (.L_HI(net1005));
 sg13g2_tiehi _29483__1006 (.L_HI(net1006));
 sg13g2_tiehi _30681__1007 (.L_HI(net1007));
 sg13g2_tiehi _29482__1008 (.L_HI(net1008));
 sg13g2_tiehi _29481__1009 (.L_HI(net1009));
 sg13g2_tiehi _29480__1010 (.L_HI(net1010));
 sg13g2_tiehi _29471__1011 (.L_HI(net1011));
 sg13g2_tiehi _29470__1012 (.L_HI(net1012));
 sg13g2_tiehi _29469__1013 (.L_HI(net1013));
 sg13g2_tiehi _29468__1014 (.L_HI(net1014));
 sg13g2_tiehi _29467__1015 (.L_HI(net1015));
 sg13g2_tiehi _29466__1016 (.L_HI(net1016));
 sg13g2_tiehi _29465__1017 (.L_HI(net1017));
 sg13g2_tiehi _29464__1018 (.L_HI(net1018));
 sg13g2_tiehi _29463__1019 (.L_HI(net1019));
 sg13g2_tiehi _29462__1020 (.L_HI(net1020));
 sg13g2_tiehi _29461__1021 (.L_HI(net1021));
 sg13g2_tiehi _29460__1022 (.L_HI(net1022));
 sg13g2_tiehi _29459__1023 (.L_HI(net1023));
 sg13g2_tiehi _29458__1024 (.L_HI(net1024));
 sg13g2_tiehi _29457__1025 (.L_HI(net1025));
 sg13g2_tiehi _29456__1026 (.L_HI(net1026));
 sg13g2_tiehi _29455__1027 (.L_HI(net1027));
 sg13g2_tiehi _29454__1028 (.L_HI(net1028));
 sg13g2_tiehi _29453__1029 (.L_HI(net1029));
 sg13g2_tiehi _29452__1030 (.L_HI(net1030));
 sg13g2_tiehi _29451__1031 (.L_HI(net1031));
 sg13g2_tiehi _29450__1032 (.L_HI(net1032));
 sg13g2_tiehi _29449__1033 (.L_HI(net1033));
 sg13g2_tiehi _29448__1034 (.L_HI(net1034));
 sg13g2_tiehi _29447__1035 (.L_HI(net1035));
 sg13g2_tiehi _29446__1036 (.L_HI(net1036));
 sg13g2_tiehi _29445__1037 (.L_HI(net1037));
 sg13g2_tiehi _29444__1038 (.L_HI(net1038));
 sg13g2_tiehi _29443__1039 (.L_HI(net1039));
 sg13g2_tiehi _29442__1040 (.L_HI(net1040));
 sg13g2_tiehi _29441__1041 (.L_HI(net1041));
 sg13g2_tiehi _29440__1042 (.L_HI(net1042));
 sg13g2_tiehi _29439__1043 (.L_HI(net1043));
 sg13g2_tiehi _29438__1044 (.L_HI(net1044));
 sg13g2_tiehi _29437__1045 (.L_HI(net1045));
 sg13g2_tiehi _29436__1046 (.L_HI(net1046));
 sg13g2_tiehi _29435__1047 (.L_HI(net1047));
 sg13g2_tiehi _29434__1048 (.L_HI(net1048));
 sg13g2_tiehi _29433__1049 (.L_HI(net1049));
 sg13g2_tiehi _29432__1050 (.L_HI(net1050));
 sg13g2_tiehi _29431__1051 (.L_HI(net1051));
 sg13g2_tiehi _29430__1052 (.L_HI(net1052));
 sg13g2_tiehi _29429__1053 (.L_HI(net1053));
 sg13g2_tiehi _29428__1054 (.L_HI(net1054));
 sg13g2_tiehi _29427__1055 (.L_HI(net1055));
 sg13g2_tiehi _29426__1056 (.L_HI(net1056));
 sg13g2_tiehi _29425__1057 (.L_HI(net1057));
 sg13g2_tiehi _29424__1058 (.L_HI(net1058));
 sg13g2_tiehi _29423__1059 (.L_HI(net1059));
 sg13g2_tiehi _29422__1060 (.L_HI(net1060));
 sg13g2_tiehi _29421__1061 (.L_HI(net1061));
 sg13g2_tiehi _29420__1062 (.L_HI(net1062));
 sg13g2_tiehi _29419__1063 (.L_HI(net1063));
 sg13g2_tiehi _29418__1064 (.L_HI(net1064));
 sg13g2_tiehi _29417__1065 (.L_HI(net1065));
 sg13g2_tiehi _29416__1066 (.L_HI(net1066));
 sg13g2_tiehi _29415__1067 (.L_HI(net1067));
 sg13g2_tiehi _29414__1068 (.L_HI(net1068));
 sg13g2_tiehi _29413__1069 (.L_HI(net1069));
 sg13g2_tiehi _29412__1070 (.L_HI(net1070));
 sg13g2_tiehi _29411__1071 (.L_HI(net1071));
 sg13g2_tiehi _29410__1072 (.L_HI(net1072));
 sg13g2_tiehi _29409__1073 (.L_HI(net1073));
 sg13g2_tiehi _29408__1074 (.L_HI(net1074));
 sg13g2_tiehi _29407__1075 (.L_HI(net1075));
 sg13g2_tiehi _29406__1076 (.L_HI(net1076));
 sg13g2_tiehi _29405__1077 (.L_HI(net1077));
 sg13g2_tiehi _29404__1078 (.L_HI(net1078));
 sg13g2_tiehi _29403__1079 (.L_HI(net1079));
 sg13g2_tiehi _29402__1080 (.L_HI(net1080));
 sg13g2_tiehi _29401__1081 (.L_HI(net1081));
 sg13g2_tiehi _29400__1082 (.L_HI(net1082));
 sg13g2_tiehi _29399__1083 (.L_HI(net1083));
 sg13g2_tiehi _29398__1084 (.L_HI(net1084));
 sg13g2_tiehi _29397__1085 (.L_HI(net1085));
 sg13g2_tiehi _29396__1086 (.L_HI(net1086));
 sg13g2_tiehi _29395__1087 (.L_HI(net1087));
 sg13g2_tiehi _29394__1088 (.L_HI(net1088));
 sg13g2_tiehi _29393__1089 (.L_HI(net1089));
 sg13g2_tiehi _29392__1090 (.L_HI(net1090));
 sg13g2_tiehi _29391__1091 (.L_HI(net1091));
 sg13g2_tiehi _29390__1092 (.L_HI(net1092));
 sg13g2_tiehi _29389__1093 (.L_HI(net1093));
 sg13g2_tiehi _29388__1094 (.L_HI(net1094));
 sg13g2_tiehi _29387__1095 (.L_HI(net1095));
 sg13g2_tiehi _29386__1096 (.L_HI(net1096));
 sg13g2_tiehi _29385__1097 (.L_HI(net1097));
 sg13g2_tiehi _29384__1098 (.L_HI(net1098));
 sg13g2_tiehi _29383__1099 (.L_HI(net1099));
 sg13g2_tiehi _29382__1100 (.L_HI(net1100));
 sg13g2_tiehi _29381__1101 (.L_HI(net1101));
 sg13g2_tiehi _29380__1102 (.L_HI(net1102));
 sg13g2_tiehi _29379__1103 (.L_HI(net1103));
 sg13g2_tiehi _29378__1104 (.L_HI(net1104));
 sg13g2_tiehi _29377__1105 (.L_HI(net1105));
 sg13g2_tiehi _29376__1106 (.L_HI(net1106));
 sg13g2_tiehi _29375__1107 (.L_HI(net1107));
 sg13g2_tiehi _29374__1108 (.L_HI(net1108));
 sg13g2_tiehi _29373__1109 (.L_HI(net1109));
 sg13g2_tiehi _29372__1110 (.L_HI(net1110));
 sg13g2_tiehi _29371__1111 (.L_HI(net1111));
 sg13g2_tiehi _29370__1112 (.L_HI(net1112));
 sg13g2_tiehi _29369__1113 (.L_HI(net1113));
 sg13g2_tiehi _29368__1114 (.L_HI(net1114));
 sg13g2_tiehi _29367__1115 (.L_HI(net1115));
 sg13g2_tiehi _29366__1116 (.L_HI(net1116));
 sg13g2_tiehi _29365__1117 (.L_HI(net1117));
 sg13g2_tiehi _29364__1118 (.L_HI(net1118));
 sg13g2_tiehi _29363__1119 (.L_HI(net1119));
 sg13g2_tiehi _29362__1120 (.L_HI(net1120));
 sg13g2_tiehi _29361__1121 (.L_HI(net1121));
 sg13g2_tiehi _29360__1122 (.L_HI(net1122));
 sg13g2_tiehi _29359__1123 (.L_HI(net1123));
 sg13g2_tiehi _29358__1124 (.L_HI(net1124));
 sg13g2_tiehi _29357__1125 (.L_HI(net1125));
 sg13g2_tiehi _29356__1126 (.L_HI(net1126));
 sg13g2_tiehi _29355__1127 (.L_HI(net1127));
 sg13g2_tiehi _29354__1128 (.L_HI(net1128));
 sg13g2_tiehi _29353__1129 (.L_HI(net1129));
 sg13g2_tiehi _29352__1130 (.L_HI(net1130));
 sg13g2_tiehi _29351__1131 (.L_HI(net1131));
 sg13g2_tiehi _29350__1132 (.L_HI(net1132));
 sg13g2_tiehi _29349__1133 (.L_HI(net1133));
 sg13g2_tiehi _29348__1134 (.L_HI(net1134));
 sg13g2_tiehi _29347__1135 (.L_HI(net1135));
 sg13g2_tiehi _29346__1136 (.L_HI(net1136));
 sg13g2_tiehi _29345__1137 (.L_HI(net1137));
 sg13g2_tiehi _29344__1138 (.L_HI(net1138));
 sg13g2_tiehi _29343__1139 (.L_HI(net1139));
 sg13g2_tiehi _29342__1140 (.L_HI(net1140));
 sg13g2_tiehi _29341__1141 (.L_HI(net1141));
 sg13g2_tiehi _29340__1142 (.L_HI(net1142));
 sg13g2_tiehi _29339__1143 (.L_HI(net1143));
 sg13g2_tiehi _29338__1144 (.L_HI(net1144));
 sg13g2_tiehi _29337__1145 (.L_HI(net1145));
 sg13g2_tiehi _29336__1146 (.L_HI(net1146));
 sg13g2_tiehi _29335__1147 (.L_HI(net1147));
 sg13g2_tiehi _29334__1148 (.L_HI(net1148));
 sg13g2_tiehi _29333__1149 (.L_HI(net1149));
 sg13g2_tiehi _29332__1150 (.L_HI(net1150));
 sg13g2_tiehi _28813__1151 (.L_HI(net1151));
 sg13g2_tiehi _28987__1152 (.L_HI(net1152));
 sg13g2_tiehi _28988__1153 (.L_HI(net1153));
 sg13g2_tiehi _28989__1154 (.L_HI(net1154));
 sg13g2_tiehi _29331__1155 (.L_HI(net1155));
 sg13g2_tiehi _29330__1156 (.L_HI(net1156));
 sg13g2_tiehi _29329__1157 (.L_HI(net1157));
 sg13g2_tiehi _29328__1158 (.L_HI(net1158));
 sg13g2_tiehi _29327__1159 (.L_HI(net1159));
 sg13g2_tiehi _29326__1160 (.L_HI(net1160));
 sg13g2_tiehi _29325__1161 (.L_HI(net1161));
 sg13g2_tiehi _29324__1162 (.L_HI(net1162));
 sg13g2_tiehi _29323__1163 (.L_HI(net1163));
 sg13g2_tiehi _29322__1164 (.L_HI(net1164));
 sg13g2_tiehi _29321__1165 (.L_HI(net1165));
 sg13g2_tiehi _29320__1166 (.L_HI(net1166));
 sg13g2_tiehi _29319__1167 (.L_HI(net1167));
 sg13g2_tiehi _29318__1168 (.L_HI(net1168));
 sg13g2_tiehi _29317__1169 (.L_HI(net1169));
 sg13g2_tiehi _29316__1170 (.L_HI(net1170));
 sg13g2_tiehi _29315__1171 (.L_HI(net1171));
 sg13g2_tiehi _29314__1172 (.L_HI(net1172));
 sg13g2_tiehi _29313__1173 (.L_HI(net1173));
 sg13g2_tiehi _29312__1174 (.L_HI(net1174));
 sg13g2_tiehi _29311__1175 (.L_HI(net1175));
 sg13g2_tiehi _29310__1176 (.L_HI(net1176));
 sg13g2_tiehi _29309__1177 (.L_HI(net1177));
 sg13g2_tiehi _29308__1178 (.L_HI(net1178));
 sg13g2_tiehi _29307__1179 (.L_HI(net1179));
 sg13g2_tiehi _29306__1180 (.L_HI(net1180));
 sg13g2_tiehi _29305__1181 (.L_HI(net1181));
 sg13g2_tiehi _29304__1182 (.L_HI(net1182));
 sg13g2_tiehi _29303__1183 (.L_HI(net1183));
 sg13g2_tiehi _29302__1184 (.L_HI(net1184));
 sg13g2_tiehi _29301__1185 (.L_HI(net1185));
 sg13g2_tiehi _29300__1186 (.L_HI(net1186));
 sg13g2_tiehi _29299__1187 (.L_HI(net1187));
 sg13g2_tiehi _28990__1188 (.L_HI(net1188));
 sg13g2_tiehi _29024__1189 (.L_HI(net1189));
 sg13g2_tiehi _29025__1190 (.L_HI(net1190));
 sg13g2_tiehi _29026__1191 (.L_HI(net1191));
 sg13g2_tiehi _29027__1192 (.L_HI(net1192));
 sg13g2_tiehi _29028__1193 (.L_HI(net1193));
 sg13g2_tiehi _29029__1194 (.L_HI(net1194));
 sg13g2_tiehi _29030__1195 (.L_HI(net1195));
 sg13g2_tiehi _29298__1196 (.L_HI(net1196));
 sg13g2_tiehi _29297__1197 (.L_HI(net1197));
 sg13g2_tiehi _29296__1198 (.L_HI(net1198));
 sg13g2_tiehi _29295__1199 (.L_HI(net1199));
 sg13g2_tiehi _29294__1200 (.L_HI(net1200));
 sg13g2_tiehi _29293__1201 (.L_HI(net1201));
 sg13g2_tiehi _29292__1202 (.L_HI(net1202));
 sg13g2_tiehi _29291__1203 (.L_HI(net1203));
 sg13g2_tiehi _29290__1204 (.L_HI(net1204));
 sg13g2_tiehi _29289__1205 (.L_HI(net1205));
 sg13g2_tiehi _29288__1206 (.L_HI(net1206));
 sg13g2_tiehi _29287__1207 (.L_HI(net1207));
 sg13g2_tiehi _29286__1208 (.L_HI(net1208));
 sg13g2_tiehi _29285__1209 (.L_HI(net1209));
 sg13g2_tiehi _29284__1210 (.L_HI(net1210));
 sg13g2_tiehi _29283__1211 (.L_HI(net1211));
 sg13g2_tiehi _29031__1212 (.L_HI(net1212));
 sg13g2_tiehi _29282__1213 (.L_HI(net1213));
 sg13g2_tiehi _29281__1214 (.L_HI(net1214));
 sg13g2_tiehi _29280__1215 (.L_HI(net1215));
 sg13g2_tiehi _29279__1216 (.L_HI(net1216));
 sg13g2_tiehi _29278__1217 (.L_HI(net1217));
 sg13g2_tiehi _29277__1218 (.L_HI(net1218));
 sg13g2_tiehi _29276__1219 (.L_HI(net1219));
 sg13g2_tiehi _29275__1220 (.L_HI(net1220));
 sg13g2_tiehi _29274__1221 (.L_HI(net1221));
 sg13g2_tiehi _29273__1222 (.L_HI(net1222));
 sg13g2_tiehi _29272__1223 (.L_HI(net1223));
 sg13g2_tiehi _29271__1224 (.L_HI(net1224));
 sg13g2_tiehi _29270__1225 (.L_HI(net1225));
 sg13g2_tiehi _29269__1226 (.L_HI(net1226));
 sg13g2_tiehi _29268__1227 (.L_HI(net1227));
 sg13g2_tiehi _29267__1228 (.L_HI(net1228));
 sg13g2_tiehi _29266__1229 (.L_HI(net1229));
 sg13g2_tiehi _29265__1230 (.L_HI(net1230));
 sg13g2_tiehi _29264__1231 (.L_HI(net1231));
 sg13g2_tiehi _29263__1232 (.L_HI(net1232));
 sg13g2_tiehi _29262__1233 (.L_HI(net1233));
 sg13g2_tiehi _29261__1234 (.L_HI(net1234));
 sg13g2_tiehi _29260__1235 (.L_HI(net1235));
 sg13g2_tiehi _29259__1236 (.L_HI(net1236));
 sg13g2_tiehi _29258__1237 (.L_HI(net1237));
 sg13g2_tiehi _29257__1238 (.L_HI(net1238));
 sg13g2_tiehi _29256__1239 (.L_HI(net1239));
 sg13g2_tiehi _29255__1240 (.L_HI(net1240));
 sg13g2_tiehi _29254__1241 (.L_HI(net1241));
 sg13g2_tiehi _29253__1242 (.L_HI(net1242));
 sg13g2_tiehi _29252__1243 (.L_HI(net1243));
 sg13g2_tiehi _29251__1244 (.L_HI(net1244));
 sg13g2_tiehi _29250__1245 (.L_HI(net1245));
 sg13g2_tiehi _29249__1246 (.L_HI(net1246));
 sg13g2_tiehi _29248__1247 (.L_HI(net1247));
 sg13g2_tiehi _29247__1248 (.L_HI(net1248));
 sg13g2_tiehi _29246__1249 (.L_HI(net1249));
 sg13g2_tiehi _29245__1250 (.L_HI(net1250));
 sg13g2_tiehi _29244__1251 (.L_HI(net1251));
 sg13g2_tiehi _29243__1252 (.L_HI(net1252));
 sg13g2_tiehi _29242__1253 (.L_HI(net1253));
 sg13g2_tiehi _29241__1254 (.L_HI(net1254));
 sg13g2_tiehi _29240__1255 (.L_HI(net1255));
 sg13g2_tiehi _29239__1256 (.L_HI(net1256));
 sg13g2_tiehi _29238__1257 (.L_HI(net1257));
 sg13g2_tiehi _29237__1258 (.L_HI(net1258));
 sg13g2_tiehi _29236__1259 (.L_HI(net1259));
 sg13g2_tiehi _29235__1260 (.L_HI(net1260));
 sg13g2_tiehi _29234__1261 (.L_HI(net1261));
 sg13g2_tiehi _29233__1262 (.L_HI(net1262));
 sg13g2_tiehi _29232__1263 (.L_HI(net1263));
 sg13g2_tiehi _29231__1264 (.L_HI(net1264));
 sg13g2_tiehi _29230__1265 (.L_HI(net1265));
 sg13g2_tiehi _29229__1266 (.L_HI(net1266));
 sg13g2_tiehi _29228__1267 (.L_HI(net1267));
 sg13g2_tiehi _29227__1268 (.L_HI(net1268));
 sg13g2_tiehi _29226__1269 (.L_HI(net1269));
 sg13g2_tiehi _29225__1270 (.L_HI(net1270));
 sg13g2_tiehi _29224__1271 (.L_HI(net1271));
 sg13g2_tiehi _29223__1272 (.L_HI(net1272));
 sg13g2_tiehi _29222__1273 (.L_HI(net1273));
 sg13g2_tiehi _29221__1274 (.L_HI(net1274));
 sg13g2_tiehi _29220__1275 (.L_HI(net1275));
 sg13g2_tiehi _29219__1276 (.L_HI(net1276));
 sg13g2_tiehi _29218__1277 (.L_HI(net1277));
 sg13g2_tiehi _29217__1278 (.L_HI(net1278));
 sg13g2_tiehi _29216__1279 (.L_HI(net1279));
 sg13g2_tiehi _29215__1280 (.L_HI(net1280));
 sg13g2_tiehi _29214__1281 (.L_HI(net1281));
 sg13g2_tiehi _29213__1282 (.L_HI(net1282));
 sg13g2_tiehi _29212__1283 (.L_HI(net1283));
 sg13g2_tiehi _29211__1284 (.L_HI(net1284));
 sg13g2_tiehi _29210__1285 (.L_HI(net1285));
 sg13g2_tiehi _29209__1286 (.L_HI(net1286));
 sg13g2_tiehi _29048__1287 (.L_HI(net1287));
 sg13g2_tiehi _29135__1288 (.L_HI(net1288));
 sg13g2_tiehi _29208__1289 (.L_HI(net1289));
 sg13g2_tiehi _29207__1290 (.L_HI(net1290));
 sg13g2_tiehi _29206__1291 (.L_HI(net1291));
 sg13g2_tiehi _29205__1292 (.L_HI(net1292));
 sg13g2_tiehi _29204__1293 (.L_HI(net1293));
 sg13g2_tiehi _29203__1294 (.L_HI(net1294));
 sg13g2_tiehi _29202__1295 (.L_HI(net1295));
 sg13g2_tiehi _29201__1296 (.L_HI(net1296));
 sg13g2_tiehi _29200__1297 (.L_HI(net1297));
 sg13g2_tiehi _29199__1298 (.L_HI(net1298));
 sg13g2_tiehi _29198__1299 (.L_HI(net1299));
 sg13g2_tiehi _29197__1300 (.L_HI(net1300));
 sg13g2_tiehi _29196__1301 (.L_HI(net1301));
 sg13g2_tiehi _29195__1302 (.L_HI(net1302));
 sg13g2_tiehi _29194__1303 (.L_HI(net1303));
 sg13g2_tiehi _29193__1304 (.L_HI(net1304));
 sg13g2_tiehi _29192__1305 (.L_HI(net1305));
 sg13g2_tiehi _29191__1306 (.L_HI(net1306));
 sg13g2_tiehi _29190__1307 (.L_HI(net1307));
 sg13g2_tiehi _29189__1308 (.L_HI(net1308));
 sg13g2_tiehi _29188__1309 (.L_HI(net1309));
 sg13g2_tiehi _29187__1310 (.L_HI(net1310));
 sg13g2_tiehi _29186__1311 (.L_HI(net1311));
 sg13g2_tiehi _29185__1312 (.L_HI(net1312));
 sg13g2_tiehi _29184__1313 (.L_HI(net1313));
 sg13g2_tiehi _29183__1314 (.L_HI(net1314));
 sg13g2_tiehi _29182__1315 (.L_HI(net1315));
 sg13g2_tiehi _29181__1316 (.L_HI(net1316));
 sg13g2_tiehi _29179__1317 (.L_HI(net1317));
 sg13g2_tiehi _29136__1318 (.L_HI(net1318));
 sg13g2_tiehi _29178__1319 (.L_HI(net1319));
 sg13g2_tiehi _29177__1320 (.L_HI(net1320));
 sg13g2_tiehi _29176__1321 (.L_HI(net1321));
 sg13g2_tiehi _29175__1322 (.L_HI(net1322));
 sg13g2_tiehi _29174__1323 (.L_HI(net1323));
 sg13g2_tiehi _29169__1324 (.L_HI(net1324));
 sg13g2_tiehi _29173__1325 (.L_HI(net1325));
 sg13g2_tiehi _29172__1326 (.L_HI(net1326));
 sg13g2_tiehi _29171__1327 (.L_HI(net1327));
 sg13g2_tiehi _29170__1328 (.L_HI(net1328));
 sg13g2_tiehi _29168__1329 (.L_HI(net1329));
 sg13g2_tiehi _29167__1330 (.L_HI(net1330));
 sg13g2_tiehi _29166__1331 (.L_HI(net1331));
 sg13g2_tiehi _29165__1332 (.L_HI(net1332));
 sg13g2_tiehi _29164__1333 (.L_HI(net1333));
 sg13g2_tiehi _29163__1334 (.L_HI(net1334));
 sg13g2_tiehi _29162__1335 (.L_HI(net1335));
 sg13g2_tiehi _29161__1336 (.L_HI(net1336));
 sg13g2_tiehi _29160__1337 (.L_HI(net1337));
 sg13g2_tiehi _29159__1338 (.L_HI(net1338));
 sg13g2_tiehi _29158__1339 (.L_HI(net1339));
 sg13g2_tiehi _29157__1340 (.L_HI(net1340));
 sg13g2_tiehi _29156__1341 (.L_HI(net1341));
 sg13g2_tiehi _29155__1342 (.L_HI(net1342));
 sg13g2_tiehi _29154__1343 (.L_HI(net1343));
 sg13g2_tiehi _29153__1344 (.L_HI(net1344));
 sg13g2_tiehi _29152__1345 (.L_HI(net1345));
 sg13g2_tiehi _29151__1346 (.L_HI(net1346));
 sg13g2_tiehi _29150__1347 (.L_HI(net1347));
 sg13g2_tiehi _29149__1348 (.L_HI(net1348));
 sg13g2_tiehi _29148__1349 (.L_HI(net1349));
 sg13g2_tiehi _29147__1350 (.L_HI(net1350));
 sg13g2_tiehi _29146__1351 (.L_HI(net1351));
 sg13g2_tiehi _29145__1352 (.L_HI(net1352));
 sg13g2_tiehi _29144__1353 (.L_HI(net1353));
 sg13g2_tiehi _29143__1354 (.L_HI(net1354));
 sg13g2_tiehi _29142__1355 (.L_HI(net1355));
 sg13g2_tiehi _29141__1356 (.L_HI(net1356));
 sg13g2_tiehi _29140__1357 (.L_HI(net1357));
 sg13g2_tiehi _29139__1358 (.L_HI(net1358));
 sg13g2_tiehi _29138__1359 (.L_HI(net1359));
 sg13g2_tiehi _29137__1360 (.L_HI(net1360));
 sg13g2_tiehi _29134__1361 (.L_HI(net1361));
 sg13g2_tiehi _29133__1362 (.L_HI(net1362));
 sg13g2_tiehi _29132__1363 (.L_HI(net1363));
 sg13g2_tiehi _29131__1364 (.L_HI(net1364));
 sg13g2_tiehi _29130__1365 (.L_HI(net1365));
 sg13g2_tiehi _29129__1366 (.L_HI(net1366));
 sg13g2_tiehi _29128__1367 (.L_HI(net1367));
 sg13g2_tiehi _29127__1368 (.L_HI(net1368));
 sg13g2_tiehi _29126__1369 (.L_HI(net1369));
 sg13g2_tiehi _29125__1370 (.L_HI(net1370));
 sg13g2_tiehi _29124__1371 (.L_HI(net1371));
 sg13g2_tiehi _29123__1372 (.L_HI(net1372));
 sg13g2_tiehi _29122__1373 (.L_HI(net1373));
 sg13g2_tiehi _29121__1374 (.L_HI(net1374));
 sg13g2_tiehi _29120__1375 (.L_HI(net1375));
 sg13g2_tiehi _29119__1376 (.L_HI(net1376));
 sg13g2_tiehi _29118__1377 (.L_HI(net1377));
 sg13g2_tiehi _29117__1378 (.L_HI(net1378));
 sg13g2_tiehi _29116__1379 (.L_HI(net1379));
 sg13g2_tiehi _29115__1380 (.L_HI(net1380));
 sg13g2_tiehi _29114__1381 (.L_HI(net1381));
 sg13g2_tiehi _29113__1382 (.L_HI(net1382));
 sg13g2_tiehi _29112__1383 (.L_HI(net1383));
 sg13g2_tiehi _29111__1384 (.L_HI(net1384));
 sg13g2_tiehi _30680__1385 (.L_HI(net1385));
 sg13g2_tiehi _29110__1386 (.L_HI(net1386));
 sg13g2_tiehi _30679__1387 (.L_HI(net1387));
 sg13g2_tiehi _29109__1388 (.L_HI(net1388));
 sg13g2_tiehi _30678__1389 (.L_HI(net1389));
 sg13g2_tiehi _29108__1390 (.L_HI(net1390));
 sg13g2_tiehi _30677__1391 (.L_HI(net1391));
 sg13g2_tiehi _29107__1392 (.L_HI(net1392));
 sg13g2_tiehi _30676__1393 (.L_HI(net1393));
 sg13g2_tiehi _29106__1394 (.L_HI(net1394));
 sg13g2_tiehi _30675__1395 (.L_HI(net1395));
 sg13g2_tiehi _29105__1396 (.L_HI(net1396));
 sg13g2_tiehi _30674__1397 (.L_HI(net1397));
 sg13g2_tiehi _29104__1398 (.L_HI(net1398));
 sg13g2_tiehi _29103__1399 (.L_HI(net1399));
 sg13g2_tiehi _29102__1400 (.L_HI(net1400));
 sg13g2_tiehi _29101__1401 (.L_HI(net1401));
 sg13g2_tiehi _29100__1402 (.L_HI(net1402));
 sg13g2_tiehi _29099__1403 (.L_HI(net1403));
 sg13g2_tiehi _29098__1404 (.L_HI(net1404));
 sg13g2_tiehi _29097__1405 (.L_HI(net1405));
 sg13g2_tiehi _29096__1406 (.L_HI(net1406));
 sg13g2_tiehi _29095__1407 (.L_HI(net1407));
 sg13g2_tiehi _29094__1408 (.L_HI(net1408));
 sg13g2_tiehi _29093__1409 (.L_HI(net1409));
 sg13g2_tiehi _29092__1410 (.L_HI(net1410));
 sg13g2_tiehi _29091__1411 (.L_HI(net1411));
 sg13g2_tiehi _29090__1412 (.L_HI(net1412));
 sg13g2_tiehi _29089__1413 (.L_HI(net1413));
 sg13g2_tiehi _29088__1414 (.L_HI(net1414));
 sg13g2_tiehi _29087__1415 (.L_HI(net1415));
 sg13g2_tiehi _29086__1416 (.L_HI(net1416));
 sg13g2_tiehi _29085__1417 (.L_HI(net1417));
 sg13g2_tiehi _29084__1418 (.L_HI(net1418));
 sg13g2_tiehi _29083__1419 (.L_HI(net1419));
 sg13g2_tiehi _29082__1420 (.L_HI(net1420));
 sg13g2_tiehi _29081__1421 (.L_HI(net1421));
 sg13g2_tiehi _29080__1422 (.L_HI(net1422));
 sg13g2_tiehi _29079__1423 (.L_HI(net1423));
 sg13g2_tiehi _29078__1424 (.L_HI(net1424));
 sg13g2_tiehi _29077__1425 (.L_HI(net1425));
 sg13g2_tiehi _29076__1426 (.L_HI(net1426));
 sg13g2_tiehi _29075__1427 (.L_HI(net1427));
 sg13g2_tiehi _29074__1428 (.L_HI(net1428));
 sg13g2_tiehi _29073__1429 (.L_HI(net1429));
 sg13g2_tiehi _29072__1430 (.L_HI(net1430));
 sg13g2_tiehi _29071__1431 (.L_HI(net1431));
 sg13g2_tiehi _29070__1432 (.L_HI(net1432));
 sg13g2_tiehi _29069__1433 (.L_HI(net1433));
 sg13g2_tiehi _29068__1434 (.L_HI(net1434));
 sg13g2_tiehi _29067__1435 (.L_HI(net1435));
 sg13g2_tiehi _29066__1436 (.L_HI(net1436));
 sg13g2_tiehi _29065__1437 (.L_HI(net1437));
 sg13g2_tiehi _29064__1438 (.L_HI(net1438));
 sg13g2_tiehi _29063__1439 (.L_HI(net1439));
 sg13g2_tiehi _29062__1440 (.L_HI(net1440));
 sg13g2_tiehi _29061__1441 (.L_HI(net1441));
 sg13g2_tiehi _29060__1442 (.L_HI(net1442));
 sg13g2_tiehi _29059__1443 (.L_HI(net1443));
 sg13g2_tiehi _29058__1444 (.L_HI(net1444));
 sg13g2_tiehi _29057__1445 (.L_HI(net1445));
 sg13g2_tiehi _29056__1446 (.L_HI(net1446));
 sg13g2_tiehi _29055__1447 (.L_HI(net1447));
 sg13g2_tiehi _29054__1448 (.L_HI(net1448));
 sg13g2_tiehi _29053__1449 (.L_HI(net1449));
 sg13g2_tiehi _29052__1450 (.L_HI(net1450));
 sg13g2_tiehi _29051__1451 (.L_HI(net1451));
 sg13g2_tiehi _29050__1452 (.L_HI(net1452));
 sg13g2_tiehi _29049__1453 (.L_HI(net1453));
 sg13g2_tiehi _29047__1454 (.L_HI(net1454));
 sg13g2_tiehi _29046__1455 (.L_HI(net1455));
 sg13g2_tiehi _29045__1456 (.L_HI(net1456));
 sg13g2_tiehi _29044__1457 (.L_HI(net1457));
 sg13g2_tiehi _29043__1458 (.L_HI(net1458));
 sg13g2_tiehi _29042__1459 (.L_HI(net1459));
 sg13g2_tiehi _29041__1460 (.L_HI(net1460));
 sg13g2_tiehi _29040__1461 (.L_HI(net1461));
 sg13g2_tiehi _29039__1462 (.L_HI(net1462));
 sg13g2_tiehi _29038__1463 (.L_HI(net1463));
 sg13g2_tiehi _29037__1464 (.L_HI(net1464));
 sg13g2_tiehi _29036__1465 (.L_HI(net1465));
 sg13g2_tiehi _29035__1466 (.L_HI(net1466));
 sg13g2_tiehi _29034__1467 (.L_HI(net1467));
 sg13g2_tiehi _29033__1468 (.L_HI(net1468));
 sg13g2_tiehi _29032__1469 (.L_HI(net1469));
 sg13g2_tiehi _29023__1470 (.L_HI(net1470));
 sg13g2_tiehi _29022__1471 (.L_HI(net1471));
 sg13g2_tiehi _29021__1472 (.L_HI(net1472));
 sg13g2_tiehi _29020__1473 (.L_HI(net1473));
 sg13g2_tiehi _29019__1474 (.L_HI(net1474));
 sg13g2_tiehi _29018__1475 (.L_HI(net1475));
 sg13g2_tiehi _29017__1476 (.L_HI(net1476));
 sg13g2_tiehi _29016__1477 (.L_HI(net1477));
 sg13g2_tiehi _29015__1478 (.L_HI(net1478));
 sg13g2_tiehi _29014__1479 (.L_HI(net1479));
 sg13g2_tiehi _29013__1480 (.L_HI(net1480));
 sg13g2_tiehi _29012__1481 (.L_HI(net1481));
 sg13g2_tiehi _29011__1482 (.L_HI(net1482));
 sg13g2_tiehi _29010__1483 (.L_HI(net1483));
 sg13g2_tiehi _29009__1484 (.L_HI(net1484));
 sg13g2_tiehi _29008__1485 (.L_HI(net1485));
 sg13g2_tiehi _29007__1486 (.L_HI(net1486));
 sg13g2_tiehi _29006__1487 (.L_HI(net1487));
 sg13g2_tiehi _29005__1488 (.L_HI(net1488));
 sg13g2_tiehi _29004__1489 (.L_HI(net1489));
 sg13g2_tiehi _29003__1490 (.L_HI(net1490));
 sg13g2_tiehi _29002__1491 (.L_HI(net1491));
 sg13g2_tiehi _29001__1492 (.L_HI(net1492));
 sg13g2_tiehi _29000__1493 (.L_HI(net1493));
 sg13g2_tiehi _28999__1494 (.L_HI(net1494));
 sg13g2_tiehi _28998__1495 (.L_HI(net1495));
 sg13g2_tiehi _28997__1496 (.L_HI(net1496));
 sg13g2_tiehi _28996__1497 (.L_HI(net1497));
 sg13g2_tiehi _28995__1498 (.L_HI(net1498));
 sg13g2_tiehi _28994__1499 (.L_HI(net1499));
 sg13g2_tiehi _28993__1500 (.L_HI(net1500));
 sg13g2_tiehi _28992__1501 (.L_HI(net1501));
 sg13g2_tiehi _28991__1502 (.L_HI(net1502));
 sg13g2_tiehi _28986__1503 (.L_HI(net1503));
 sg13g2_tiehi _28985__1504 (.L_HI(net1504));
 sg13g2_tiehi _28984__1505 (.L_HI(net1505));
 sg13g2_tiehi _28983__1506 (.L_HI(net1506));
 sg13g2_tiehi _28982__1507 (.L_HI(net1507));
 sg13g2_tiehi _28981__1508 (.L_HI(net1508));
 sg13g2_tiehi _28980__1509 (.L_HI(net1509));
 sg13g2_tiehi _28979__1510 (.L_HI(net1510));
 sg13g2_tiehi _28978__1511 (.L_HI(net1511));
 sg13g2_tiehi _28977__1512 (.L_HI(net1512));
 sg13g2_tiehi _28976__1513 (.L_HI(net1513));
 sg13g2_tiehi _28975__1514 (.L_HI(net1514));
 sg13g2_tiehi _28974__1515 (.L_HI(net1515));
 sg13g2_tiehi _28973__1516 (.L_HI(net1516));
 sg13g2_tiehi _28972__1517 (.L_HI(net1517));
 sg13g2_tiehi _28971__1518 (.L_HI(net1518));
 sg13g2_tiehi _28970__1519 (.L_HI(net1519));
 sg13g2_tiehi _28969__1520 (.L_HI(net1520));
 sg13g2_tiehi _28968__1521 (.L_HI(net1521));
 sg13g2_tiehi _28967__1522 (.L_HI(net1522));
 sg13g2_tiehi _28966__1523 (.L_HI(net1523));
 sg13g2_tiehi _28965__1524 (.L_HI(net1524));
 sg13g2_tiehi _28964__1525 (.L_HI(net1525));
 sg13g2_tiehi _28963__1526 (.L_HI(net1526));
 sg13g2_tiehi _28962__1527 (.L_HI(net1527));
 sg13g2_tiehi _28961__1528 (.L_HI(net1528));
 sg13g2_tiehi _28960__1529 (.L_HI(net1529));
 sg13g2_tiehi _28959__1530 (.L_HI(net1530));
 sg13g2_tiehi _28958__1531 (.L_HI(net1531));
 sg13g2_tiehi _28957__1532 (.L_HI(net1532));
 sg13g2_tiehi _28956__1533 (.L_HI(net1533));
 sg13g2_tiehi _28955__1534 (.L_HI(net1534));
 sg13g2_tiehi _28954__1535 (.L_HI(net1535));
 sg13g2_tiehi _28953__1536 (.L_HI(net1536));
 sg13g2_tiehi _28952__1537 (.L_HI(net1537));
 sg13g2_tiehi _28951__1538 (.L_HI(net1538));
 sg13g2_tiehi _28950__1539 (.L_HI(net1539));
 sg13g2_tiehi _28949__1540 (.L_HI(net1540));
 sg13g2_tiehi _28948__1541 (.L_HI(net1541));
 sg13g2_tiehi _28947__1542 (.L_HI(net1542));
 sg13g2_tiehi _28946__1543 (.L_HI(net1543));
 sg13g2_tiehi _28945__1544 (.L_HI(net1544));
 sg13g2_tiehi _28944__1545 (.L_HI(net1545));
 sg13g2_tiehi _28943__1546 (.L_HI(net1546));
 sg13g2_tiehi _28942__1547 (.L_HI(net1547));
 sg13g2_tiehi _28941__1548 (.L_HI(net1548));
 sg13g2_tiehi _28940__1549 (.L_HI(net1549));
 sg13g2_tiehi _28939__1550 (.L_HI(net1550));
 sg13g2_tiehi _28938__1551 (.L_HI(net1551));
 sg13g2_tiehi _28937__1552 (.L_HI(net1552));
 sg13g2_tiehi _28936__1553 (.L_HI(net1553));
 sg13g2_tiehi _28935__1554 (.L_HI(net1554));
 sg13g2_tiehi _28934__1555 (.L_HI(net1555));
 sg13g2_tiehi _28933__1556 (.L_HI(net1556));
 sg13g2_tiehi _28932__1557 (.L_HI(net1557));
 sg13g2_tiehi _28931__1558 (.L_HI(net1558));
 sg13g2_tiehi _28930__1559 (.L_HI(net1559));
 sg13g2_tiehi _28929__1560 (.L_HI(net1560));
 sg13g2_tiehi _28928__1561 (.L_HI(net1561));
 sg13g2_tiehi _28927__1562 (.L_HI(net1562));
 sg13g2_tiehi _28926__1563 (.L_HI(net1563));
 sg13g2_tiehi _28925__1564 (.L_HI(net1564));
 sg13g2_tiehi _28924__1565 (.L_HI(net1565));
 sg13g2_tiehi _28923__1566 (.L_HI(net1566));
 sg13g2_tiehi _28922__1567 (.L_HI(net1567));
 sg13g2_tiehi _28921__1568 (.L_HI(net1568));
 sg13g2_tiehi _28920__1569 (.L_HI(net1569));
 sg13g2_tiehi _28919__1570 (.L_HI(net1570));
 sg13g2_tiehi _28918__1571 (.L_HI(net1571));
 sg13g2_tiehi _28917__1572 (.L_HI(net1572));
 sg13g2_tiehi _28916__1573 (.L_HI(net1573));
 sg13g2_tiehi _28915__1574 (.L_HI(net1574));
 sg13g2_tiehi _28914__1575 (.L_HI(net1575));
 sg13g2_tiehi _28913__1576 (.L_HI(net1576));
 sg13g2_tiehi _28912__1577 (.L_HI(net1577));
 sg13g2_tiehi _28911__1578 (.L_HI(net1578));
 sg13g2_tiehi _28910__1579 (.L_HI(net1579));
 sg13g2_tiehi _28909__1580 (.L_HI(net1580));
 sg13g2_tiehi _28908__1581 (.L_HI(net1581));
 sg13g2_tiehi _28907__1582 (.L_HI(net1582));
 sg13g2_tiehi _29180__1583 (.L_HI(net1583));
 sg13g2_tiehi _29472__1584 (.L_HI(net1584));
 sg13g2_tiehi _29473__1585 (.L_HI(net1585));
 sg13g2_tiehi _29474__1586 (.L_HI(net1586));
 sg13g2_tiehi _29475__1587 (.L_HI(net1587));
 sg13g2_tiehi _29476__1588 (.L_HI(net1588));
 sg13g2_tiehi _29477__1589 (.L_HI(net1589));
 sg13g2_tiehi _29478__1590 (.L_HI(net1590));
 sg13g2_tiehi _28906__1591 (.L_HI(net1591));
 sg13g2_tiehi _28905__1592 (.L_HI(net1592));
 sg13g2_tiehi _28904__1593 (.L_HI(net1593));
 sg13g2_tiehi _28903__1594 (.L_HI(net1594));
 sg13g2_tiehi _28902__1595 (.L_HI(net1595));
 sg13g2_tiehi _28901__1596 (.L_HI(net1596));
 sg13g2_tiehi _28900__1597 (.L_HI(net1597));
 sg13g2_tiehi _28899__1598 (.L_HI(net1598));
 sg13g2_tiehi _28898__1599 (.L_HI(net1599));
 sg13g2_tiehi _28897__1600 (.L_HI(net1600));
 sg13g2_tiehi _28896__1601 (.L_HI(net1601));
 sg13g2_tiehi _28895__1602 (.L_HI(net1602));
 sg13g2_tiehi _28894__1603 (.L_HI(net1603));
 sg13g2_tiehi _28893__1604 (.L_HI(net1604));
 sg13g2_tiehi _28892__1605 (.L_HI(net1605));
 sg13g2_tiehi _28891__1606 (.L_HI(net1606));
 sg13g2_tiehi _28890__1607 (.L_HI(net1607));
 sg13g2_tiehi _28889__1608 (.L_HI(net1608));
 sg13g2_tiehi _28888__1609 (.L_HI(net1609));
 sg13g2_tiehi _28887__1610 (.L_HI(net1610));
 sg13g2_tiehi _28886__1611 (.L_HI(net1611));
 sg13g2_tiehi _28885__1612 (.L_HI(net1612));
 sg13g2_tiehi _28884__1613 (.L_HI(net1613));
 sg13g2_tiehi _28883__1614 (.L_HI(net1614));
 sg13g2_tiehi _28882__1615 (.L_HI(net1615));
 sg13g2_tiehi _28881__1616 (.L_HI(net1616));
 sg13g2_tiehi _28880__1617 (.L_HI(net1617));
 sg13g2_tiehi _28879__1618 (.L_HI(net1618));
 sg13g2_tiehi _28878__1619 (.L_HI(net1619));
 sg13g2_tiehi _28877__1620 (.L_HI(net1620));
 sg13g2_tiehi _28876__1621 (.L_HI(net1621));
 sg13g2_tiehi _28875__1622 (.L_HI(net1622));
 sg13g2_tiehi _28874__1623 (.L_HI(net1623));
 sg13g2_tiehi _28873__1624 (.L_HI(net1624));
 sg13g2_tiehi _28872__1625 (.L_HI(net1625));
 sg13g2_tiehi _28871__1626 (.L_HI(net1626));
 sg13g2_tiehi _28870__1627 (.L_HI(net1627));
 sg13g2_tiehi _28869__1628 (.L_HI(net1628));
 sg13g2_tiehi _28868__1629 (.L_HI(net1629));
 sg13g2_tiehi _28867__1630 (.L_HI(net1630));
 sg13g2_tiehi _28866__1631 (.L_HI(net1631));
 sg13g2_tiehi _28865__1632 (.L_HI(net1632));
 sg13g2_tiehi _28864__1633 (.L_HI(net1633));
 sg13g2_tiehi _28863__1634 (.L_HI(net1634));
 sg13g2_tiehi _28862__1635 (.L_HI(net1635));
 sg13g2_tiehi _28861__1636 (.L_HI(net1636));
 sg13g2_tiehi _28860__1637 (.L_HI(net1637));
 sg13g2_tiehi _28859__1638 (.L_HI(net1638));
 sg13g2_tiehi _28858__1639 (.L_HI(net1639));
 sg13g2_tiehi _28857__1640 (.L_HI(net1640));
 sg13g2_tiehi _28856__1641 (.L_HI(net1641));
 sg13g2_tiehi _28855__1642 (.L_HI(net1642));
 sg13g2_tiehi _28854__1643 (.L_HI(net1643));
 sg13g2_tiehi _28853__1644 (.L_HI(net1644));
 sg13g2_tiehi _28852__1645 (.L_HI(net1645));
 sg13g2_tiehi _28851__1646 (.L_HI(net1646));
 sg13g2_tiehi _28850__1647 (.L_HI(net1647));
 sg13g2_tiehi _28849__1648 (.L_HI(net1648));
 sg13g2_tiehi _28848__1649 (.L_HI(net1649));
 sg13g2_tiehi _28847__1650 (.L_HI(net1650));
 sg13g2_tiehi _28846__1651 (.L_HI(net1651));
 sg13g2_tiehi _28845__1652 (.L_HI(net1652));
 sg13g2_tiehi _28844__1653 (.L_HI(net1653));
 sg13g2_tiehi _28843__1654 (.L_HI(net1654));
 sg13g2_tiehi _28842__1655 (.L_HI(net1655));
 sg13g2_tiehi _28841__1656 (.L_HI(net1656));
 sg13g2_tiehi _28840__1657 (.L_HI(net1657));
 sg13g2_tiehi _28839__1658 (.L_HI(net1658));
 sg13g2_tiehi _28838__1659 (.L_HI(net1659));
 sg13g2_tiehi _28837__1660 (.L_HI(net1660));
 sg13g2_tiehi _28836__1661 (.L_HI(net1661));
 sg13g2_tiehi _28835__1662 (.L_HI(net1662));
 sg13g2_tiehi _28834__1663 (.L_HI(net1663));
 sg13g2_tiehi _30673__1664 (.L_HI(net1664));
 sg13g2_tiehi _28833__1665 (.L_HI(net1665));
 sg13g2_tiehi _30672__1666 (.L_HI(net1666));
 sg13g2_tiehi _28832__1667 (.L_HI(net1667));
 sg13g2_tiehi _30671__1668 (.L_HI(net1668));
 sg13g2_tiehi _28831__1669 (.L_HI(net1669));
 sg13g2_tiehi _30670__1670 (.L_HI(net1670));
 sg13g2_tiehi _28830__1671 (.L_HI(net1671));
 sg13g2_tiehi _30669__1672 (.L_HI(net1672));
 sg13g2_tiehi _28829__1673 (.L_HI(net1673));
 sg13g2_tiehi _30668__1674 (.L_HI(net1674));
 sg13g2_tiehi _28828__1675 (.L_HI(net1675));
 sg13g2_tiehi _30667__1676 (.L_HI(net1676));
 sg13g2_tiehi _28827__1677 (.L_HI(net1677));
 sg13g2_tiehi _28826__1678 (.L_HI(net1678));
 sg13g2_tiehi _28825__1679 (.L_HI(net1679));
 sg13g2_tiehi _28824__1680 (.L_HI(net1680));
 sg13g2_tiehi _28823__1681 (.L_HI(net1681));
 sg13g2_tiehi _28822__1682 (.L_HI(net1682));
 sg13g2_tiehi _28821__1683 (.L_HI(net1683));
 sg13g2_tiehi _28820__1684 (.L_HI(net1684));
 sg13g2_tiehi _28819__1685 (.L_HI(net1685));
 sg13g2_tiehi _28818__1686 (.L_HI(net1686));
 sg13g2_tiehi _28817__1687 (.L_HI(net1687));
 sg13g2_tiehi _28816__1688 (.L_HI(net1688));
 sg13g2_tiehi _28815__1689 (.L_HI(net1689));
 sg13g2_tiehi _28814__1690 (.L_HI(net1690));
 sg13g2_tiehi _28798__1691 (.L_HI(net1691));
 sg13g2_tiehi _28797__1692 (.L_HI(net1692));
 sg13g2_tiehi _28796__1693 (.L_HI(net1693));
 sg13g2_tiehi _28795__1694 (.L_HI(net1694));
 sg13g2_tiehi _28794__1695 (.L_HI(net1695));
 sg13g2_tiehi _28793__1696 (.L_HI(net1696));
 sg13g2_tiehi _28792__1697 (.L_HI(net1697));
 sg13g2_tiehi _28791__1698 (.L_HI(net1698));
 sg13g2_tiehi _28790__1699 (.L_HI(net1699));
 sg13g2_tiehi _28789__1700 (.L_HI(net1700));
 sg13g2_tiehi _28788__1701 (.L_HI(net1701));
 sg13g2_tiehi _28787__1702 (.L_HI(net1702));
 sg13g2_tiehi _28786__1703 (.L_HI(net1703));
 sg13g2_tiehi _28785__1704 (.L_HI(net1704));
 sg13g2_tiehi _28784__1705 (.L_HI(net1705));
 sg13g2_tiehi _28783__1706 (.L_HI(net1706));
 sg13g2_tiehi _28782__1707 (.L_HI(net1707));
 sg13g2_tiehi _28781__1708 (.L_HI(net1708));
 sg13g2_tiehi _28780__1709 (.L_HI(net1709));
 sg13g2_tiehi _28779__1710 (.L_HI(net1710));
 sg13g2_tiehi _28778__1711 (.L_HI(net1711));
 sg13g2_tiehi _28777__1712 (.L_HI(net1712));
 sg13g2_tiehi _28776__1713 (.L_HI(net1713));
 sg13g2_tiehi _28775__1714 (.L_HI(net1714));
 sg13g2_tiehi _28774__1715 (.L_HI(net1715));
 sg13g2_tiehi _28773__1716 (.L_HI(net1716));
 sg13g2_tiehi _28772__1717 (.L_HI(net1717));
 sg13g2_tiehi _28771__1718 (.L_HI(net1718));
 sg13g2_tiehi _28770__1719 (.L_HI(net1719));
 sg13g2_tiehi _28769__1720 (.L_HI(net1720));
 sg13g2_tiehi _28768__1721 (.L_HI(net1721));
 sg13g2_tiehi _28767__1722 (.L_HI(net1722));
 sg13g2_tiehi _28766__1723 (.L_HI(net1723));
 sg13g2_tiehi _28765__1724 (.L_HI(net1724));
 sg13g2_tiehi _28764__1725 (.L_HI(net1725));
 sg13g2_tiehi _28763__1726 (.L_HI(net1726));
 sg13g2_tiehi _28762__1727 (.L_HI(net1727));
 sg13g2_tiehi _28761__1728 (.L_HI(net1728));
 sg13g2_tiehi _28760__1729 (.L_HI(net1729));
 sg13g2_tiehi _28759__1730 (.L_HI(net1730));
 sg13g2_tiehi _28758__1731 (.L_HI(net1731));
 sg13g2_tiehi _28757__1732 (.L_HI(net1732));
 sg13g2_tiehi _28756__1733 (.L_HI(net1733));
 sg13g2_tiehi _28755__1734 (.L_HI(net1734));
 sg13g2_tiehi _28754__1735 (.L_HI(net1735));
 sg13g2_tiehi _28753__1736 (.L_HI(net1736));
 sg13g2_tiehi _28752__1737 (.L_HI(net1737));
 sg13g2_tiehi _28751__1738 (.L_HI(net1738));
 sg13g2_tiehi _28750__1739 (.L_HI(net1739));
 sg13g2_tiehi _28749__1740 (.L_HI(net1740));
 sg13g2_tiehi _30666__1741 (.L_HI(net1741));
 sg13g2_tiehi _28748__1742 (.L_HI(net1742));
 sg13g2_tiehi _30665__1743 (.L_HI(net1743));
 sg13g2_tiehi _28747__1744 (.L_HI(net1744));
 sg13g2_tiehi _30664__1745 (.L_HI(net1745));
 sg13g2_tiehi _28746__1746 (.L_HI(net1746));
 sg13g2_tiehi _30663__1747 (.L_HI(net1747));
 sg13g2_tiehi _28745__1748 (.L_HI(net1748));
 sg13g2_tiehi _30662__1749 (.L_HI(net1749));
 sg13g2_tiehi _28744__1750 (.L_HI(net1750));
 sg13g2_tiehi _30661__1751 (.L_HI(net1751));
 sg13g2_tiehi _28743__1752 (.L_HI(net1752));
 sg13g2_tiehi _30660__1753 (.L_HI(net1753));
 sg13g2_tiehi _28742__1754 (.L_HI(net1754));
 sg13g2_tiehi _28741__1755 (.L_HI(net1755));
 sg13g2_tiehi _28740__1756 (.L_HI(net1756));
 sg13g2_tiehi _28739__1757 (.L_HI(net1757));
 sg13g2_tiehi _28738__1758 (.L_HI(net1758));
 sg13g2_tiehi _28737__1759 (.L_HI(net1759));
 sg13g2_tiehi _28736__1760 (.L_HI(net1760));
 sg13g2_tiehi _28735__1761 (.L_HI(net1761));
 sg13g2_tiehi _28734__1762 (.L_HI(net1762));
 sg13g2_tiehi _28733__1763 (.L_HI(net1763));
 sg13g2_tiehi _28732__1764 (.L_HI(net1764));
 sg13g2_tiehi _28731__1765 (.L_HI(net1765));
 sg13g2_tiehi _28730__1766 (.L_HI(net1766));
 sg13g2_tiehi _28729__1767 (.L_HI(net1767));
 sg13g2_tiehi _28728__1768 (.L_HI(net1768));
 sg13g2_tiehi _28727__1769 (.L_HI(net1769));
 sg13g2_tiehi _28726__1770 (.L_HI(net1770));
 sg13g2_tiehi _28725__1771 (.L_HI(net1771));
 sg13g2_tiehi _28724__1772 (.L_HI(net1772));
 sg13g2_tiehi _28723__1773 (.L_HI(net1773));
 sg13g2_tiehi _28722__1774 (.L_HI(net1774));
 sg13g2_tiehi _28721__1775 (.L_HI(net1775));
 sg13g2_tiehi _28720__1776 (.L_HI(net1776));
 sg13g2_tiehi _28719__1777 (.L_HI(net1777));
 sg13g2_tiehi _28718__1778 (.L_HI(net1778));
 sg13g2_tiehi _28717__1779 (.L_HI(net1779));
 sg13g2_tiehi _28716__1780 (.L_HI(net1780));
 sg13g2_tiehi _28715__1781 (.L_HI(net1781));
 sg13g2_tiehi _28714__1782 (.L_HI(net1782));
 sg13g2_tiehi _28713__1783 (.L_HI(net1783));
 sg13g2_tiehi _28712__1784 (.L_HI(net1784));
 sg13g2_tiehi _28711__1785 (.L_HI(net1785));
 sg13g2_tiehi _28710__1786 (.L_HI(net1786));
 sg13g2_tiehi _28709__1787 (.L_HI(net1787));
 sg13g2_tiehi _28708__1788 (.L_HI(net1788));
 sg13g2_tiehi _28707__1789 (.L_HI(net1789));
 sg13g2_tiehi _28706__1790 (.L_HI(net1790));
 sg13g2_tiehi _28705__1791 (.L_HI(net1791));
 sg13g2_tiehi _28704__1792 (.L_HI(net1792));
 sg13g2_tiehi _28703__1793 (.L_HI(net1793));
 sg13g2_tiehi _28702__1794 (.L_HI(net1794));
 sg13g2_tiehi _28701__1795 (.L_HI(net1795));
 sg13g2_tiehi _28700__1796 (.L_HI(net1796));
 sg13g2_tiehi _28699__1797 (.L_HI(net1797));
 sg13g2_tiehi _28698__1798 (.L_HI(net1798));
 sg13g2_tiehi _28697__1799 (.L_HI(net1799));
 sg13g2_tiehi _28696__1800 (.L_HI(net1800));
 sg13g2_tiehi _28695__1801 (.L_HI(net1801));
 sg13g2_tiehi _28694__1802 (.L_HI(net1802));
 sg13g2_tiehi _28693__1803 (.L_HI(net1803));
 sg13g2_tiehi _28692__1804 (.L_HI(net1804));
 sg13g2_tiehi _28691__1805 (.L_HI(net1805));
 sg13g2_tiehi _28690__1806 (.L_HI(net1806));
 sg13g2_tiehi _28689__1807 (.L_HI(net1807));
 sg13g2_tiehi _28688__1808 (.L_HI(net1808));
 sg13g2_tiehi _28687__1809 (.L_HI(net1809));
 sg13g2_tiehi _28686__1810 (.L_HI(net1810));
 sg13g2_tiehi _28685__1811 (.L_HI(net1811));
 sg13g2_tiehi _28684__1812 (.L_HI(net1812));
 sg13g2_tiehi _28683__1813 (.L_HI(net1813));
 sg13g2_tiehi _28682__1814 (.L_HI(net1814));
 sg13g2_tiehi _28681__1815 (.L_HI(net1815));
 sg13g2_tiehi _28680__1816 (.L_HI(net1816));
 sg13g2_tiehi _28679__1817 (.L_HI(net1817));
 sg13g2_tiehi _28678__1818 (.L_HI(net1818));
 sg13g2_tiehi _28677__1819 (.L_HI(net1819));
 sg13g2_tiehi _28676__1820 (.L_HI(net1820));
 sg13g2_tiehi _28675__1821 (.L_HI(net1821));
 sg13g2_tiehi _28674__1822 (.L_HI(net1822));
 sg13g2_tiehi _28673__1823 (.L_HI(net1823));
 sg13g2_tiehi _28672__1824 (.L_HI(net1824));
 sg13g2_tiehi _28671__1825 (.L_HI(net1825));
 sg13g2_tiehi _28670__1826 (.L_HI(net1826));
 sg13g2_tiehi _28669__1827 (.L_HI(net1827));
 sg13g2_tiehi _28668__1828 (.L_HI(net1828));
 sg13g2_tiehi _28667__1829 (.L_HI(net1829));
 sg13g2_tiehi _28666__1830 (.L_HI(net1830));
 sg13g2_tiehi _28665__1831 (.L_HI(net1831));
 sg13g2_tiehi _28664__1832 (.L_HI(net1832));
 sg13g2_tiehi _30659__1833 (.L_HI(net1833));
 sg13g2_tiehi _28663__1834 (.L_HI(net1834));
 sg13g2_tiehi _28662__1835 (.L_HI(net1835));
 sg13g2_tiehi _28661__1836 (.L_HI(net1836));
 sg13g2_tiehi _28660__1837 (.L_HI(net1837));
 sg13g2_tiehi _30658__1838 (.L_HI(net1838));
 sg13g2_tiehi _28659__1839 (.L_HI(net1839));
 sg13g2_tiehi _30657__1840 (.L_HI(net1840));
 sg13g2_tiehi _28658__1841 (.L_HI(net1841));
 sg13g2_tiehi _30656__1842 (.L_HI(net1842));
 sg13g2_tiehi _28657__1843 (.L_HI(net1843));
 sg13g2_tiehi _30655__1844 (.L_HI(net1844));
 sg13g2_tiehi _28639__1845 (.L_HI(net1845));
 sg13g2_tiehi _30654__1846 (.L_HI(net1846));
 sg13g2_tiehi _28638__1847 (.L_HI(net1847));
 sg13g2_tiehi _30653__1848 (.L_HI(net1848));
 sg13g2_tiehi _28637__1849 (.L_HI(net1849));
 sg13g2_tiehi _28636__1850 (.L_HI(net1850));
 sg13g2_tiehi _28635__1851 (.L_HI(net1851));
 sg13g2_tiehi _28634__1852 (.L_HI(net1852));
 sg13g2_tiehi _28633__1853 (.L_HI(net1853));
 sg13g2_tiehi _28632__1854 (.L_HI(net1854));
 sg13g2_tiehi _28631__1855 (.L_HI(net1855));
 sg13g2_tiehi _28630__1856 (.L_HI(net1856));
 sg13g2_tiehi _28629__1857 (.L_HI(net1857));
 sg13g2_tiehi _28628__1858 (.L_HI(net1858));
 sg13g2_tiehi _28627__1859 (.L_HI(net1859));
 sg13g2_tiehi _28626__1860 (.L_HI(net1860));
 sg13g2_tiehi _28625__1861 (.L_HI(net1861));
 sg13g2_tiehi _28624__1862 (.L_HI(net1862));
 sg13g2_tiehi _28623__1863 (.L_HI(net1863));
 sg13g2_tiehi _28622__1864 (.L_HI(net1864));
 sg13g2_tiehi _28621__1865 (.L_HI(net1865));
 sg13g2_tiehi _28620__1866 (.L_HI(net1866));
 sg13g2_tiehi _28619__1867 (.L_HI(net1867));
 sg13g2_tiehi _28618__1868 (.L_HI(net1868));
 sg13g2_tiehi _28617__1869 (.L_HI(net1869));
 sg13g2_tiehi _28616__1870 (.L_HI(net1870));
 sg13g2_tiehi _28615__1871 (.L_HI(net1871));
 sg13g2_tiehi _28614__1872 (.L_HI(net1872));
 sg13g2_tiehi _28613__1873 (.L_HI(net1873));
 sg13g2_tiehi _28612__1874 (.L_HI(net1874));
 sg13g2_tiehi _28611__1875 (.L_HI(net1875));
 sg13g2_tiehi _28610__1876 (.L_HI(net1876));
 sg13g2_tiehi _28609__1877 (.L_HI(net1877));
 sg13g2_tiehi _28608__1878 (.L_HI(net1878));
 sg13g2_tiehi _28607__1879 (.L_HI(net1879));
 sg13g2_tiehi _28606__1880 (.L_HI(net1880));
 sg13g2_tiehi _28605__1881 (.L_HI(net1881));
 sg13g2_tiehi _28604__1882 (.L_HI(net1882));
 sg13g2_tiehi _28603__1883 (.L_HI(net1883));
 sg13g2_tiehi _28602__1884 (.L_HI(net1884));
 sg13g2_tiehi _28601__1885 (.L_HI(net1885));
 sg13g2_tiehi _28600__1886 (.L_HI(net1886));
 sg13g2_tiehi _28599__1887 (.L_HI(net1887));
 sg13g2_tiehi _28598__1888 (.L_HI(net1888));
 sg13g2_tiehi _28597__1889 (.L_HI(net1889));
 sg13g2_tiehi _28596__1890 (.L_HI(net1890));
 sg13g2_tiehi _28595__1891 (.L_HI(net1891));
 sg13g2_tiehi _28594__1892 (.L_HI(net1892));
 sg13g2_tiehi _28593__1893 (.L_HI(net1893));
 sg13g2_tiehi _28592__1894 (.L_HI(net1894));
 sg13g2_tiehi _28591__1895 (.L_HI(net1895));
 sg13g2_tiehi _28590__1896 (.L_HI(net1896));
 sg13g2_tiehi _28589__1897 (.L_HI(net1897));
 sg13g2_tiehi _28588__1898 (.L_HI(net1898));
 sg13g2_tiehi _28587__1899 (.L_HI(net1899));
 sg13g2_tiehi _28586__1900 (.L_HI(net1900));
 sg13g2_tiehi _28585__1901 (.L_HI(net1901));
 sg13g2_tiehi _28584__1902 (.L_HI(net1902));
 sg13g2_tiehi _28583__1903 (.L_HI(net1903));
 sg13g2_tiehi _28582__1904 (.L_HI(net1904));
 sg13g2_tiehi _28581__1905 (.L_HI(net1905));
 sg13g2_tiehi _28580__1906 (.L_HI(net1906));
 sg13g2_tiehi _28579__1907 (.L_HI(net1907));
 sg13g2_tiehi _28578__1908 (.L_HI(net1908));
 sg13g2_tiehi _28577__1909 (.L_HI(net1909));
 sg13g2_tiehi _28576__1910 (.L_HI(net1910));
 sg13g2_tiehi _28575__1911 (.L_HI(net1911));
 sg13g2_tiehi _28574__1912 (.L_HI(net1912));
 sg13g2_tiehi _28573__1913 (.L_HI(net1913));
 sg13g2_tiehi _28572__1914 (.L_HI(net1914));
 sg13g2_tiehi _28571__1915 (.L_HI(net1915));
 sg13g2_tiehi _28570__1916 (.L_HI(net1916));
 sg13g2_tiehi _28569__1917 (.L_HI(net1917));
 sg13g2_tiehi _28568__1918 (.L_HI(net1918));
 sg13g2_tiehi _28567__1919 (.L_HI(net1919));
 sg13g2_tiehi _28566__1920 (.L_HI(net1920));
 sg13g2_tiehi _28565__1921 (.L_HI(net1921));
 sg13g2_tiehi _28564__1922 (.L_HI(net1922));
 sg13g2_tiehi _28563__1923 (.L_HI(net1923));
 sg13g2_tiehi _28562__1924 (.L_HI(net1924));
 sg13g2_tiehi _28561__1925 (.L_HI(net1925));
 sg13g2_tiehi _28560__1926 (.L_HI(net1926));
 sg13g2_tiehi _28559__1927 (.L_HI(net1927));
 sg13g2_tiehi _28558__1928 (.L_HI(net1928));
 sg13g2_tiehi _28557__1929 (.L_HI(net1929));
 sg13g2_tiehi _28556__1930 (.L_HI(net1930));
 sg13g2_tiehi _28555__1931 (.L_HI(net1931));
 sg13g2_tiehi _28554__1932 (.L_HI(net1932));
 sg13g2_tiehi _28553__1933 (.L_HI(net1933));
 sg13g2_tiehi _28552__1934 (.L_HI(net1934));
 sg13g2_tiehi _28551__1935 (.L_HI(net1935));
 sg13g2_tiehi _28550__1936 (.L_HI(net1936));
 sg13g2_tiehi _28549__1937 (.L_HI(net1937));
 sg13g2_tiehi _28548__1938 (.L_HI(net1938));
 sg13g2_tiehi _28547__1939 (.L_HI(net1939));
 sg13g2_tiehi _28546__1940 (.L_HI(net1940));
 sg13g2_tiehi _28545__1941 (.L_HI(net1941));
 sg13g2_tiehi _28544__1942 (.L_HI(net1942));
 sg13g2_tiehi _28543__1943 (.L_HI(net1943));
 sg13g2_tiehi _28542__1944 (.L_HI(net1944));
 sg13g2_tiehi _30652__1945 (.L_HI(net1945));
 sg13g2_tiehi _28541__1946 (.L_HI(net1946));
 sg13g2_tiehi _30651__1947 (.L_HI(net1947));
 sg13g2_tiehi _28540__1948 (.L_HI(net1948));
 sg13g2_tiehi _30650__1949 (.L_HI(net1949));
 sg13g2_tiehi _28539__1950 (.L_HI(net1950));
 sg13g2_tiehi _30649__1951 (.L_HI(net1951));
 sg13g2_tiehi _28538__1952 (.L_HI(net1952));
 sg13g2_tiehi _28537__1953 (.L_HI(net1953));
 sg13g2_tiehi _28536__1954 (.L_HI(net1954));
 sg13g2_tiehi _28535__1955 (.L_HI(net1955));
 sg13g2_tiehi _28534__1956 (.L_HI(net1956));
 sg13g2_tiehi _28533__1957 (.L_HI(net1957));
 sg13g2_tiehi _28532__1958 (.L_HI(net1958));
 sg13g2_tiehi _28531__1959 (.L_HI(net1959));
 sg13g2_tiehi _28530__1960 (.L_HI(net1960));
 sg13g2_tiehi _28529__1961 (.L_HI(net1961));
 sg13g2_tiehi _28528__1962 (.L_HI(net1962));
 sg13g2_tiehi _28527__1963 (.L_HI(net1963));
 sg13g2_tiehi _28526__1964 (.L_HI(net1964));
 sg13g2_tiehi _28525__1965 (.L_HI(net1965));
 sg13g2_tiehi _28524__1966 (.L_HI(net1966));
 sg13g2_tiehi _28523__1967 (.L_HI(net1967));
 sg13g2_tiehi _28522__1968 (.L_HI(net1968));
 sg13g2_tiehi _28521__1969 (.L_HI(net1969));
 sg13g2_tiehi _28520__1970 (.L_HI(net1970));
 sg13g2_tiehi _28519__1971 (.L_HI(net1971));
 sg13g2_tiehi _28518__1972 (.L_HI(net1972));
 sg13g2_tiehi _28517__1973 (.L_HI(net1973));
 sg13g2_tiehi _28516__1974 (.L_HI(net1974));
 sg13g2_tiehi _28515__1975 (.L_HI(net1975));
 sg13g2_tiehi _28514__1976 (.L_HI(net1976));
 sg13g2_tiehi _28513__1977 (.L_HI(net1977));
 sg13g2_tiehi _30648__1978 (.L_HI(net1978));
 sg13g2_tiehi _28512__1979 (.L_HI(net1979));
 sg13g2_tiehi _30647__1980 (.L_HI(net1980));
 sg13g2_tiehi _28511__1981 (.L_HI(net1981));
 sg13g2_tiehi _30646__1982 (.L_HI(net1982));
 sg13g2_tiehi _28510__1983 (.L_HI(net1983));
 sg13g2_tiehi _28509__1984 (.L_HI(net1984));
 sg13g2_tiehi _28508__1985 (.L_HI(net1985));
 sg13g2_tiehi _28507__1986 (.L_HI(net1986));
 sg13g2_tiehi _28506__1987 (.L_HI(net1987));
 sg13g2_tiehi _28505__1988 (.L_HI(net1988));
 sg13g2_tiehi _28504__1989 (.L_HI(net1989));
 sg13g2_tiehi _28503__1990 (.L_HI(net1990));
 sg13g2_tiehi _28502__1991 (.L_HI(net1991));
 sg13g2_tiehi _28501__1992 (.L_HI(net1992));
 sg13g2_tiehi _28500__1993 (.L_HI(net1993));
 sg13g2_tiehi _28499__1994 (.L_HI(net1994));
 sg13g2_tiehi _28498__1995 (.L_HI(net1995));
 sg13g2_tiehi _28497__1996 (.L_HI(net1996));
 sg13g2_tiehi _28496__1997 (.L_HI(net1997));
 sg13g2_tiehi _28495__1998 (.L_HI(net1998));
 sg13g2_tiehi _28494__1999 (.L_HI(net1999));
 sg13g2_tiehi _28493__2000 (.L_HI(net2000));
 sg13g2_tiehi _28492__2001 (.L_HI(net2001));
 sg13g2_tiehi _28491__2002 (.L_HI(net2002));
 sg13g2_tiehi _28490__2003 (.L_HI(net2003));
 sg13g2_tiehi _28489__2004 (.L_HI(net2004));
 sg13g2_tiehi _28488__2005 (.L_HI(net2005));
 sg13g2_tiehi _28487__2006 (.L_HI(net2006));
 sg13g2_tiehi _28486__2007 (.L_HI(net2007));
 sg13g2_tiehi _28485__2008 (.L_HI(net2008));
 sg13g2_tiehi _28484__2009 (.L_HI(net2009));
 sg13g2_tiehi _28483__2010 (.L_HI(net2010));
 sg13g2_tiehi _28482__2011 (.L_HI(net2011));
 sg13g2_tiehi _28481__2012 (.L_HI(net2012));
 sg13g2_tiehi _28480__2013 (.L_HI(net2013));
 sg13g2_tiehi _28479__2014 (.L_HI(net2014));
 sg13g2_tiehi _28478__2015 (.L_HI(net2015));
 sg13g2_tiehi _28477__2016 (.L_HI(net2016));
 sg13g2_tiehi _28476__2017 (.L_HI(net2017));
 sg13g2_tiehi _28475__2018 (.L_HI(net2018));
 sg13g2_tiehi _28474__2019 (.L_HI(net2019));
 sg13g2_tiehi _28473__2020 (.L_HI(net2020));
 sg13g2_tiehi _28472__2021 (.L_HI(net2021));
 sg13g2_tiehi _28471__2022 (.L_HI(net2022));
 sg13g2_tiehi _28470__2023 (.L_HI(net2023));
 sg13g2_tiehi _28469__2024 (.L_HI(net2024));
 sg13g2_tiehi _28468__2025 (.L_HI(net2025));
 sg13g2_tiehi _28467__2026 (.L_HI(net2026));
 sg13g2_tiehi _28466__2027 (.L_HI(net2027));
 sg13g2_tiehi _28465__2028 (.L_HI(net2028));
 sg13g2_tiehi _28464__2029 (.L_HI(net2029));
 sg13g2_tiehi _28463__2030 (.L_HI(net2030));
 sg13g2_tiehi _28462__2031 (.L_HI(net2031));
 sg13g2_tiehi _28461__2032 (.L_HI(net2032));
 sg13g2_tiehi _28460__2033 (.L_HI(net2033));
 sg13g2_tiehi _28459__2034 (.L_HI(net2034));
 sg13g2_tiehi _28458__2035 (.L_HI(net2035));
 sg13g2_tiehi _28457__2036 (.L_HI(net2036));
 sg13g2_tiehi _28456__2037 (.L_HI(net2037));
 sg13g2_tiehi _28455__2038 (.L_HI(net2038));
 sg13g2_tiehi _28454__2039 (.L_HI(net2039));
 sg13g2_tiehi _28453__2040 (.L_HI(net2040));
 sg13g2_tiehi _28452__2041 (.L_HI(net2041));
 sg13g2_tiehi _28451__2042 (.L_HI(net2042));
 sg13g2_tiehi _28450__2043 (.L_HI(net2043));
 sg13g2_tiehi _28449__2044 (.L_HI(net2044));
 sg13g2_tiehi _28448__2045 (.L_HI(net2045));
 sg13g2_tiehi _28447__2046 (.L_HI(net2046));
 sg13g2_tiehi _28446__2047 (.L_HI(net2047));
 sg13g2_tiehi _28445__2048 (.L_HI(net2048));
 sg13g2_tiehi _28444__2049 (.L_HI(net2049));
 sg13g2_tiehi _28443__2050 (.L_HI(net2050));
 sg13g2_tiehi _28442__2051 (.L_HI(net2051));
 sg13g2_tiehi _28441__2052 (.L_HI(net2052));
 sg13g2_tiehi _28440__2053 (.L_HI(net2053));
 sg13g2_tiehi _28439__2054 (.L_HI(net2054));
 sg13g2_tiehi _28438__2055 (.L_HI(net2055));
 sg13g2_tiehi _28437__2056 (.L_HI(net2056));
 sg13g2_tiehi _28436__2057 (.L_HI(net2057));
 sg13g2_tiehi _28435__2058 (.L_HI(net2058));
 sg13g2_tiehi _28434__2059 (.L_HI(net2059));
 sg13g2_tiehi _28433__2060 (.L_HI(net2060));
 sg13g2_tiehi _28432__2061 (.L_HI(net2061));
 sg13g2_tiehi _28431__2062 (.L_HI(net2062));
 sg13g2_tiehi _28430__2063 (.L_HI(net2063));
 sg13g2_tiehi _28429__2064 (.L_HI(net2064));
 sg13g2_tiehi _28428__2065 (.L_HI(net2065));
 sg13g2_tiehi _28427__2066 (.L_HI(net2066));
 sg13g2_tiehi _28426__2067 (.L_HI(net2067));
 sg13g2_tiehi _28425__2068 (.L_HI(net2068));
 sg13g2_tiehi _28424__2069 (.L_HI(net2069));
 sg13g2_tiehi _28423__2070 (.L_HI(net2070));
 sg13g2_tiehi _28422__2071 (.L_HI(net2071));
 sg13g2_tiehi _28421__2072 (.L_HI(net2072));
 sg13g2_tiehi _28420__2073 (.L_HI(net2073));
 sg13g2_tiehi _28419__2074 (.L_HI(net2074));
 sg13g2_tiehi _28418__2075 (.L_HI(net2075));
 sg13g2_tiehi _28417__2076 (.L_HI(net2076));
 sg13g2_tiehi _28416__2077 (.L_HI(net2077));
 sg13g2_tiehi _28415__2078 (.L_HI(net2078));
 sg13g2_tiehi _28414__2079 (.L_HI(net2079));
 sg13g2_tiehi _28413__2080 (.L_HI(net2080));
 sg13g2_tiehi _28412__2081 (.L_HI(net2081));
 sg13g2_tiehi _28411__2082 (.L_HI(net2082));
 sg13g2_tiehi _28410__2083 (.L_HI(net2083));
 sg13g2_tiehi _28409__2084 (.L_HI(net2084));
 sg13g2_tiehi _28408__2085 (.L_HI(net2085));
 sg13g2_tiehi _28407__2086 (.L_HI(net2086));
 sg13g2_tiehi _28406__2087 (.L_HI(net2087));
 sg13g2_tiehi _28405__2088 (.L_HI(net2088));
 sg13g2_tiehi _28404__2089 (.L_HI(net2089));
 sg13g2_tiehi _28403__2090 (.L_HI(net2090));
 sg13g2_tiehi _28402__2091 (.L_HI(net2091));
 sg13g2_tiehi _28401__2092 (.L_HI(net2092));
 sg13g2_tiehi _28400__2093 (.L_HI(net2093));
 sg13g2_tiehi _28399__2094 (.L_HI(net2094));
 sg13g2_tiehi _28398__2095 (.L_HI(net2095));
 sg13g2_tiehi _28397__2096 (.L_HI(net2096));
 sg13g2_tiehi _28396__2097 (.L_HI(net2097));
 sg13g2_tiehi _28395__2098 (.L_HI(net2098));
 sg13g2_tiehi _28394__2099 (.L_HI(net2099));
 sg13g2_tiehi _28393__2100 (.L_HI(net2100));
 sg13g2_tiehi _28392__2101 (.L_HI(net2101));
 sg13g2_tiehi _28391__2102 (.L_HI(net2102));
 sg13g2_tiehi _28390__2103 (.L_HI(net2103));
 sg13g2_tiehi _28389__2104 (.L_HI(net2104));
 sg13g2_tiehi _28388__2105 (.L_HI(net2105));
 sg13g2_tiehi _28387__2106 (.L_HI(net2106));
 sg13g2_tiehi _28386__2107 (.L_HI(net2107));
 sg13g2_tiehi _28385__2108 (.L_HI(net2108));
 sg13g2_tiehi _28384__2109 (.L_HI(net2109));
 sg13g2_tiehi _28383__2110 (.L_HI(net2110));
 sg13g2_tiehi _28382__2111 (.L_HI(net2111));
 sg13g2_tiehi _28381__2112 (.L_HI(net2112));
 sg13g2_tiehi _28380__2113 (.L_HI(net2113));
 sg13g2_tiehi _28379__2114 (.L_HI(net2114));
 sg13g2_tiehi _28378__2115 (.L_HI(net2115));
 sg13g2_tiehi _28377__2116 (.L_HI(net2116));
 sg13g2_tiehi _28376__2117 (.L_HI(net2117));
 sg13g2_tiehi _28375__2118 (.L_HI(net2118));
 sg13g2_tiehi _28374__2119 (.L_HI(net2119));
 sg13g2_tiehi _28373__2120 (.L_HI(net2120));
 sg13g2_tiehi _28372__2121 (.L_HI(net2121));
 sg13g2_tiehi _28371__2122 (.L_HI(net2122));
 sg13g2_tiehi _28370__2123 (.L_HI(net2123));
 sg13g2_tiehi _28369__2124 (.L_HI(net2124));
 sg13g2_tiehi _28368__2125 (.L_HI(net2125));
 sg13g2_tiehi _28367__2126 (.L_HI(net2126));
 sg13g2_tiehi _28366__2127 (.L_HI(net2127));
 sg13g2_tiehi _28365__2128 (.L_HI(net2128));
 sg13g2_tiehi _28364__2129 (.L_HI(net2129));
 sg13g2_tiehi _28363__2130 (.L_HI(net2130));
 sg13g2_tiehi _28362__2131 (.L_HI(net2131));
 sg13g2_tiehi _28361__2132 (.L_HI(net2132));
 sg13g2_tiehi _28360__2133 (.L_HI(net2133));
 sg13g2_tiehi _28359__2134 (.L_HI(net2134));
 sg13g2_tiehi _28358__2135 (.L_HI(net2135));
 sg13g2_tiehi _28357__2136 (.L_HI(net2136));
 sg13g2_tiehi _28356__2137 (.L_HI(net2137));
 sg13g2_tiehi _28355__2138 (.L_HI(net2138));
 sg13g2_tiehi _28354__2139 (.L_HI(net2139));
 sg13g2_tiehi _28353__2140 (.L_HI(net2140));
 sg13g2_tiehi _28352__2141 (.L_HI(net2141));
 sg13g2_tiehi _28351__2142 (.L_HI(net2142));
 sg13g2_tiehi _28350__2143 (.L_HI(net2143));
 sg13g2_tiehi _28349__2144 (.L_HI(net2144));
 sg13g2_tiehi _28348__2145 (.L_HI(net2145));
 sg13g2_tiehi _28347__2146 (.L_HI(net2146));
 sg13g2_tiehi _28346__2147 (.L_HI(net2147));
 sg13g2_tiehi _28345__2148 (.L_HI(net2148));
 sg13g2_tiehi _28344__2149 (.L_HI(net2149));
 sg13g2_tiehi _28343__2150 (.L_HI(net2150));
 sg13g2_tiehi _28342__2151 (.L_HI(net2151));
 sg13g2_tiehi _28341__2152 (.L_HI(net2152));
 sg13g2_tiehi _28340__2153 (.L_HI(net2153));
 sg13g2_tiehi _28339__2154 (.L_HI(net2154));
 sg13g2_tiehi _28338__2155 (.L_HI(net2155));
 sg13g2_tiehi _28337__2156 (.L_HI(net2156));
 sg13g2_tiehi _28336__2157 (.L_HI(net2157));
 sg13g2_tiehi _28335__2158 (.L_HI(net2158));
 sg13g2_tiehi _28334__2159 (.L_HI(net2159));
 sg13g2_tiehi _28333__2160 (.L_HI(net2160));
 sg13g2_tiehi _28332__2161 (.L_HI(net2161));
 sg13g2_tiehi _28331__2162 (.L_HI(net2162));
 sg13g2_tiehi _28330__2163 (.L_HI(net2163));
 sg13g2_tiehi _28329__2164 (.L_HI(net2164));
 sg13g2_tiehi _28328__2165 (.L_HI(net2165));
 sg13g2_tiehi _28327__2166 (.L_HI(net2166));
 sg13g2_tiehi _28326__2167 (.L_HI(net2167));
 sg13g2_tiehi _28325__2168 (.L_HI(net2168));
 sg13g2_tiehi _28324__2169 (.L_HI(net2169));
 sg13g2_tiehi _28323__2170 (.L_HI(net2170));
 sg13g2_tiehi _28322__2171 (.L_HI(net2171));
 sg13g2_tiehi _28321__2172 (.L_HI(net2172));
 sg13g2_tiehi _28320__2173 (.L_HI(net2173));
 sg13g2_tiehi _28319__2174 (.L_HI(net2174));
 sg13g2_tiehi _28318__2175 (.L_HI(net2175));
 sg13g2_tiehi _28317__2176 (.L_HI(net2176));
 sg13g2_tiehi _28316__2177 (.L_HI(net2177));
 sg13g2_tiehi _28315__2178 (.L_HI(net2178));
 sg13g2_tiehi _28314__2179 (.L_HI(net2179));
 sg13g2_tiehi _28313__2180 (.L_HI(net2180));
 sg13g2_tiehi _28312__2181 (.L_HI(net2181));
 sg13g2_tiehi _28311__2182 (.L_HI(net2182));
 sg13g2_tiehi _28310__2183 (.L_HI(net2183));
 sg13g2_tiehi _28309__2184 (.L_HI(net2184));
 sg13g2_tiehi _28308__2185 (.L_HI(net2185));
 sg13g2_tiehi _28307__2186 (.L_HI(net2186));
 sg13g2_tiehi _28306__2187 (.L_HI(net2187));
 sg13g2_tiehi _28305__2188 (.L_HI(net2188));
 sg13g2_tiehi _28304__2189 (.L_HI(net2189));
 sg13g2_tiehi _28303__2190 (.L_HI(net2190));
 sg13g2_tiehi _28302__2191 (.L_HI(net2191));
 sg13g2_tiehi _28301__2192 (.L_HI(net2192));
 sg13g2_tiehi _28300__2193 (.L_HI(net2193));
 sg13g2_tiehi _28299__2194 (.L_HI(net2194));
 sg13g2_tiehi _28298__2195 (.L_HI(net2195));
 sg13g2_tiehi _28297__2196 (.L_HI(net2196));
 sg13g2_tiehi _28296__2197 (.L_HI(net2197));
 sg13g2_tiehi _28295__2198 (.L_HI(net2198));
 sg13g2_tiehi _28294__2199 (.L_HI(net2199));
 sg13g2_tiehi _28293__2200 (.L_HI(net2200));
 sg13g2_tiehi _28292__2201 (.L_HI(net2201));
 sg13g2_tiehi _28291__2202 (.L_HI(net2202));
 sg13g2_tiehi _28290__2203 (.L_HI(net2203));
 sg13g2_tiehi _28289__2204 (.L_HI(net2204));
 sg13g2_tiehi _28288__2205 (.L_HI(net2205));
 sg13g2_tiehi _28287__2206 (.L_HI(net2206));
 sg13g2_tiehi _28286__2207 (.L_HI(net2207));
 sg13g2_tiehi _28285__2208 (.L_HI(net2208));
 sg13g2_tiehi _28284__2209 (.L_HI(net2209));
 sg13g2_tiehi _28283__2210 (.L_HI(net2210));
 sg13g2_tiehi _28282__2211 (.L_HI(net2211));
 sg13g2_tiehi _28281__2212 (.L_HI(net2212));
 sg13g2_tiehi _28280__2213 (.L_HI(net2213));
 sg13g2_tiehi _28279__2214 (.L_HI(net2214));
 sg13g2_tiehi _28278__2215 (.L_HI(net2215));
 sg13g2_tiehi _28277__2216 (.L_HI(net2216));
 sg13g2_tiehi _28276__2217 (.L_HI(net2217));
 sg13g2_tiehi _28275__2218 (.L_HI(net2218));
 sg13g2_tiehi _28274__2219 (.L_HI(net2219));
 sg13g2_tiehi _28273__2220 (.L_HI(net2220));
 sg13g2_tiehi _28272__2221 (.L_HI(net2221));
 sg13g2_tiehi _28271__2222 (.L_HI(net2222));
 sg13g2_tiehi _28270__2223 (.L_HI(net2223));
 sg13g2_tiehi _28269__2224 (.L_HI(net2224));
 sg13g2_tiehi _28268__2225 (.L_HI(net2225));
 sg13g2_tiehi _28267__2226 (.L_HI(net2226));
 sg13g2_tiehi _28266__2227 (.L_HI(net2227));
 sg13g2_tiehi _28265__2228 (.L_HI(net2228));
 sg13g2_tiehi _28264__2229 (.L_HI(net2229));
 sg13g2_tiehi _28263__2230 (.L_HI(net2230));
 sg13g2_tiehi _28262__2231 (.L_HI(net2231));
 sg13g2_tiehi _28261__2232 (.L_HI(net2232));
 sg13g2_tiehi _28260__2233 (.L_HI(net2233));
 sg13g2_tiehi _28259__2234 (.L_HI(net2234));
 sg13g2_tiehi _28258__2235 (.L_HI(net2235));
 sg13g2_tiehi _28257__2236 (.L_HI(net2236));
 sg13g2_tiehi _28256__2237 (.L_HI(net2237));
 sg13g2_tiehi _28255__2238 (.L_HI(net2238));
 sg13g2_tiehi _28254__2239 (.L_HI(net2239));
 sg13g2_tiehi _28253__2240 (.L_HI(net2240));
 sg13g2_tiehi _28252__2241 (.L_HI(net2241));
 sg13g2_tiehi _28251__2242 (.L_HI(net2242));
 sg13g2_tiehi _28250__2243 (.L_HI(net2243));
 sg13g2_tiehi _28249__2244 (.L_HI(net2244));
 sg13g2_tiehi _28248__2245 (.L_HI(net2245));
 sg13g2_tiehi _28247__2246 (.L_HI(net2246));
 sg13g2_tiehi _28246__2247 (.L_HI(net2247));
 sg13g2_tiehi _28245__2248 (.L_HI(net2248));
 sg13g2_tiehi _28244__2249 (.L_HI(net2249));
 sg13g2_tiehi _28243__2250 (.L_HI(net2250));
 sg13g2_tiehi _28242__2251 (.L_HI(net2251));
 sg13g2_tiehi _28241__2252 (.L_HI(net2252));
 sg13g2_tiehi _28240__2253 (.L_HI(net2253));
 sg13g2_tiehi _28239__2254 (.L_HI(net2254));
 sg13g2_tiehi _28238__2255 (.L_HI(net2255));
 sg13g2_tiehi _28237__2256 (.L_HI(net2256));
 sg13g2_tiehi _28236__2257 (.L_HI(net2257));
 sg13g2_tiehi _28235__2258 (.L_HI(net2258));
 sg13g2_tiehi _28234__2259 (.L_HI(net2259));
 sg13g2_tiehi _28233__2260 (.L_HI(net2260));
 sg13g2_tiehi _28232__2261 (.L_HI(net2261));
 sg13g2_tiehi _28231__2262 (.L_HI(net2262));
 sg13g2_tiehi _28230__2263 (.L_HI(net2263));
 sg13g2_tiehi _28229__2264 (.L_HI(net2264));
 sg13g2_tiehi _28228__2265 (.L_HI(net2265));
 sg13g2_tiehi _28227__2266 (.L_HI(net2266));
 sg13g2_tiehi _28226__2267 (.L_HI(net2267));
 sg13g2_tiehi _28225__2268 (.L_HI(net2268));
 sg13g2_tiehi _28224__2269 (.L_HI(net2269));
 sg13g2_tiehi _28223__2270 (.L_HI(net2270));
 sg13g2_tiehi _28222__2271 (.L_HI(net2271));
 sg13g2_tiehi _28221__2272 (.L_HI(net2272));
 sg13g2_tiehi _28220__2273 (.L_HI(net2273));
 sg13g2_tiehi _28219__2274 (.L_HI(net2274));
 sg13g2_tiehi _28218__2275 (.L_HI(net2275));
 sg13g2_tiehi _28217__2276 (.L_HI(net2276));
 sg13g2_tiehi _28216__2277 (.L_HI(net2277));
 sg13g2_tiehi _28215__2278 (.L_HI(net2278));
 sg13g2_tiehi _28214__2279 (.L_HI(net2279));
 sg13g2_tiehi _28213__2280 (.L_HI(net2280));
 sg13g2_tiehi _28212__2281 (.L_HI(net2281));
 sg13g2_tiehi _28211__2282 (.L_HI(net2282));
 sg13g2_tiehi _28210__2283 (.L_HI(net2283));
 sg13g2_tiehi _28209__2284 (.L_HI(net2284));
 sg13g2_tiehi _28208__2285 (.L_HI(net2285));
 sg13g2_tiehi _28207__2286 (.L_HI(net2286));
 sg13g2_tiehi _28206__2287 (.L_HI(net2287));
 sg13g2_tiehi _28205__2288 (.L_HI(net2288));
 sg13g2_tiehi _28204__2289 (.L_HI(net2289));
 sg13g2_tiehi _28203__2290 (.L_HI(net2290));
 sg13g2_tiehi _28202__2291 (.L_HI(net2291));
 sg13g2_tiehi _28201__2292 (.L_HI(net2292));
 sg13g2_tiehi _28200__2293 (.L_HI(net2293));
 sg13g2_tiehi _28199__2294 (.L_HI(net2294));
 sg13g2_tiehi _28198__2295 (.L_HI(net2295));
 sg13g2_tiehi _28197__2296 (.L_HI(net2296));
 sg13g2_tiehi _28196__2297 (.L_HI(net2297));
 sg13g2_tiehi _28195__2298 (.L_HI(net2298));
 sg13g2_tiehi _28194__2299 (.L_HI(net2299));
 sg13g2_tiehi _28193__2300 (.L_HI(net2300));
 sg13g2_tiehi _28192__2301 (.L_HI(net2301));
 sg13g2_tiehi _28191__2302 (.L_HI(net2302));
 sg13g2_tiehi _28190__2303 (.L_HI(net2303));
 sg13g2_tiehi _28189__2304 (.L_HI(net2304));
 sg13g2_tiehi _28188__2305 (.L_HI(net2305));
 sg13g2_tiehi _28187__2306 (.L_HI(net2306));
 sg13g2_tiehi _28186__2307 (.L_HI(net2307));
 sg13g2_tiehi _28185__2308 (.L_HI(net2308));
 sg13g2_tiehi _28184__2309 (.L_HI(net2309));
 sg13g2_tiehi _28183__2310 (.L_HI(net2310));
 sg13g2_tiehi _28182__2311 (.L_HI(net2311));
 sg13g2_tiehi _28181__2312 (.L_HI(net2312));
 sg13g2_tiehi _28180__2313 (.L_HI(net2313));
 sg13g2_tiehi _28179__2314 (.L_HI(net2314));
 sg13g2_tiehi _28178__2315 (.L_HI(net2315));
 sg13g2_tiehi _28177__2316 (.L_HI(net2316));
 sg13g2_tiehi _28176__2317 (.L_HI(net2317));
 sg13g2_tiehi _28175__2318 (.L_HI(net2318));
 sg13g2_tiehi _28174__2319 (.L_HI(net2319));
 sg13g2_tiehi _28173__2320 (.L_HI(net2320));
 sg13g2_tiehi _28172__2321 (.L_HI(net2321));
 sg13g2_tiehi _28171__2322 (.L_HI(net2322));
 sg13g2_tiehi _28170__2323 (.L_HI(net2323));
 sg13g2_tiehi _28169__2324 (.L_HI(net2324));
 sg13g2_tiehi _28168__2325 (.L_HI(net2325));
 sg13g2_tiehi _28167__2326 (.L_HI(net2326));
 sg13g2_tiehi _28166__2327 (.L_HI(net2327));
 sg13g2_tiehi _28165__2328 (.L_HI(net2328));
 sg13g2_tiehi _28164__2329 (.L_HI(net2329));
 sg13g2_tiehi _28163__2330 (.L_HI(net2330));
 sg13g2_tiehi _28162__2331 (.L_HI(net2331));
 sg13g2_tiehi _28161__2332 (.L_HI(net2332));
 sg13g2_tiehi _28160__2333 (.L_HI(net2333));
 sg13g2_tiehi _28159__2334 (.L_HI(net2334));
 sg13g2_tiehi _28158__2335 (.L_HI(net2335));
 sg13g2_tiehi _28157__2336 (.L_HI(net2336));
 sg13g2_tiehi _28156__2337 (.L_HI(net2337));
 sg13g2_tiehi _28155__2338 (.L_HI(net2338));
 sg13g2_tiehi _28154__2339 (.L_HI(net2339));
 sg13g2_tiehi _28153__2340 (.L_HI(net2340));
 sg13g2_tiehi _28152__2341 (.L_HI(net2341));
 sg13g2_tiehi _28151__2342 (.L_HI(net2342));
 sg13g2_tiehi _28150__2343 (.L_HI(net2343));
 sg13g2_tiehi _28149__2344 (.L_HI(net2344));
 sg13g2_tiehi _28148__2345 (.L_HI(net2345));
 sg13g2_tiehi _28147__2346 (.L_HI(net2346));
 sg13g2_tiehi _28146__2347 (.L_HI(net2347));
 sg13g2_tiehi _28145__2348 (.L_HI(net2348));
 sg13g2_tiehi _28144__2349 (.L_HI(net2349));
 sg13g2_tiehi _28143__2350 (.L_HI(net2350));
 sg13g2_tiehi _28142__2351 (.L_HI(net2351));
 sg13g2_tiehi _28141__2352 (.L_HI(net2352));
 sg13g2_tiehi _28140__2353 (.L_HI(net2353));
 sg13g2_tiehi _28139__2354 (.L_HI(net2354));
 sg13g2_tiehi _28138__2355 (.L_HI(net2355));
 sg13g2_tiehi _28137__2356 (.L_HI(net2356));
 sg13g2_tiehi _28136__2357 (.L_HI(net2357));
 sg13g2_tiehi _28135__2358 (.L_HI(net2358));
 sg13g2_tiehi _28134__2359 (.L_HI(net2359));
 sg13g2_tiehi _28133__2360 (.L_HI(net2360));
 sg13g2_tiehi _28132__2361 (.L_HI(net2361));
 sg13g2_tiehi _28131__2362 (.L_HI(net2362));
 sg13g2_tiehi _28130__2363 (.L_HI(net2363));
 sg13g2_tiehi _28129__2364 (.L_HI(net2364));
 sg13g2_tiehi _28128__2365 (.L_HI(net2365));
 sg13g2_tiehi _28127__2366 (.L_HI(net2366));
 sg13g2_tiehi _28126__2367 (.L_HI(net2367));
 sg13g2_tiehi _28125__2368 (.L_HI(net2368));
 sg13g2_tiehi _28124__2369 (.L_HI(net2369));
 sg13g2_tiehi _28123__2370 (.L_HI(net2370));
 sg13g2_tiehi _28122__2371 (.L_HI(net2371));
 sg13g2_tiehi _28121__2372 (.L_HI(net2372));
 sg13g2_tiehi _28120__2373 (.L_HI(net2373));
 sg13g2_tiehi _28119__2374 (.L_HI(net2374));
 sg13g2_tiehi _28118__2375 (.L_HI(net2375));
 sg13g2_tiehi _28117__2376 (.L_HI(net2376));
 sg13g2_tiehi _28116__2377 (.L_HI(net2377));
 sg13g2_tiehi _28115__2378 (.L_HI(net2378));
 sg13g2_tiehi _28114__2379 (.L_HI(net2379));
 sg13g2_tiehi _28113__2380 (.L_HI(net2380));
 sg13g2_tiehi _28112__2381 (.L_HI(net2381));
 sg13g2_tiehi _28111__2382 (.L_HI(net2382));
 sg13g2_tiehi _28110__2383 (.L_HI(net2383));
 sg13g2_tiehi _28109__2384 (.L_HI(net2384));
 sg13g2_tiehi _28108__2385 (.L_HI(net2385));
 sg13g2_tiehi _28107__2386 (.L_HI(net2386));
 sg13g2_tiehi _28106__2387 (.L_HI(net2387));
 sg13g2_tiehi _28105__2388 (.L_HI(net2388));
 sg13g2_tiehi _28104__2389 (.L_HI(net2389));
 sg13g2_tiehi _28103__2390 (.L_HI(net2390));
 sg13g2_tiehi _28102__2391 (.L_HI(net2391));
 sg13g2_tiehi _28101__2392 (.L_HI(net2392));
 sg13g2_tiehi _28100__2393 (.L_HI(net2393));
 sg13g2_tiehi _28099__2394 (.L_HI(net2394));
 sg13g2_tiehi _28098__2395 (.L_HI(net2395));
 sg13g2_tiehi _28097__2396 (.L_HI(net2396));
 sg13g2_tiehi _28096__2397 (.L_HI(net2397));
 sg13g2_tiehi _28095__2398 (.L_HI(net2398));
 sg13g2_tiehi _28094__2399 (.L_HI(net2399));
 sg13g2_tiehi _28093__2400 (.L_HI(net2400));
 sg13g2_tiehi _28092__2401 (.L_HI(net2401));
 sg13g2_tiehi _28091__2402 (.L_HI(net2402));
 sg13g2_tiehi _28090__2403 (.L_HI(net2403));
 sg13g2_tiehi _28089__2404 (.L_HI(net2404));
 sg13g2_tiehi _28088__2405 (.L_HI(net2405));
 sg13g2_tiehi _28087__2406 (.L_HI(net2406));
 sg13g2_tiehi _28086__2407 (.L_HI(net2407));
 sg13g2_tiehi _28085__2408 (.L_HI(net2408));
 sg13g2_tiehi _28084__2409 (.L_HI(net2409));
 sg13g2_tiehi _28083__2410 (.L_HI(net2410));
 sg13g2_tiehi _28082__2411 (.L_HI(net2411));
 sg13g2_tiehi _28081__2412 (.L_HI(net2412));
 sg13g2_tiehi _28080__2413 (.L_HI(net2413));
 sg13g2_tiehi _28079__2414 (.L_HI(net2414));
 sg13g2_tiehi _28078__2415 (.L_HI(net2415));
 sg13g2_tiehi _28077__2416 (.L_HI(net2416));
 sg13g2_tiehi _28076__2417 (.L_HI(net2417));
 sg13g2_tiehi _28075__2418 (.L_HI(net2418));
 sg13g2_tiehi _28074__2419 (.L_HI(net2419));
 sg13g2_tiehi _28073__2420 (.L_HI(net2420));
 sg13g2_tiehi _28064__2421 (.L_HI(net2421));
 sg13g2_tiehi _28063__2422 (.L_HI(net2422));
 sg13g2_tiehi _28062__2423 (.L_HI(net2423));
 sg13g2_tiehi _28061__2424 (.L_HI(net2424));
 sg13g2_tiehi _28060__2425 (.L_HI(net2425));
 sg13g2_tiehi _28059__2426 (.L_HI(net2426));
 sg13g2_tiehi _28058__2427 (.L_HI(net2427));
 sg13g2_tiehi _28057__2428 (.L_HI(net2428));
 sg13g2_tiehi _28056__2429 (.L_HI(net2429));
 sg13g2_tiehi _28055__2430 (.L_HI(net2430));
 sg13g2_tiehi _28054__2431 (.L_HI(net2431));
 sg13g2_tiehi _28053__2432 (.L_HI(net2432));
 sg13g2_tiehi _28052__2433 (.L_HI(net2433));
 sg13g2_tiehi _28051__2434 (.L_HI(net2434));
 sg13g2_tiehi _28050__2435 (.L_HI(net2435));
 sg13g2_tiehi _28049__2436 (.L_HI(net2436));
 sg13g2_tiehi _28048__2437 (.L_HI(net2437));
 sg13g2_tiehi _28047__2438 (.L_HI(net2438));
 sg13g2_tiehi _28046__2439 (.L_HI(net2439));
 sg13g2_tiehi _28045__2440 (.L_HI(net2440));
 sg13g2_tiehi _28044__2441 (.L_HI(net2441));
 sg13g2_tiehi _28043__2442 (.L_HI(net2442));
 sg13g2_tiehi _28042__2443 (.L_HI(net2443));
 sg13g2_tiehi _28041__2444 (.L_HI(net2444));
 sg13g2_tiehi _28040__2445 (.L_HI(net2445));
 sg13g2_tiehi _28039__2446 (.L_HI(net2446));
 sg13g2_tiehi _28038__2447 (.L_HI(net2447));
 sg13g2_tiehi _28037__2448 (.L_HI(net2448));
 sg13g2_tiehi _28036__2449 (.L_HI(net2449));
 sg13g2_tiehi _28035__2450 (.L_HI(net2450));
 sg13g2_tiehi _28034__2451 (.L_HI(net2451));
 sg13g2_tiehi _28033__2452 (.L_HI(net2452));
 sg13g2_tiehi _28032__2453 (.L_HI(net2453));
 sg13g2_tiehi _28031__2454 (.L_HI(net2454));
 sg13g2_tiehi _28030__2455 (.L_HI(net2455));
 sg13g2_tiehi _28029__2456 (.L_HI(net2456));
 sg13g2_tiehi _28028__2457 (.L_HI(net2457));
 sg13g2_tiehi _28027__2458 (.L_HI(net2458));
 sg13g2_tiehi _28026__2459 (.L_HI(net2459));
 sg13g2_tiehi _28025__2460 (.L_HI(net2460));
 sg13g2_tiehi _28024__2461 (.L_HI(net2461));
 sg13g2_tiehi _28023__2462 (.L_HI(net2462));
 sg13g2_tiehi _28022__2463 (.L_HI(net2463));
 sg13g2_tiehi _28021__2464 (.L_HI(net2464));
 sg13g2_tiehi _28020__2465 (.L_HI(net2465));
 sg13g2_tiehi _28019__2466 (.L_HI(net2466));
 sg13g2_tiehi _28018__2467 (.L_HI(net2467));
 sg13g2_tiehi _28017__2468 (.L_HI(net2468));
 sg13g2_tiehi _28016__2469 (.L_HI(net2469));
 sg13g2_tiehi _28015__2470 (.L_HI(net2470));
 sg13g2_tiehi _28014__2471 (.L_HI(net2471));
 sg13g2_tiehi _28013__2472 (.L_HI(net2472));
 sg13g2_tiehi _28012__2473 (.L_HI(net2473));
 sg13g2_tiehi _28011__2474 (.L_HI(net2474));
 sg13g2_tiehi _28010__2475 (.L_HI(net2475));
 sg13g2_tiehi _28009__2476 (.L_HI(net2476));
 sg13g2_tiehi _28008__2477 (.L_HI(net2477));
 sg13g2_tiehi _28007__2478 (.L_HI(net2478));
 sg13g2_tiehi _28006__2479 (.L_HI(net2479));
 sg13g2_tiehi _28005__2480 (.L_HI(net2480));
 sg13g2_tiehi _28004__2481 (.L_HI(net2481));
 sg13g2_tiehi _28003__2482 (.L_HI(net2482));
 sg13g2_tiehi _28002__2483 (.L_HI(net2483));
 sg13g2_tiehi _28001__2484 (.L_HI(net2484));
 sg13g2_tiehi _28000__2485 (.L_HI(net2485));
 sg13g2_tiehi _27999__2486 (.L_HI(net2486));
 sg13g2_tiehi _27998__2487 (.L_HI(net2487));
 sg13g2_tiehi _27997__2488 (.L_HI(net2488));
 sg13g2_tiehi _27996__2489 (.L_HI(net2489));
 sg13g2_tiehi _27995__2490 (.L_HI(net2490));
 sg13g2_tiehi _27994__2491 (.L_HI(net2491));
 sg13g2_tiehi _27993__2492 (.L_HI(net2492));
 sg13g2_tiehi _27992__2493 (.L_HI(net2493));
 sg13g2_tiehi _27991__2494 (.L_HI(net2494));
 sg13g2_tiehi _27990__2495 (.L_HI(net2495));
 sg13g2_tiehi _27989__2496 (.L_HI(net2496));
 sg13g2_tiehi _27988__2497 (.L_HI(net2497));
 sg13g2_tiehi _27987__2498 (.L_HI(net2498));
 sg13g2_tiehi _27986__2499 (.L_HI(net2499));
 sg13g2_tiehi _27978__2500 (.L_HI(net2500));
 sg13g2_tiehi _27977__2501 (.L_HI(net2501));
 sg13g2_tiehi _27976__2502 (.L_HI(net2502));
 sg13g2_tiehi _27975__2503 (.L_HI(net2503));
 sg13g2_tiehi _27974__2504 (.L_HI(net2504));
 sg13g2_tiehi _27973__2505 (.L_HI(net2505));
 sg13g2_tiehi _27972__2506 (.L_HI(net2506));
 sg13g2_tiehi _27971__2507 (.L_HI(net2507));
 sg13g2_tiehi _27970__2508 (.L_HI(net2508));
 sg13g2_tiehi _27969__2509 (.L_HI(net2509));
 sg13g2_tiehi _27968__2510 (.L_HI(net2510));
 sg13g2_tiehi _27967__2511 (.L_HI(net2511));
 sg13g2_tiehi _27966__2512 (.L_HI(net2512));
 sg13g2_tiehi _27965__2513 (.L_HI(net2513));
 sg13g2_tiehi _27964__2514 (.L_HI(net2514));
 sg13g2_tiehi _27963__2515 (.L_HI(net2515));
 sg13g2_tiehi _27962__2516 (.L_HI(net2516));
 sg13g2_tiehi _27961__2517 (.L_HI(net2517));
 sg13g2_tiehi _27960__2518 (.L_HI(net2518));
 sg13g2_tiehi _27959__2519 (.L_HI(net2519));
 sg13g2_tiehi _27958__2520 (.L_HI(net2520));
 sg13g2_tiehi _27957__2521 (.L_HI(net2521));
 sg13g2_tiehi _27956__2522 (.L_HI(net2522));
 sg13g2_tiehi _27955__2523 (.L_HI(net2523));
 sg13g2_tiehi _27954__2524 (.L_HI(net2524));
 sg13g2_tiehi _27953__2525 (.L_HI(net2525));
 sg13g2_tiehi _27952__2526 (.L_HI(net2526));
 sg13g2_tiehi _27951__2527 (.L_HI(net2527));
 sg13g2_tiehi _27950__2528 (.L_HI(net2528));
 sg13g2_tiehi _27948__2529 (.L_HI(net2529));
 sg13g2_tiehi _27947__2530 (.L_HI(net2530));
 sg13g2_tiehi _27946__2531 (.L_HI(net2531));
 sg13g2_tiehi _27945__2532 (.L_HI(net2532));
 sg13g2_tiehi _27944__2533 (.L_HI(net2533));
 sg13g2_tiehi _27943__2534 (.L_HI(net2534));
 sg13g2_tiehi _27942__2535 (.L_HI(net2535));
 sg13g2_tiehi _27941__2536 (.L_HI(net2536));
 sg13g2_tiehi _27940__2537 (.L_HI(net2537));
 sg13g2_tiehi _27939__2538 (.L_HI(net2538));
 sg13g2_tiehi _27938__2539 (.L_HI(net2539));
 sg13g2_tiehi _27937__2540 (.L_HI(net2540));
 sg13g2_tiehi _27936__2541 (.L_HI(net2541));
 sg13g2_tiehi _27935__2542 (.L_HI(net2542));
 sg13g2_tiehi _27934__2543 (.L_HI(net2543));
 sg13g2_tiehi _27933__2544 (.L_HI(net2544));
 sg13g2_tiehi _27932__2545 (.L_HI(net2545));
 sg13g2_tiehi _27931__2546 (.L_HI(net2546));
 sg13g2_tiehi _27930__2547 (.L_HI(net2547));
 sg13g2_tiehi _27929__2548 (.L_HI(net2548));
 sg13g2_tiehi _27928__2549 (.L_HI(net2549));
 sg13g2_tiehi _27927__2550 (.L_HI(net2550));
 sg13g2_tiehi _27926__2551 (.L_HI(net2551));
 sg13g2_tiehi _27925__2552 (.L_HI(net2552));
 sg13g2_tiehi _27924__2553 (.L_HI(net2553));
 sg13g2_tiehi _27923__2554 (.L_HI(net2554));
 sg13g2_tiehi _27922__2555 (.L_HI(net2555));
 sg13g2_tiehi _27921__2556 (.L_HI(net2556));
 sg13g2_tiehi _27920__2557 (.L_HI(net2557));
 sg13g2_tiehi _27919__2558 (.L_HI(net2558));
 sg13g2_tiehi _27918__2559 (.L_HI(net2559));
 sg13g2_tiehi _27917__2560 (.L_HI(net2560));
 sg13g2_tiehi _27916__2561 (.L_HI(net2561));
 sg13g2_tiehi _27915__2562 (.L_HI(net2562));
 sg13g2_tiehi _27914__2563 (.L_HI(net2563));
 sg13g2_tiehi _27913__2564 (.L_HI(net2564));
 sg13g2_tiehi _27912__2565 (.L_HI(net2565));
 sg13g2_tiehi _27911__2566 (.L_HI(net2566));
 sg13g2_tiehi _27910__2567 (.L_HI(net2567));
 sg13g2_tiehi _27909__2568 (.L_HI(net2568));
 sg13g2_tiehi _27908__2569 (.L_HI(net2569));
 sg13g2_tiehi _27907__2570 (.L_HI(net2570));
 sg13g2_tiehi _27906__2571 (.L_HI(net2571));
 sg13g2_tiehi _27905__2572 (.L_HI(net2572));
 sg13g2_tiehi _27904__2573 (.L_HI(net2573));
 sg13g2_tiehi _27903__2574 (.L_HI(net2574));
 sg13g2_tiehi _27902__2575 (.L_HI(net2575));
 sg13g2_tiehi _27901__2576 (.L_HI(net2576));
 sg13g2_tiehi _27900__2577 (.L_HI(net2577));
 sg13g2_tiehi _27899__2578 (.L_HI(net2578));
 sg13g2_tiehi _27898__2579 (.L_HI(net2579));
 sg13g2_tiehi _27897__2580 (.L_HI(net2580));
 sg13g2_tiehi _27896__2581 (.L_HI(net2581));
 sg13g2_tiehi _27895__2582 (.L_HI(net2582));
 sg13g2_tiehi _27894__2583 (.L_HI(net2583));
 sg13g2_tiehi _27893__2584 (.L_HI(net2584));
 sg13g2_tiehi _27892__2585 (.L_HI(net2585));
 sg13g2_tiehi _27891__2586 (.L_HI(net2586));
 sg13g2_tiehi _27890__2587 (.L_HI(net2587));
 sg13g2_tiehi _27889__2588 (.L_HI(net2588));
 sg13g2_tiehi _27888__2589 (.L_HI(net2589));
 sg13g2_tiehi _27887__2590 (.L_HI(net2590));
 sg13g2_tiehi _27886__2591 (.L_HI(net2591));
 sg13g2_tiehi _27885__2592 (.L_HI(net2592));
 sg13g2_tiehi _27884__2593 (.L_HI(net2593));
 sg13g2_tiehi _27883__2594 (.L_HI(net2594));
 sg13g2_tiehi _27882__2595 (.L_HI(net2595));
 sg13g2_tiehi _27881__2596 (.L_HI(net2596));
 sg13g2_tiehi _27880__2597 (.L_HI(net2597));
 sg13g2_tiehi _27879__2598 (.L_HI(net2598));
 sg13g2_tiehi _27878__2599 (.L_HI(net2599));
 sg13g2_tiehi _27877__2600 (.L_HI(net2600));
 sg13g2_tiehi _27876__2601 (.L_HI(net2601));
 sg13g2_tiehi _27875__2602 (.L_HI(net2602));
 sg13g2_tiehi _27874__2603 (.L_HI(net2603));
 sg13g2_tiehi _27873__2604 (.L_HI(net2604));
 sg13g2_tiehi _27872__2605 (.L_HI(net2605));
 sg13g2_tiehi _27871__2606 (.L_HI(net2606));
 sg13g2_tiehi _27870__2607 (.L_HI(net2607));
 sg13g2_tiehi _27869__2608 (.L_HI(net2608));
 sg13g2_tiehi _27868__2609 (.L_HI(net2609));
 sg13g2_tiehi _27867__2610 (.L_HI(net2610));
 sg13g2_tiehi _27866__2611 (.L_HI(net2611));
 sg13g2_tiehi _27865__2612 (.L_HI(net2612));
 sg13g2_tiehi _27864__2613 (.L_HI(net2613));
 sg13g2_tiehi _27863__2614 (.L_HI(net2614));
 sg13g2_tiehi _27862__2615 (.L_HI(net2615));
 sg13g2_tiehi _27861__2616 (.L_HI(net2616));
 sg13g2_tiehi _27858__2617 (.L_HI(net2617));
 sg13g2_tiehi _27857__2618 (.L_HI(net2618));
 sg13g2_tiehi _27856__2619 (.L_HI(net2619));
 sg13g2_tiehi _27855__2620 (.L_HI(net2620));
 sg13g2_tiehi _27854__2621 (.L_HI(net2621));
 sg13g2_tiehi _27853__2622 (.L_HI(net2622));
 sg13g2_tiehi _27852__2623 (.L_HI(net2623));
 sg13g2_tiehi _27851__2624 (.L_HI(net2624));
 sg13g2_tiehi _27850__2625 (.L_HI(net2625));
 sg13g2_tiehi _27849__2626 (.L_HI(net2626));
 sg13g2_tiehi _27848__2627 (.L_HI(net2627));
 sg13g2_tiehi _27847__2628 (.L_HI(net2628));
 sg13g2_tiehi _27846__2629 (.L_HI(net2629));
 sg13g2_tiehi _27845__2630 (.L_HI(net2630));
 sg13g2_tiehi _27844__2631 (.L_HI(net2631));
 sg13g2_tiehi _27843__2632 (.L_HI(net2632));
 sg13g2_tiehi _27842__2633 (.L_HI(net2633));
 sg13g2_tiehi _27841__2634 (.L_HI(net2634));
 sg13g2_tiehi _27840__2635 (.L_HI(net2635));
 sg13g2_tiehi _27839__2636 (.L_HI(net2636));
 sg13g2_tiehi _27838__2637 (.L_HI(net2637));
 sg13g2_tiehi _27837__2638 (.L_HI(net2638));
 sg13g2_tiehi _27836__2639 (.L_HI(net2639));
 sg13g2_tiehi _27835__2640 (.L_HI(net2640));
 sg13g2_tiehi _27834__2641 (.L_HI(net2641));
 sg13g2_tiehi _27833__2642 (.L_HI(net2642));
 sg13g2_tiehi _27832__2643 (.L_HI(net2643));
 sg13g2_tiehi _27831__2644 (.L_HI(net2644));
 sg13g2_tiehi _27830__2645 (.L_HI(net2645));
 sg13g2_tiehi _27829__2646 (.L_HI(net2646));
 sg13g2_tiehi _27828__2647 (.L_HI(net2647));
 sg13g2_tiehi _27827__2648 (.L_HI(net2648));
 sg13g2_tiehi _27826__2649 (.L_HI(net2649));
 sg13g2_tiehi _27825__2650 (.L_HI(net2650));
 sg13g2_tiehi _27824__2651 (.L_HI(net2651));
 sg13g2_tiehi _27823__2652 (.L_HI(net2652));
 sg13g2_tiehi _27822__2653 (.L_HI(net2653));
 sg13g2_tiehi _27821__2654 (.L_HI(net2654));
 sg13g2_tiehi _27820__2655 (.L_HI(net2655));
 sg13g2_tiehi _27819__2656 (.L_HI(net2656));
 sg13g2_tiehi _27818__2657 (.L_HI(net2657));
 sg13g2_tiehi _27817__2658 (.L_HI(net2658));
 sg13g2_tiehi _27816__2659 (.L_HI(net2659));
 sg13g2_tiehi _27815__2660 (.L_HI(net2660));
 sg13g2_tiehi _27814__2661 (.L_HI(net2661));
 sg13g2_tiehi _27813__2662 (.L_HI(net2662));
 sg13g2_tiehi _27812__2663 (.L_HI(net2663));
 sg13g2_tiehi _27811__2664 (.L_HI(net2664));
 sg13g2_tiehi _27810__2665 (.L_HI(net2665));
 sg13g2_tiehi _27809__2666 (.L_HI(net2666));
 sg13g2_tiehi _27808__2667 (.L_HI(net2667));
 sg13g2_tiehi _27807__2668 (.L_HI(net2668));
 sg13g2_tiehi _27806__2669 (.L_HI(net2669));
 sg13g2_tiehi _27805__2670 (.L_HI(net2670));
 sg13g2_tiehi _27804__2671 (.L_HI(net2671));
 sg13g2_tiehi _27803__2672 (.L_HI(net2672));
 sg13g2_tiehi _27802__2673 (.L_HI(net2673));
 sg13g2_tiehi _27801__2674 (.L_HI(net2674));
 sg13g2_tiehi _27800__2675 (.L_HI(net2675));
 sg13g2_tiehi _27799__2676 (.L_HI(net2676));
 sg13g2_tiehi _27798__2677 (.L_HI(net2677));
 sg13g2_tiehi _27797__2678 (.L_HI(net2678));
 sg13g2_tiehi _27796__2679 (.L_HI(net2679));
 sg13g2_tiehi _27795__2680 (.L_HI(net2680));
 sg13g2_tiehi _27794__2681 (.L_HI(net2681));
 sg13g2_tiehi _27793__2682 (.L_HI(net2682));
 sg13g2_tiehi _27792__2683 (.L_HI(net2683));
 sg13g2_tiehi _27791__2684 (.L_HI(net2684));
 sg13g2_tiehi _27790__2685 (.L_HI(net2685));
 sg13g2_tiehi _27789__2686 (.L_HI(net2686));
 sg13g2_tiehi _27788__2687 (.L_HI(net2687));
 sg13g2_tiehi _27787__2688 (.L_HI(net2688));
 sg13g2_tiehi _27786__2689 (.L_HI(net2689));
 sg13g2_tiehi _27785__2690 (.L_HI(net2690));
 sg13g2_tiehi _27784__2691 (.L_HI(net2691));
 sg13g2_tiehi _27783__2692 (.L_HI(net2692));
 sg13g2_tiehi _27782__2693 (.L_HI(net2693));
 sg13g2_tiehi _27781__2694 (.L_HI(net2694));
 sg13g2_tiehi _27780__2695 (.L_HI(net2695));
 sg13g2_tiehi _27779__2696 (.L_HI(net2696));
 sg13g2_tiehi _27778__2697 (.L_HI(net2697));
 sg13g2_tiehi _27777__2698 (.L_HI(net2698));
 sg13g2_tiehi _27776__2699 (.L_HI(net2699));
 sg13g2_tiehi _30645__2700 (.L_HI(net2700));
 sg13g2_tiehi _30644__2701 (.L_HI(net2701));
 sg13g2_tiehi _30643__2702 (.L_HI(net2702));
 sg13g2_tiehi _30642__2703 (.L_HI(net2703));
 sg13g2_tiehi _30641__2704 (.L_HI(net2704));
 sg13g2_tiehi _30640__2705 (.L_HI(net2705));
 sg13g2_tiehi _30639__2706 (.L_HI(net2706));
 sg13g2_tiehi _30638__2707 (.L_HI(net2707));
 sg13g2_tiehi _30637__2708 (.L_HI(net2708));
 sg13g2_tiehi _30636__2709 (.L_HI(net2709));
 sg13g2_tiehi _30635__2710 (.L_HI(net2710));
 sg13g2_tiehi _30634__2711 (.L_HI(net2711));
 sg13g2_tiehi _30633__2712 (.L_HI(net2712));
 sg13g2_tiehi _30632__2713 (.L_HI(net2713));
 sg13g2_tiehi _30631__2714 (.L_HI(net2714));
 sg13g2_tiehi _30630__2715 (.L_HI(net2715));
 sg13g2_tiehi _30629__2716 (.L_HI(net2716));
 sg13g2_tiehi _30628__2717 (.L_HI(net2717));
 sg13g2_tiehi _30627__2718 (.L_HI(net2718));
 sg13g2_tiehi _30626__2719 (.L_HI(net2719));
 sg13g2_tiehi _30625__2720 (.L_HI(net2720));
 sg13g2_tiehi _30624__2721 (.L_HI(net2721));
 sg13g2_tiehi _30623__2722 (.L_HI(net2722));
 sg13g2_tiehi _30622__2723 (.L_HI(net2723));
 sg13g2_tiehi _30621__2724 (.L_HI(net2724));
 sg13g2_tiehi _30620__2725 (.L_HI(net2725));
 sg13g2_tiehi _30619__2726 (.L_HI(net2726));
 sg13g2_tiehi _30618__2727 (.L_HI(net2727));
 sg13g2_tiehi _30617__2728 (.L_HI(net2728));
 sg13g2_tiehi _30616__2729 (.L_HI(net2729));
 sg13g2_tiehi _30615__2730 (.L_HI(net2730));
 sg13g2_tiehi _30614__2731 (.L_HI(net2731));
 sg13g2_tiehi _30613__2732 (.L_HI(net2732));
 sg13g2_tiehi _30612__2733 (.L_HI(net2733));
 sg13g2_tiehi _30611__2734 (.L_HI(net2734));
 sg13g2_tiehi _30610__2735 (.L_HI(net2735));
 sg13g2_tiehi _30609__2736 (.L_HI(net2736));
 sg13g2_tiehi _30608__2737 (.L_HI(net2737));
 sg13g2_tiehi _30607__2738 (.L_HI(net2738));
 sg13g2_tiehi _30606__2739 (.L_HI(net2739));
 sg13g2_tiehi _30605__2740 (.L_HI(net2740));
 sg13g2_tiehi _30604__2741 (.L_HI(net2741));
 sg13g2_tiehi _30603__2742 (.L_HI(net2742));
 sg13g2_tiehi _30602__2743 (.L_HI(net2743));
 sg13g2_tiehi _30601__2744 (.L_HI(net2744));
 sg13g2_tiehi _30600__2745 (.L_HI(net2745));
 sg13g2_tiehi _30599__2746 (.L_HI(net2746));
 sg13g2_tiehi _30598__2747 (.L_HI(net2747));
 sg13g2_tiehi _30597__2748 (.L_HI(net2748));
 sg13g2_tiehi _30596__2749 (.L_HI(net2749));
 sg13g2_tiehi _30595__2750 (.L_HI(net2750));
 sg13g2_tiehi _30594__2751 (.L_HI(net2751));
 sg13g2_tiehi _30593__2752 (.L_HI(net2752));
 sg13g2_tiehi _30592__2753 (.L_HI(net2753));
 sg13g2_tiehi _30591__2754 (.L_HI(net2754));
 sg13g2_tiehi _30590__2755 (.L_HI(net2755));
 sg13g2_tiehi _30589__2756 (.L_HI(net2756));
 sg13g2_tiehi _30588__2757 (.L_HI(net2757));
 sg13g2_tiehi _30587__2758 (.L_HI(net2758));
 sg13g2_tiehi _30586__2759 (.L_HI(net2759));
 sg13g2_tiehi _30585__2760 (.L_HI(net2760));
 sg13g2_tiehi _30584__2761 (.L_HI(net2761));
 sg13g2_tiehi _30583__2762 (.L_HI(net2762));
 sg13g2_tiehi _30582__2763 (.L_HI(net2763));
 sg13g2_tiehi _30581__2764 (.L_HI(net2764));
 sg13g2_tiehi _30580__2765 (.L_HI(net2765));
 sg13g2_tiehi _30579__2766 (.L_HI(net2766));
 sg13g2_tiehi _30578__2767 (.L_HI(net2767));
 sg13g2_tiehi _30577__2768 (.L_HI(net2768));
 sg13g2_tiehi _30576__2769 (.L_HI(net2769));
 sg13g2_tiehi _30575__2770 (.L_HI(net2770));
 sg13g2_tiehi _30574__2771 (.L_HI(net2771));
 sg13g2_tiehi _30573__2772 (.L_HI(net2772));
 sg13g2_tiehi _30572__2773 (.L_HI(net2773));
 sg13g2_tiehi _30571__2774 (.L_HI(net2774));
 sg13g2_tiehi _30570__2775 (.L_HI(net2775));
 sg13g2_tiehi _30569__2776 (.L_HI(net2776));
 sg13g2_tiehi _30568__2777 (.L_HI(net2777));
 sg13g2_tiehi _30567__2778 (.L_HI(net2778));
 sg13g2_tiehi _30566__2779 (.L_HI(net2779));
 sg13g2_tiehi _30565__2780 (.L_HI(net2780));
 sg13g2_tiehi _30564__2781 (.L_HI(net2781));
 sg13g2_tiehi _30563__2782 (.L_HI(net2782));
 sg13g2_tiehi _30562__2783 (.L_HI(net2783));
 sg13g2_tiehi _30561__2784 (.L_HI(net2784));
 sg13g2_tiehi _30560__2785 (.L_HI(net2785));
 sg13g2_tiehi _30559__2786 (.L_HI(net2786));
 sg13g2_tiehi _30558__2787 (.L_HI(net2787));
 sg13g2_tiehi _30557__2788 (.L_HI(net2788));
 sg13g2_tiehi _30556__2789 (.L_HI(net2789));
 sg13g2_tiehi _30555__2790 (.L_HI(net2790));
 sg13g2_tiehi _30554__2791 (.L_HI(net2791));
 sg13g2_tiehi _30553__2792 (.L_HI(net2792));
 sg13g2_tiehi _30552__2793 (.L_HI(net2793));
 sg13g2_tiehi _30551__2794 (.L_HI(net2794));
 sg13g2_tiehi _30550__2795 (.L_HI(net2795));
 sg13g2_tiehi _30549__2796 (.L_HI(net2796));
 sg13g2_tiehi _30548__2797 (.L_HI(net2797));
 sg13g2_tiehi _30547__2798 (.L_HI(net2798));
 sg13g2_tiehi _30546__2799 (.L_HI(net2799));
 sg13g2_tiehi _30545__2800 (.L_HI(net2800));
 sg13g2_tiehi _30544__2801 (.L_HI(net2801));
 sg13g2_tiehi _30543__2802 (.L_HI(net2802));
 sg13g2_tiehi _30542__2803 (.L_HI(net2803));
 sg13g2_tiehi _30541__2804 (.L_HI(net2804));
 sg13g2_tiehi _30540__2805 (.L_HI(net2805));
 sg13g2_tiehi _30539__2806 (.L_HI(net2806));
 sg13g2_tiehi _30538__2807 (.L_HI(net2807));
 sg13g2_tiehi _30537__2808 (.L_HI(net2808));
 sg13g2_tiehi _30536__2809 (.L_HI(net2809));
 sg13g2_tiehi _30535__2810 (.L_HI(net2810));
 sg13g2_tiehi _30534__2811 (.L_HI(net2811));
 sg13g2_tiehi _30533__2812 (.L_HI(net2812));
 sg13g2_tiehi _30532__2813 (.L_HI(net2813));
 sg13g2_tiehi _30531__2814 (.L_HI(net2814));
 sg13g2_tiehi _30530__2815 (.L_HI(net2815));
 sg13g2_tiehi _30529__2816 (.L_HI(net2816));
 sg13g2_tiehi _30528__2817 (.L_HI(net2817));
 sg13g2_tiehi _30527__2818 (.L_HI(net2818));
 sg13g2_tiehi _30526__2819 (.L_HI(net2819));
 sg13g2_tiehi _30525__2820 (.L_HI(net2820));
 sg13g2_tiehi _30524__2821 (.L_HI(net2821));
 sg13g2_tiehi _30523__2822 (.L_HI(net2822));
 sg13g2_tiehi _30522__2823 (.L_HI(net2823));
 sg13g2_tiehi _30521__2824 (.L_HI(net2824));
 sg13g2_tiehi _30520__2825 (.L_HI(net2825));
 sg13g2_tiehi _30519__2826 (.L_HI(net2826));
 sg13g2_tiehi _30518__2827 (.L_HI(net2827));
 sg13g2_tiehi _30517__2828 (.L_HI(net2828));
 sg13g2_tiehi _30516__2829 (.L_HI(net2829));
 sg13g2_tiehi _30515__2830 (.L_HI(net2830));
 sg13g2_tiehi _30514__2831 (.L_HI(net2831));
 sg13g2_tiehi _30513__2832 (.L_HI(net2832));
 sg13g2_tiehi _30512__2833 (.L_HI(net2833));
 sg13g2_tiehi _30511__2834 (.L_HI(net2834));
 sg13g2_tiehi _30510__2835 (.L_HI(net2835));
 sg13g2_tiehi _30509__2836 (.L_HI(net2836));
 sg13g2_tiehi _30508__2837 (.L_HI(net2837));
 sg13g2_tiehi _30507__2838 (.L_HI(net2838));
 sg13g2_tiehi _30506__2839 (.L_HI(net2839));
 sg13g2_tiehi _30505__2840 (.L_HI(net2840));
 sg13g2_tiehi _30504__2841 (.L_HI(net2841));
 sg13g2_tiehi _30503__2842 (.L_HI(net2842));
 sg13g2_tiehi _30502__2843 (.L_HI(net2843));
 sg13g2_tiehi _30501__2844 (.L_HI(net2844));
 sg13g2_tiehi _30500__2845 (.L_HI(net2845));
 sg13g2_tiehi _30499__2846 (.L_HI(net2846));
 sg13g2_tiehi _30498__2847 (.L_HI(net2847));
 sg13g2_tiehi _30497__2848 (.L_HI(net2848));
 sg13g2_tiehi _30496__2849 (.L_HI(net2849));
 sg13g2_tiehi _30495__2850 (.L_HI(net2850));
 sg13g2_tiehi _30494__2851 (.L_HI(net2851));
 sg13g2_tiehi _30493__2852 (.L_HI(net2852));
 sg13g2_tiehi _30492__2853 (.L_HI(net2853));
 sg13g2_tiehi _30491__2854 (.L_HI(net2854));
 sg13g2_tiehi _30490__2855 (.L_HI(net2855));
 sg13g2_tiehi _30489__2856 (.L_HI(net2856));
 sg13g2_tiehi _30488__2857 (.L_HI(net2857));
 sg13g2_tiehi _30487__2858 (.L_HI(net2858));
 sg13g2_tiehi _30486__2859 (.L_HI(net2859));
 sg13g2_tiehi _30485__2860 (.L_HI(net2860));
 sg13g2_tiehi _30484__2861 (.L_HI(net2861));
 sg13g2_tiehi _30483__2862 (.L_HI(net2862));
 sg13g2_tiehi _30482__2863 (.L_HI(net2863));
 sg13g2_tiehi _30481__2864 (.L_HI(net2864));
 sg13g2_tiehi _30480__2865 (.L_HI(net2865));
 sg13g2_tiehi _30479__2866 (.L_HI(net2866));
 sg13g2_tiehi _30478__2867 (.L_HI(net2867));
 sg13g2_tiehi _30477__2868 (.L_HI(net2868));
 sg13g2_tiehi _30476__2869 (.L_HI(net2869));
 sg13g2_tiehi _30475__2870 (.L_HI(net2870));
 sg13g2_tiehi _30474__2871 (.L_HI(net2871));
 sg13g2_tiehi _30473__2872 (.L_HI(net2872));
 sg13g2_tiehi _30472__2873 (.L_HI(net2873));
 sg13g2_tiehi _30471__2874 (.L_HI(net2874));
 sg13g2_tiehi _30470__2875 (.L_HI(net2875));
 sg13g2_tiehi _30469__2876 (.L_HI(net2876));
 sg13g2_tiehi _30468__2877 (.L_HI(net2877));
 sg13g2_tiehi _30467__2878 (.L_HI(net2878));
 sg13g2_tiehi _30466__2879 (.L_HI(net2879));
 sg13g2_tiehi _30465__2880 (.L_HI(net2880));
 sg13g2_tiehi _30464__2881 (.L_HI(net2881));
 sg13g2_tiehi _30463__2882 (.L_HI(net2882));
 sg13g2_tiehi _30462__2883 (.L_HI(net2883));
 sg13g2_tiehi _30461__2884 (.L_HI(net2884));
 sg13g2_tiehi _30460__2885 (.L_HI(net2885));
 sg13g2_tiehi _30459__2886 (.L_HI(net2886));
 sg13g2_tiehi _30458__2887 (.L_HI(net2887));
 sg13g2_tiehi _30457__2888 (.L_HI(net2888));
 sg13g2_tiehi _30456__2889 (.L_HI(net2889));
 sg13g2_tiehi _30455__2890 (.L_HI(net2890));
 sg13g2_tiehi _30454__2891 (.L_HI(net2891));
 sg13g2_tiehi _30453__2892 (.L_HI(net2892));
 sg13g2_tiehi _30452__2893 (.L_HI(net2893));
 sg13g2_tiehi _30451__2894 (.L_HI(net2894));
 sg13g2_tiehi _30450__2895 (.L_HI(net2895));
 sg13g2_tiehi _30449__2896 (.L_HI(net2896));
 sg13g2_tiehi _30448__2897 (.L_HI(net2897));
 sg13g2_tiehi _30447__2898 (.L_HI(net2898));
 sg13g2_tiehi _30446__2899 (.L_HI(net2899));
 sg13g2_tiehi _30445__2900 (.L_HI(net2900));
 sg13g2_tiehi _30444__2901 (.L_HI(net2901));
 sg13g2_tiehi _30443__2902 (.L_HI(net2902));
 sg13g2_tiehi _30442__2903 (.L_HI(net2903));
 sg13g2_tiehi _30441__2904 (.L_HI(net2904));
 sg13g2_tiehi _30440__2905 (.L_HI(net2905));
 sg13g2_tiehi _30439__2906 (.L_HI(net2906));
 sg13g2_tiehi _30438__2907 (.L_HI(net2907));
 sg13g2_tiehi _30437__2908 (.L_HI(net2908));
 sg13g2_tiehi _30436__2909 (.L_HI(net2909));
 sg13g2_tiehi _30435__2910 (.L_HI(net2910));
 sg13g2_tiehi _30434__2911 (.L_HI(net2911));
 sg13g2_tiehi _30433__2912 (.L_HI(net2912));
 sg13g2_tiehi _30432__2913 (.L_HI(net2913));
 sg13g2_tiehi _30431__2914 (.L_HI(net2914));
 sg13g2_tiehi _30430__2915 (.L_HI(net2915));
 sg13g2_tiehi _30429__2916 (.L_HI(net2916));
 sg13g2_tiehi _30428__2917 (.L_HI(net2917));
 sg13g2_tiehi _30427__2918 (.L_HI(net2918));
 sg13g2_tiehi _30426__2919 (.L_HI(net2919));
 sg13g2_tiehi _30425__2920 (.L_HI(net2920));
 sg13g2_tiehi _30424__2921 (.L_HI(net2921));
 sg13g2_tiehi _30423__2922 (.L_HI(net2922));
 sg13g2_tiehi tt_um_rejunity_atari2600_2923 (.L_HI(net2923));
 sg13g2_tiehi tt_um_rejunity_atari2600_2924 (.L_HI(net2924));
 sg13g2_tiehi tt_um_rejunity_atari2600_2925 (.L_HI(net2925));
 sg13g2_tiehi tt_um_rejunity_atari2600_2926 (.L_HI(net2926));
 sg13g2_tiehi tt_um_rejunity_atari2600_2927 (.L_HI(net2927));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _33606_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _33607_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _33608_ (.A(\flash_rom.spi_select ),
    .X(uio_out[0]));
 sg13g2_buf_1 _33609_ (.A(\flash_rom.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_1 _33610_ (.A(audio_pwm),
    .X(uio_out[7]));
 sg13g2_buf_2 _33611_ (.A(\hvsync_gen.vga.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _33612_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout4961 (.A(_07225_),
    .X(net4961));
 sg13g2_buf_2 fanout4962 (.A(_07225_),
    .X(net4962));
 sg13g2_buf_2 fanout4963 (.A(_06457_),
    .X(net4963));
 sg13g2_buf_2 fanout4964 (.A(_06457_),
    .X(net4964));
 sg13g2_buf_2 fanout4965 (.A(_05996_),
    .X(net4965));
 sg13g2_buf_2 fanout4966 (.A(_05996_),
    .X(net4966));
 sg13g2_buf_4 fanout4967 (.X(net4967),
    .A(net4968));
 sg13g2_buf_2 fanout4968 (.A(_07224_),
    .X(net4968));
 sg13g2_buf_2 fanout4969 (.A(_07160_),
    .X(net4969));
 sg13g2_buf_1 fanout4970 (.A(_07160_),
    .X(net4970));
 sg13g2_buf_2 fanout4971 (.A(net4974),
    .X(net4971));
 sg13g2_buf_1 fanout4972 (.A(net4974),
    .X(net4972));
 sg13g2_buf_2 fanout4973 (.A(net4974),
    .X(net4973));
 sg13g2_buf_2 fanout4974 (.A(_07160_),
    .X(net4974));
 sg13g2_buf_2 fanout4975 (.A(_03208_),
    .X(net4975));
 sg13g2_buf_2 fanout4976 (.A(_03208_),
    .X(net4976));
 sg13g2_buf_2 fanout4977 (.A(net4981),
    .X(net4977));
 sg13g2_buf_1 fanout4978 (.A(net4981),
    .X(net4978));
 sg13g2_buf_2 fanout4979 (.A(net4981),
    .X(net4979));
 sg13g2_buf_2 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_1 fanout4981 (.A(_03207_),
    .X(net4981));
 sg13g2_buf_4 fanout4982 (.X(net4982),
    .A(_03205_));
 sg13g2_buf_2 fanout4983 (.A(_03205_),
    .X(net4983));
 sg13g2_buf_2 fanout4984 (.A(net4990),
    .X(net4984));
 sg13g2_buf_1 fanout4985 (.A(net4990),
    .X(net4985));
 sg13g2_buf_2 fanout4986 (.A(net4990),
    .X(net4986));
 sg13g2_buf_2 fanout4987 (.A(net4990),
    .X(net4987));
 sg13g2_buf_2 fanout4988 (.A(net4989),
    .X(net4988));
 sg13g2_buf_2 fanout4989 (.A(net4990),
    .X(net4989));
 sg13g2_buf_2 fanout4990 (.A(_03204_),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(_05381_),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(net4993),
    .X(net4992));
 sg13g2_buf_2 fanout4993 (.A(_08219_),
    .X(net4993));
 sg13g2_buf_2 fanout4994 (.A(net4995),
    .X(net4994));
 sg13g2_buf_2 fanout4995 (.A(_08186_),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(_08177_),
    .X(net4996));
 sg13g2_buf_2 fanout4997 (.A(_08177_),
    .X(net4997));
 sg13g2_buf_2 fanout4998 (.A(_08168_),
    .X(net4998));
 sg13g2_buf_2 fanout4999 (.A(_08168_),
    .X(net4999));
 sg13g2_buf_2 fanout5000 (.A(_08159_),
    .X(net5000));
 sg13g2_buf_2 fanout5001 (.A(_08159_),
    .X(net5001));
 sg13g2_buf_2 fanout5002 (.A(_08149_),
    .X(net5002));
 sg13g2_buf_2 fanout5003 (.A(_08149_),
    .X(net5003));
 sg13g2_buf_2 fanout5004 (.A(_08097_),
    .X(net5004));
 sg13g2_buf_2 fanout5005 (.A(_08097_),
    .X(net5005));
 sg13g2_buf_2 fanout5006 (.A(_08087_),
    .X(net5006));
 sg13g2_buf_2 fanout5007 (.A(_08087_),
    .X(net5007));
 sg13g2_buf_2 fanout5008 (.A(_08078_),
    .X(net5008));
 sg13g2_buf_2 fanout5009 (.A(_08078_),
    .X(net5009));
 sg13g2_buf_2 fanout5010 (.A(net5011),
    .X(net5010));
 sg13g2_buf_2 fanout5011 (.A(_08069_),
    .X(net5011));
 sg13g2_buf_2 fanout5012 (.A(net5013),
    .X(net5012));
 sg13g2_buf_2 fanout5013 (.A(_08060_),
    .X(net5013));
 sg13g2_buf_2 fanout5014 (.A(_08051_),
    .X(net5014));
 sg13g2_buf_2 fanout5015 (.A(_08051_),
    .X(net5015));
 sg13g2_buf_2 fanout5016 (.A(_08033_),
    .X(net5016));
 sg13g2_buf_2 fanout5017 (.A(_08033_),
    .X(net5017));
 sg13g2_buf_2 fanout5018 (.A(_07959_),
    .X(net5018));
 sg13g2_buf_2 fanout5019 (.A(_07959_),
    .X(net5019));
 sg13g2_buf_2 fanout5020 (.A(net5021),
    .X(net5020));
 sg13g2_buf_2 fanout5021 (.A(_07911_),
    .X(net5021));
 sg13g2_buf_2 fanout5022 (.A(net5023),
    .X(net5022));
 sg13g2_buf_2 fanout5023 (.A(_07898_),
    .X(net5023));
 sg13g2_buf_2 fanout5024 (.A(_07889_),
    .X(net5024));
 sg13g2_buf_2 fanout5025 (.A(_07889_),
    .X(net5025));
 sg13g2_buf_2 fanout5026 (.A(net5027),
    .X(net5026));
 sg13g2_buf_2 fanout5027 (.A(_07880_),
    .X(net5027));
 sg13g2_buf_2 fanout5028 (.A(net5029),
    .X(net5028));
 sg13g2_buf_2 fanout5029 (.A(_07844_),
    .X(net5029));
 sg13g2_buf_2 fanout5030 (.A(net5031),
    .X(net5030));
 sg13g2_buf_2 fanout5031 (.A(_07816_),
    .X(net5031));
 sg13g2_buf_2 fanout5032 (.A(net5034),
    .X(net5032));
 sg13g2_buf_1 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_2 fanout5034 (.A(_07807_),
    .X(net5034));
 sg13g2_buf_2 fanout5035 (.A(_07791_),
    .X(net5035));
 sg13g2_buf_2 fanout5036 (.A(_07791_),
    .X(net5036));
 sg13g2_buf_2 fanout5037 (.A(net5038),
    .X(net5037));
 sg13g2_buf_2 fanout5038 (.A(_07782_),
    .X(net5038));
 sg13g2_buf_2 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_2 fanout5040 (.A(_07362_),
    .X(net5040));
 sg13g2_buf_2 fanout5041 (.A(net5042),
    .X(net5041));
 sg13g2_buf_2 fanout5042 (.A(_07353_),
    .X(net5042));
 sg13g2_buf_2 fanout5043 (.A(net5044),
    .X(net5043));
 sg13g2_buf_2 fanout5044 (.A(_07323_),
    .X(net5044));
 sg13g2_buf_2 fanout5045 (.A(_07311_),
    .X(net5045));
 sg13g2_buf_2 fanout5046 (.A(_07311_),
    .X(net5046));
 sg13g2_buf_2 fanout5047 (.A(_07293_),
    .X(net5047));
 sg13g2_buf_2 fanout5048 (.A(_07293_),
    .X(net5048));
 sg13g2_buf_2 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_2 fanout5050 (.A(_07013_),
    .X(net5050));
 sg13g2_buf_2 fanout5051 (.A(net5052),
    .X(net5051));
 sg13g2_buf_4 fanout5052 (.X(net5052),
    .A(_06946_));
 sg13g2_buf_2 fanout5053 (.A(_06874_),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(net5055),
    .X(net5054));
 sg13g2_buf_4 fanout5055 (.X(net5055),
    .A(_06824_));
 sg13g2_buf_2 fanout5056 (.A(_06756_),
    .X(net5056));
 sg13g2_buf_1 fanout5057 (.A(_06756_),
    .X(net5057));
 sg13g2_buf_2 fanout5058 (.A(net5059),
    .X(net5058));
 sg13g2_buf_2 fanout5059 (.A(_05604_),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net5062),
    .X(net5060));
 sg13g2_buf_1 fanout5061 (.A(net5062),
    .X(net5061));
 sg13g2_buf_2 fanout5062 (.A(_05173_),
    .X(net5062));
 sg13g2_buf_2 fanout5063 (.A(net5064),
    .X(net5063));
 sg13g2_buf_2 fanout5064 (.A(_04985_),
    .X(net5064));
 sg13g2_buf_2 fanout5065 (.A(_04909_),
    .X(net5065));
 sg13g2_buf_2 fanout5066 (.A(_04909_),
    .X(net5066));
 sg13g2_buf_2 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_2 fanout5068 (.A(_04871_),
    .X(net5068));
 sg13g2_buf_2 fanout5069 (.A(net5070),
    .X(net5069));
 sg13g2_buf_2 fanout5070 (.A(_04838_),
    .X(net5070));
 sg13g2_buf_2 fanout5071 (.A(net5072),
    .X(net5071));
 sg13g2_buf_2 fanout5072 (.A(_03144_),
    .X(net5072));
 sg13g2_buf_2 fanout5073 (.A(net5075),
    .X(net5073));
 sg13g2_buf_1 fanout5074 (.A(net5075),
    .X(net5074));
 sg13g2_buf_2 fanout5075 (.A(_03135_),
    .X(net5075));
 sg13g2_buf_2 fanout5076 (.A(_03070_),
    .X(net5076));
 sg13g2_buf_2 fanout5077 (.A(_03070_),
    .X(net5077));
 sg13g2_buf_2 fanout5078 (.A(_10066_),
    .X(net5078));
 sg13g2_buf_4 fanout5079 (.X(net5079),
    .A(_09205_));
 sg13g2_buf_4 fanout5080 (.X(net5080),
    .A(_09174_));
 sg13g2_buf_2 fanout5081 (.A(net5082),
    .X(net5081));
 sg13g2_buf_2 fanout5082 (.A(_08042_),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(_08024_),
    .X(net5083));
 sg13g2_buf_2 fanout5084 (.A(_08024_),
    .X(net5084));
 sg13g2_buf_2 fanout5085 (.A(net5086),
    .X(net5085));
 sg13g2_buf_2 fanout5086 (.A(_08014_),
    .X(net5086));
 sg13g2_buf_2 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(_08005_),
    .X(net5088));
 sg13g2_buf_2 fanout5089 (.A(net5090),
    .X(net5089));
 sg13g2_buf_2 fanout5090 (.A(_07996_),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(_07986_),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(_07986_),
    .X(net5092));
 sg13g2_buf_2 fanout5093 (.A(net5094),
    .X(net5093));
 sg13g2_buf_2 fanout5094 (.A(_07977_),
    .X(net5094));
 sg13g2_buf_2 fanout5095 (.A(_07968_),
    .X(net5095));
 sg13g2_buf_2 fanout5096 (.A(_07968_),
    .X(net5096));
 sg13g2_buf_2 fanout5097 (.A(net5098),
    .X(net5097));
 sg13g2_buf_2 fanout5098 (.A(_07950_),
    .X(net5098));
 sg13g2_buf_2 fanout5099 (.A(net5100),
    .X(net5099));
 sg13g2_buf_2 fanout5100 (.A(_07941_),
    .X(net5100));
 sg13g2_buf_2 fanout5101 (.A(net5102),
    .X(net5101));
 sg13g2_buf_2 fanout5102 (.A(_07932_),
    .X(net5102));
 sg13g2_buf_2 fanout5103 (.A(net5104),
    .X(net5103));
 sg13g2_buf_2 fanout5104 (.A(_07835_),
    .X(net5104));
 sg13g2_buf_2 fanout5105 (.A(_07340_),
    .X(net5105));
 sg13g2_buf_2 fanout5106 (.A(_07340_),
    .X(net5106));
 sg13g2_buf_2 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_2 fanout5108 (.A(_07266_),
    .X(net5108));
 sg13g2_buf_2 fanout5109 (.A(net5110),
    .X(net5109));
 sg13g2_buf_2 fanout5110 (.A(_07251_),
    .X(net5110));
 sg13g2_buf_2 fanout5111 (.A(_07136_),
    .X(net5111));
 sg13g2_buf_2 fanout5112 (.A(net5113),
    .X(net5112));
 sg13g2_buf_2 fanout5113 (.A(_07059_),
    .X(net5113));
 sg13g2_buf_2 fanout5114 (.A(net5116),
    .X(net5114));
 sg13g2_buf_2 fanout5115 (.A(net5116),
    .X(net5115));
 sg13g2_buf_2 fanout5116 (.A(_06618_),
    .X(net5116));
 sg13g2_buf_2 fanout5117 (.A(_06581_),
    .X(net5117));
 sg13g2_buf_2 fanout5118 (.A(_06581_),
    .X(net5118));
 sg13g2_buf_2 fanout5119 (.A(_06573_),
    .X(net5119));
 sg13g2_buf_2 fanout5120 (.A(_06573_),
    .X(net5120));
 sg13g2_buf_2 fanout5121 (.A(_06564_),
    .X(net5121));
 sg13g2_buf_2 fanout5122 (.A(_06564_),
    .X(net5122));
 sg13g2_buf_2 fanout5123 (.A(_06556_),
    .X(net5123));
 sg13g2_buf_2 fanout5124 (.A(_06556_),
    .X(net5124));
 sg13g2_buf_2 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_2 fanout5126 (.A(_05539_),
    .X(net5126));
 sg13g2_buf_2 fanout5127 (.A(net5128),
    .X(net5127));
 sg13g2_buf_2 fanout5128 (.A(_05507_),
    .X(net5128));
 sg13g2_buf_2 fanout5129 (.A(net5130),
    .X(net5129));
 sg13g2_buf_2 fanout5130 (.A(_05494_),
    .X(net5130));
 sg13g2_buf_2 fanout5131 (.A(net5132),
    .X(net5131));
 sg13g2_buf_2 fanout5132 (.A(_05467_),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(_05466_),
    .X(net5133));
 sg13g2_buf_2 fanout5134 (.A(_05376_),
    .X(net5134));
 sg13g2_buf_2 fanout5135 (.A(net5136),
    .X(net5135));
 sg13g2_buf_2 fanout5136 (.A(_05223_),
    .X(net5136));
 sg13g2_buf_2 fanout5137 (.A(net5138),
    .X(net5137));
 sg13g2_buf_2 fanout5138 (.A(_05203_),
    .X(net5138));
 sg13g2_buf_2 fanout5139 (.A(net5140),
    .X(net5139));
 sg13g2_buf_2 fanout5140 (.A(_05193_),
    .X(net5140));
 sg13g2_buf_2 fanout5141 (.A(_05183_),
    .X(net5141));
 sg13g2_buf_2 fanout5142 (.A(_05183_),
    .X(net5142));
 sg13g2_buf_2 fanout5143 (.A(_05117_),
    .X(net5143));
 sg13g2_buf_2 fanout5144 (.A(_05117_),
    .X(net5144));
 sg13g2_buf_2 fanout5145 (.A(_05108_),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(_05108_),
    .X(net5146));
 sg13g2_buf_2 fanout5147 (.A(_05099_),
    .X(net5147));
 sg13g2_buf_2 fanout5148 (.A(_05099_),
    .X(net5148));
 sg13g2_buf_2 fanout5149 (.A(_05090_),
    .X(net5149));
 sg13g2_buf_2 fanout5150 (.A(_05090_),
    .X(net5150));
 sg13g2_buf_2 fanout5151 (.A(_05080_),
    .X(net5151));
 sg13g2_buf_2 fanout5152 (.A(_05080_),
    .X(net5152));
 sg13g2_buf_2 fanout5153 (.A(_05071_),
    .X(net5153));
 sg13g2_buf_2 fanout5154 (.A(_05071_),
    .X(net5154));
 sg13g2_buf_2 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_2 fanout5156 (.A(_05062_),
    .X(net5156));
 sg13g2_buf_2 fanout5157 (.A(_05034_),
    .X(net5157));
 sg13g2_buf_2 fanout5158 (.A(_05034_),
    .X(net5158));
 sg13g2_buf_2 fanout5159 (.A(_05015_),
    .X(net5159));
 sg13g2_buf_2 fanout5160 (.A(_05015_),
    .X(net5160));
 sg13g2_buf_2 fanout5161 (.A(_04976_),
    .X(net5161));
 sg13g2_buf_2 fanout5162 (.A(_04976_),
    .X(net5162));
 sg13g2_buf_2 fanout5163 (.A(_04957_),
    .X(net5163));
 sg13g2_buf_2 fanout5164 (.A(_04957_),
    .X(net5164));
 sg13g2_buf_2 fanout5165 (.A(_04936_),
    .X(net5165));
 sg13g2_buf_2 fanout5166 (.A(_04936_),
    .X(net5166));
 sg13g2_buf_2 fanout5167 (.A(_04927_),
    .X(net5167));
 sg13g2_buf_2 fanout5168 (.A(_04927_),
    .X(net5168));
 sg13g2_buf_2 fanout5169 (.A(net5170),
    .X(net5169));
 sg13g2_buf_2 fanout5170 (.A(_04918_),
    .X(net5170));
 sg13g2_buf_2 fanout5171 (.A(_04900_),
    .X(net5171));
 sg13g2_buf_2 fanout5172 (.A(_04900_),
    .X(net5172));
 sg13g2_buf_2 fanout5173 (.A(_04891_),
    .X(net5173));
 sg13g2_buf_2 fanout5174 (.A(_04891_),
    .X(net5174));
 sg13g2_buf_2 fanout5175 (.A(net5176),
    .X(net5175));
 sg13g2_buf_2 fanout5176 (.A(_04882_),
    .X(net5176));
 sg13g2_buf_2 fanout5177 (.A(net5178),
    .X(net5177));
 sg13g2_buf_2 fanout5178 (.A(_04847_),
    .X(net5178));
 sg13g2_buf_2 fanout5179 (.A(net5180),
    .X(net5179));
 sg13g2_buf_2 fanout5180 (.A(_04829_),
    .X(net5180));
 sg13g2_buf_2 fanout5181 (.A(_04820_),
    .X(net5181));
 sg13g2_buf_2 fanout5182 (.A(_04820_),
    .X(net5182));
 sg13g2_buf_2 fanout5183 (.A(net5184),
    .X(net5183));
 sg13g2_buf_2 fanout5184 (.A(_04811_),
    .X(net5184));
 sg13g2_buf_2 fanout5185 (.A(_04802_),
    .X(net5185));
 sg13g2_buf_2 fanout5186 (.A(_04802_),
    .X(net5186));
 sg13g2_buf_2 fanout5187 (.A(net5188),
    .X(net5187));
 sg13g2_buf_2 fanout5188 (.A(_04793_),
    .X(net5188));
 sg13g2_buf_2 fanout5189 (.A(_04783_),
    .X(net5189));
 sg13g2_buf_2 fanout5190 (.A(_04783_),
    .X(net5190));
 sg13g2_buf_2 fanout5191 (.A(net5192),
    .X(net5191));
 sg13g2_buf_2 fanout5192 (.A(_04768_),
    .X(net5192));
 sg13g2_buf_2 fanout5193 (.A(_03113_),
    .X(net5193));
 sg13g2_buf_2 fanout5194 (.A(_03113_),
    .X(net5194));
 sg13g2_buf_2 fanout5195 (.A(_03104_),
    .X(net5195));
 sg13g2_buf_2 fanout5196 (.A(_03104_),
    .X(net5196));
 sg13g2_buf_2 fanout5197 (.A(net5198),
    .X(net5197));
 sg13g2_buf_2 fanout5198 (.A(_03094_),
    .X(net5198));
 sg13g2_buf_2 fanout5199 (.A(_03082_),
    .X(net5199));
 sg13g2_buf_2 fanout5200 (.A(_03082_),
    .X(net5200));
 sg13g2_buf_2 fanout5201 (.A(net5202),
    .X(net5201));
 sg13g2_buf_2 fanout5202 (.A(_03028_),
    .X(net5202));
 sg13g2_buf_4 fanout5203 (.X(net5203),
    .A(_09414_));
 sg13g2_buf_2 fanout5204 (.A(net5205),
    .X(net5204));
 sg13g2_buf_2 fanout5205 (.A(_07922_),
    .X(net5205));
 sg13g2_buf_2 fanout5206 (.A(_07302_),
    .X(net5206));
 sg13g2_buf_2 fanout5207 (.A(_07302_),
    .X(net5207));
 sg13g2_buf_2 fanout5208 (.A(_07284_),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(_07284_),
    .X(net5209));
 sg13g2_buf_2 fanout5210 (.A(_07275_),
    .X(net5210));
 sg13g2_buf_2 fanout5211 (.A(_07275_),
    .X(net5211));
 sg13g2_buf_4 fanout5212 (.X(net5212),
    .A(_07145_));
 sg13g2_buf_4 fanout5213 (.X(net5213),
    .A(_06944_));
 sg13g2_buf_2 fanout5214 (.A(_06871_),
    .X(net5214));
 sg13g2_buf_2 fanout5215 (.A(_05579_),
    .X(net5215));
 sg13g2_buf_2 fanout5216 (.A(_05579_),
    .X(net5216));
 sg13g2_buf_4 fanout5217 (.X(net5217),
    .A(_05504_));
 sg13g2_buf_2 fanout5218 (.A(_05503_),
    .X(net5218));
 sg13g2_buf_2 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_2 fanout5220 (.A(_05213_),
    .X(net5220));
 sg13g2_buf_2 fanout5221 (.A(net5223),
    .X(net5221));
 sg13g2_buf_1 fanout5222 (.A(net5223),
    .X(net5222));
 sg13g2_buf_2 fanout5223 (.A(_05052_),
    .X(net5223));
 sg13g2_buf_2 fanout5224 (.A(_05043_),
    .X(net5224));
 sg13g2_buf_2 fanout5225 (.A(_05043_),
    .X(net5225));
 sg13g2_buf_2 fanout5226 (.A(_05024_),
    .X(net5226));
 sg13g2_buf_2 fanout5227 (.A(_05024_),
    .X(net5227));
 sg13g2_buf_2 fanout5228 (.A(_05006_),
    .X(net5228));
 sg13g2_buf_2 fanout5229 (.A(_05006_),
    .X(net5229));
 sg13g2_buf_2 fanout5230 (.A(_04994_),
    .X(net5230));
 sg13g2_buf_2 fanout5231 (.A(_04994_),
    .X(net5231));
 sg13g2_buf_2 fanout5232 (.A(_04966_),
    .X(net5232));
 sg13g2_buf_2 fanout5233 (.A(_04966_),
    .X(net5233));
 sg13g2_buf_2 fanout5234 (.A(_04948_),
    .X(net5234));
 sg13g2_buf_2 fanout5235 (.A(_04948_),
    .X(net5235));
 sg13g2_buf_8 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(_04767_),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(_03093_),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(_03093_),
    .X(net5239));
 sg13g2_buf_2 fanout5240 (.A(net5245),
    .X(net5240));
 sg13g2_buf_2 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_2 fanout5242 (.A(net5245),
    .X(net5242));
 sg13g2_buf_2 fanout5243 (.A(net5244),
    .X(net5243));
 sg13g2_buf_2 fanout5244 (.A(net5245),
    .X(net5244));
 sg13g2_buf_2 fanout5245 (.A(_09364_),
    .X(net5245));
 sg13g2_buf_4 fanout5246 (.X(net5246),
    .A(_09128_));
 sg13g2_buf_2 fanout5247 (.A(_05367_),
    .X(net5247));
 sg13g2_buf_8 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(_04792_),
    .X(net5249));
 sg13g2_buf_4 fanout5250 (.X(net5250),
    .A(_04781_));
 sg13g2_buf_8 fanout5251 (.A(_04781_),
    .X(net5251));
 sg13g2_buf_8 fanout5252 (.A(net5253),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(_03125_),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5255),
    .X(net5254));
 sg13g2_buf_8 fanout5255 (.A(_03103_),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(net5257),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(_03081_),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(net5259),
    .X(net5258));
 sg13g2_buf_8 fanout5259 (.A(_03027_),
    .X(net5259));
 sg13g2_buf_2 fanout5260 (.A(net5262),
    .X(net5260));
 sg13g2_buf_1 fanout5261 (.A(net5262),
    .X(net5261));
 sg13g2_buf_2 fanout5262 (.A(_09641_),
    .X(net5262));
 sg13g2_buf_4 fanout5263 (.X(net5263),
    .A(_09436_));
 sg13g2_buf_2 fanout5264 (.A(net5265),
    .X(net5264));
 sg13g2_buf_2 fanout5265 (.A(net5267),
    .X(net5265));
 sg13g2_buf_2 fanout5266 (.A(net5267),
    .X(net5266));
 sg13g2_buf_4 fanout5267 (.X(net5267),
    .A(_09320_));
 sg13g2_buf_4 fanout5268 (.X(net5268),
    .A(_09302_));
 sg13g2_buf_4 fanout5269 (.X(net5269),
    .A(_09302_));
 sg13g2_buf_2 fanout5270 (.A(net5272),
    .X(net5270));
 sg13g2_buf_4 fanout5271 (.X(net5271),
    .A(net5272));
 sg13g2_buf_4 fanout5272 (.X(net5272),
    .A(_09106_));
 sg13g2_buf_2 fanout5273 (.A(_05364_),
    .X(net5273));
 sg13g2_buf_2 fanout5274 (.A(_05364_),
    .X(net5274));
 sg13g2_buf_8 fanout5275 (.A(net5278),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5278),
    .X(net5276));
 sg13g2_buf_1 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_4 fanout5278 (.X(net5278),
    .A(_09094_));
 sg13g2_buf_4 fanout5279 (.X(net5279),
    .A(net5280));
 sg13g2_buf_8 fanout5280 (.A(_09093_),
    .X(net5280));
 sg13g2_buf_8 fanout5281 (.A(net5283),
    .X(net5281));
 sg13g2_buf_2 fanout5282 (.A(net5283),
    .X(net5282));
 sg13g2_buf_4 fanout5283 (.X(net5283),
    .A(_09093_));
 sg13g2_buf_2 fanout5284 (.A(net5286),
    .X(net5284));
 sg13g2_buf_2 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_4 fanout5286 (.X(net5286),
    .A(_09936_));
 sg13g2_buf_2 fanout5287 (.A(net5289),
    .X(net5287));
 sg13g2_buf_2 fanout5288 (.A(net5289),
    .X(net5288));
 sg13g2_buf_2 fanout5289 (.A(_09877_),
    .X(net5289));
 sg13g2_buf_2 fanout5290 (.A(net5292),
    .X(net5290));
 sg13g2_buf_1 fanout5291 (.A(net5292),
    .X(net5291));
 sg13g2_buf_4 fanout5292 (.X(net5292),
    .A(_09814_));
 sg13g2_buf_4 fanout5293 (.X(net5293),
    .A(net5294));
 sg13g2_buf_4 fanout5294 (.X(net5294),
    .A(net5295));
 sg13g2_buf_4 fanout5295 (.X(net5295),
    .A(net5305));
 sg13g2_buf_4 fanout5296 (.X(net5296),
    .A(net5297));
 sg13g2_buf_4 fanout5297 (.X(net5297),
    .A(net5305));
 sg13g2_buf_4 fanout5298 (.X(net5298),
    .A(net5302));
 sg13g2_buf_2 fanout5299 (.A(net5302),
    .X(net5299));
 sg13g2_buf_4 fanout5300 (.X(net5300),
    .A(net5302));
 sg13g2_buf_2 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_2 fanout5302 (.A(net5305),
    .X(net5302));
 sg13g2_buf_4 fanout5303 (.X(net5303),
    .A(net5305));
 sg13g2_buf_2 fanout5304 (.A(net5305),
    .X(net5304));
 sg13g2_buf_4 fanout5305 (.X(net5305),
    .A(_09304_));
 sg13g2_buf_4 fanout5306 (.X(net5306),
    .A(net5308));
 sg13g2_buf_4 fanout5307 (.X(net5307),
    .A(net5308));
 sg13g2_buf_4 fanout5308 (.X(net5308),
    .A(net5311));
 sg13g2_buf_4 fanout5309 (.X(net5309),
    .A(net5310));
 sg13g2_buf_4 fanout5310 (.X(net5310),
    .A(net5311));
 sg13g2_buf_2 fanout5311 (.A(_09304_),
    .X(net5311));
 sg13g2_buf_4 fanout5312 (.X(net5312),
    .A(net5315));
 sg13g2_buf_2 fanout5313 (.A(net5315),
    .X(net5313));
 sg13g2_buf_4 fanout5314 (.X(net5314),
    .A(net5315));
 sg13g2_buf_2 fanout5315 (.A(net5318),
    .X(net5315));
 sg13g2_buf_4 fanout5316 (.X(net5316),
    .A(net5318));
 sg13g2_buf_4 fanout5317 (.X(net5317),
    .A(net5318));
 sg13g2_buf_2 fanout5318 (.A(net5337),
    .X(net5318));
 sg13g2_buf_4 fanout5319 (.X(net5319),
    .A(net5321));
 sg13g2_buf_4 fanout5320 (.X(net5320),
    .A(net5321));
 sg13g2_buf_2 fanout5321 (.A(net5337),
    .X(net5321));
 sg13g2_buf_4 fanout5322 (.X(net5322),
    .A(net5325));
 sg13g2_buf_4 fanout5323 (.X(net5323),
    .A(net5325));
 sg13g2_buf_2 fanout5324 (.A(net5325),
    .X(net5324));
 sg13g2_buf_2 fanout5325 (.A(net5337),
    .X(net5325));
 sg13g2_buf_4 fanout5326 (.X(net5326),
    .A(net5327));
 sg13g2_buf_4 fanout5327 (.X(net5327),
    .A(net5336));
 sg13g2_buf_4 fanout5328 (.X(net5328),
    .A(net5330));
 sg13g2_buf_4 fanout5329 (.X(net5329),
    .A(net5330));
 sg13g2_buf_4 fanout5330 (.X(net5330),
    .A(net5336));
 sg13g2_buf_4 fanout5331 (.X(net5331),
    .A(net5332));
 sg13g2_buf_4 fanout5332 (.X(net5332),
    .A(net5336));
 sg13g2_buf_4 fanout5333 (.X(net5333),
    .A(net5335));
 sg13g2_buf_2 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_4 fanout5335 (.X(net5335),
    .A(net5336));
 sg13g2_buf_4 fanout5336 (.X(net5336),
    .A(net5337));
 sg13g2_buf_4 fanout5337 (.X(net5337),
    .A(_09304_));
 sg13g2_buf_4 fanout5338 (.X(net5338),
    .A(_09299_));
 sg13g2_buf_4 fanout5339 (.X(net5339),
    .A(_09299_));
 sg13g2_buf_4 fanout5340 (.X(net5340),
    .A(net5341));
 sg13g2_buf_4 fanout5341 (.X(net5341),
    .A(net5343));
 sg13g2_buf_4 fanout5342 (.X(net5342),
    .A(net5343));
 sg13g2_buf_2 fanout5343 (.A(net5352),
    .X(net5343));
 sg13g2_buf_4 fanout5344 (.X(net5344),
    .A(net5352));
 sg13g2_buf_2 fanout5345 (.A(net5352),
    .X(net5345));
 sg13g2_buf_4 fanout5346 (.X(net5346),
    .A(net5348));
 sg13g2_buf_4 fanout5347 (.X(net5347),
    .A(net5348));
 sg13g2_buf_2 fanout5348 (.A(net5352),
    .X(net5348));
 sg13g2_buf_4 fanout5349 (.X(net5349),
    .A(net5351));
 sg13g2_buf_4 fanout5350 (.X(net5350),
    .A(net5351));
 sg13g2_buf_2 fanout5351 (.A(net5352),
    .X(net5351));
 sg13g2_buf_4 fanout5352 (.X(net5352),
    .A(_09298_));
 sg13g2_buf_4 fanout5353 (.X(net5353),
    .A(net5354));
 sg13g2_buf_4 fanout5354 (.X(net5354),
    .A(net5355));
 sg13g2_buf_4 fanout5355 (.X(net5355),
    .A(net5358));
 sg13g2_buf_4 fanout5356 (.X(net5356),
    .A(net5357));
 sg13g2_buf_4 fanout5357 (.X(net5357),
    .A(net5358));
 sg13g2_buf_2 fanout5358 (.A(_09298_),
    .X(net5358));
 sg13g2_buf_4 fanout5359 (.X(net5359),
    .A(net5361));
 sg13g2_buf_4 fanout5360 (.X(net5360),
    .A(net5364));
 sg13g2_buf_2 fanout5361 (.A(net5364),
    .X(net5361));
 sg13g2_buf_4 fanout5362 (.X(net5362),
    .A(net5363));
 sg13g2_buf_4 fanout5363 (.X(net5363),
    .A(net5364));
 sg13g2_buf_4 fanout5364 (.X(net5364),
    .A(net5383));
 sg13g2_buf_4 fanout5365 (.X(net5365),
    .A(net5367));
 sg13g2_buf_2 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_4 fanout5367 (.X(net5367),
    .A(net5370));
 sg13g2_buf_4 fanout5368 (.X(net5368),
    .A(net5369));
 sg13g2_buf_4 fanout5369 (.X(net5369),
    .A(net5370));
 sg13g2_buf_4 fanout5370 (.X(net5370),
    .A(net5383));
 sg13g2_buf_4 fanout5371 (.X(net5371),
    .A(net5372));
 sg13g2_buf_4 fanout5372 (.X(net5372),
    .A(net5376));
 sg13g2_buf_4 fanout5373 (.X(net5373),
    .A(net5374));
 sg13g2_buf_4 fanout5374 (.X(net5374),
    .A(net5376));
 sg13g2_buf_2 fanout5375 (.A(net5376),
    .X(net5375));
 sg13g2_buf_2 fanout5376 (.A(net5383),
    .X(net5376));
 sg13g2_buf_4 fanout5377 (.X(net5377),
    .A(net5379));
 sg13g2_buf_4 fanout5378 (.X(net5378),
    .A(net5379));
 sg13g2_buf_2 fanout5379 (.A(net5382),
    .X(net5379));
 sg13g2_buf_4 fanout5380 (.X(net5380),
    .A(net5381));
 sg13g2_buf_4 fanout5381 (.X(net5381),
    .A(net5382));
 sg13g2_buf_2 fanout5382 (.A(net5383),
    .X(net5382));
 sg13g2_buf_4 fanout5383 (.X(net5383),
    .A(_09298_));
 sg13g2_buf_8 fanout5384 (.A(_09210_),
    .X(net5384));
 sg13g2_buf_4 fanout5385 (.X(net5385),
    .A(net5388));
 sg13g2_buf_2 fanout5386 (.A(net5388),
    .X(net5386));
 sg13g2_buf_4 fanout5387 (.X(net5387),
    .A(net5388));
 sg13g2_buf_2 fanout5388 (.A(net5397),
    .X(net5388));
 sg13g2_buf_4 fanout5389 (.X(net5389),
    .A(net5397));
 sg13g2_buf_2 fanout5390 (.A(net5397),
    .X(net5390));
 sg13g2_buf_4 fanout5391 (.X(net5391),
    .A(net5393));
 sg13g2_buf_4 fanout5392 (.X(net5392),
    .A(net5393));
 sg13g2_buf_2 fanout5393 (.A(net5397),
    .X(net5393));
 sg13g2_buf_4 fanout5394 (.X(net5394),
    .A(net5396));
 sg13g2_buf_4 fanout5395 (.X(net5395),
    .A(net5396));
 sg13g2_buf_2 fanout5396 (.A(net5397),
    .X(net5396));
 sg13g2_buf_2 fanout5397 (.A(net5431),
    .X(net5397));
 sg13g2_buf_4 fanout5398 (.X(net5398),
    .A(net5400));
 sg13g2_buf_4 fanout5399 (.X(net5399),
    .A(net5400));
 sg13g2_buf_2 fanout5400 (.A(net5401),
    .X(net5400));
 sg13g2_buf_2 fanout5401 (.A(net5431),
    .X(net5401));
 sg13g2_buf_4 fanout5402 (.X(net5402),
    .A(net5404));
 sg13g2_buf_1 fanout5403 (.A(net5404),
    .X(net5403));
 sg13g2_buf_4 fanout5404 (.X(net5404),
    .A(net5405));
 sg13g2_buf_2 fanout5405 (.A(net5431),
    .X(net5405));
 sg13g2_buf_4 fanout5406 (.X(net5406),
    .A(net5411));
 sg13g2_buf_2 fanout5407 (.A(net5411),
    .X(net5407));
 sg13g2_buf_4 fanout5408 (.X(net5408),
    .A(net5410));
 sg13g2_buf_4 fanout5409 (.X(net5409),
    .A(net5410));
 sg13g2_buf_2 fanout5410 (.A(net5411),
    .X(net5410));
 sg13g2_buf_2 fanout5411 (.A(net5431),
    .X(net5411));
 sg13g2_buf_2 fanout5412 (.A(net5414),
    .X(net5412));
 sg13g2_buf_2 fanout5413 (.A(net5414),
    .X(net5413));
 sg13g2_buf_2 fanout5414 (.A(net5418),
    .X(net5414));
 sg13g2_buf_2 fanout5415 (.A(net5417),
    .X(net5415));
 sg13g2_buf_4 fanout5416 (.X(net5416),
    .A(net5418));
 sg13g2_buf_2 fanout5417 (.A(net5418),
    .X(net5417));
 sg13g2_buf_2 fanout5418 (.A(net5431),
    .X(net5418));
 sg13g2_buf_2 fanout5419 (.A(net5420),
    .X(net5419));
 sg13g2_buf_4 fanout5420 (.X(net5420),
    .A(net5424));
 sg13g2_buf_2 fanout5421 (.A(net5423),
    .X(net5421));
 sg13g2_buf_2 fanout5422 (.A(net5423),
    .X(net5422));
 sg13g2_buf_2 fanout5423 (.A(net5424),
    .X(net5423));
 sg13g2_buf_2 fanout5424 (.A(net5430),
    .X(net5424));
 sg13g2_buf_4 fanout5425 (.X(net5425),
    .A(net5427));
 sg13g2_buf_4 fanout5426 (.X(net5426),
    .A(net5427));
 sg13g2_buf_2 fanout5427 (.A(net5430),
    .X(net5427));
 sg13g2_buf_2 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_4 fanout5429 (.X(net5429),
    .A(net5430));
 sg13g2_buf_2 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_4 fanout5431 (.X(net5431),
    .A(_09209_));
 sg13g2_buf_8 fanout5432 (.A(_09169_),
    .X(net5432));
 sg13g2_buf_2 fanout5433 (.A(net5434),
    .X(net5433));
 sg13g2_buf_4 fanout5434 (.X(net5434),
    .A(net5435));
 sg13g2_buf_4 fanout5435 (.X(net5435),
    .A(net5445));
 sg13g2_buf_4 fanout5436 (.X(net5436),
    .A(net5437));
 sg13g2_buf_4 fanout5437 (.X(net5437),
    .A(net5445));
 sg13g2_buf_4 fanout5438 (.X(net5438),
    .A(net5442));
 sg13g2_buf_1 fanout5439 (.A(net5442),
    .X(net5439));
 sg13g2_buf_2 fanout5440 (.A(net5442),
    .X(net5440));
 sg13g2_buf_2 fanout5441 (.A(net5442),
    .X(net5441));
 sg13g2_buf_2 fanout5442 (.A(net5445),
    .X(net5442));
 sg13g2_buf_4 fanout5443 (.X(net5443),
    .A(net5445));
 sg13g2_buf_2 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_4 fanout5445 (.X(net5445),
    .A(_09168_));
 sg13g2_buf_4 fanout5446 (.X(net5446),
    .A(net5448));
 sg13g2_buf_4 fanout5447 (.X(net5447),
    .A(net5448));
 sg13g2_buf_4 fanout5448 (.X(net5448),
    .A(net5451));
 sg13g2_buf_4 fanout5449 (.X(net5449),
    .A(net5451));
 sg13g2_buf_2 fanout5450 (.A(net5451),
    .X(net5450));
 sg13g2_buf_2 fanout5451 (.A(_09168_),
    .X(net5451));
 sg13g2_buf_4 fanout5452 (.X(net5452),
    .A(net5454));
 sg13g2_buf_4 fanout5453 (.X(net5453),
    .A(net5454));
 sg13g2_buf_2 fanout5454 (.A(net5457),
    .X(net5454));
 sg13g2_buf_4 fanout5455 (.X(net5455),
    .A(net5457));
 sg13g2_buf_4 fanout5456 (.X(net5456),
    .A(net5457));
 sg13g2_buf_2 fanout5457 (.A(net5476),
    .X(net5457));
 sg13g2_buf_4 fanout5458 (.X(net5458),
    .A(net5460));
 sg13g2_buf_2 fanout5459 (.A(net5460),
    .X(net5459));
 sg13g2_buf_2 fanout5460 (.A(net5476),
    .X(net5460));
 sg13g2_buf_2 fanout5461 (.A(net5464),
    .X(net5461));
 sg13g2_buf_2 fanout5462 (.A(net5464),
    .X(net5462));
 sg13g2_buf_1 fanout5463 (.A(net5464),
    .X(net5463));
 sg13g2_buf_2 fanout5464 (.A(net5476),
    .X(net5464));
 sg13g2_buf_2 fanout5465 (.A(net5466),
    .X(net5465));
 sg13g2_buf_2 fanout5466 (.A(net5475),
    .X(net5466));
 sg13g2_buf_2 fanout5467 (.A(net5469),
    .X(net5467));
 sg13g2_buf_4 fanout5468 (.X(net5468),
    .A(net5469));
 sg13g2_buf_2 fanout5469 (.A(net5475),
    .X(net5469));
 sg13g2_buf_2 fanout5470 (.A(net5471),
    .X(net5470));
 sg13g2_buf_4 fanout5471 (.X(net5471),
    .A(net5475));
 sg13g2_buf_4 fanout5472 (.X(net5472),
    .A(net5474));
 sg13g2_buf_2 fanout5473 (.A(net5474),
    .X(net5473));
 sg13g2_buf_2 fanout5474 (.A(net5475),
    .X(net5474));
 sg13g2_buf_4 fanout5475 (.X(net5475),
    .A(net5476));
 sg13g2_buf_4 fanout5476 (.X(net5476),
    .A(_09168_));
 sg13g2_buf_4 fanout5477 (.X(net5477),
    .A(net5478));
 sg13g2_buf_4 fanout5478 (.X(net5478),
    .A(net5481));
 sg13g2_buf_2 fanout5479 (.A(net5481),
    .X(net5479));
 sg13g2_buf_4 fanout5480 (.X(net5480),
    .A(net5481));
 sg13g2_buf_4 fanout5481 (.X(net5481),
    .A(_09341_));
 sg13g2_buf_4 fanout5482 (.X(net5482),
    .A(net5484));
 sg13g2_buf_2 fanout5483 (.A(net5484),
    .X(net5483));
 sg13g2_buf_4 fanout5484 (.X(net5484),
    .A(net5487));
 sg13g2_buf_2 fanout5485 (.A(net5486),
    .X(net5485));
 sg13g2_buf_4 fanout5486 (.X(net5486),
    .A(net5487));
 sg13g2_buf_2 fanout5487 (.A(_09341_),
    .X(net5487));
 sg13g2_buf_4 fanout5488 (.X(net5488),
    .A(net5489));
 sg13g2_buf_2 fanout5489 (.A(net5493),
    .X(net5489));
 sg13g2_buf_4 fanout5490 (.X(net5490),
    .A(net5493));
 sg13g2_buf_4 fanout5491 (.X(net5491),
    .A(net5492));
 sg13g2_buf_8 fanout5492 (.A(net5493),
    .X(net5492));
 sg13g2_buf_8 fanout5493 (.A(_09315_),
    .X(net5493));
 sg13g2_buf_4 fanout5494 (.X(net5494),
    .A(net5500));
 sg13g2_buf_2 fanout5495 (.A(net5500),
    .X(net5495));
 sg13g2_buf_4 fanout5496 (.X(net5496),
    .A(net5497));
 sg13g2_buf_4 fanout5497 (.X(net5497),
    .A(net5500));
 sg13g2_buf_4 fanout5498 (.X(net5498),
    .A(net5499));
 sg13g2_buf_4 fanout5499 (.X(net5499),
    .A(net5500));
 sg13g2_buf_8 fanout5500 (.A(_09315_),
    .X(net5500));
 sg13g2_buf_4 fanout5501 (.X(net5501),
    .A(net5503));
 sg13g2_buf_1 fanout5502 (.A(net5503),
    .X(net5502));
 sg13g2_buf_4 fanout5503 (.X(net5503),
    .A(net5507));
 sg13g2_buf_4 fanout5504 (.X(net5504),
    .A(net5506));
 sg13g2_buf_2 fanout5505 (.A(net5506),
    .X(net5505));
 sg13g2_buf_8 fanout5506 (.A(net5507),
    .X(net5506));
 sg13g2_buf_2 fanout5507 (.A(net5513),
    .X(net5507));
 sg13g2_buf_4 fanout5508 (.X(net5508),
    .A(net5509));
 sg13g2_buf_2 fanout5509 (.A(net5510),
    .X(net5509));
 sg13g2_buf_4 fanout5510 (.X(net5510),
    .A(net5513));
 sg13g2_buf_4 fanout5511 (.X(net5511),
    .A(net5513));
 sg13g2_buf_2 fanout5512 (.A(net5513),
    .X(net5512));
 sg13g2_buf_2 fanout5513 (.A(_09292_),
    .X(net5513));
 sg13g2_buf_4 fanout5514 (.X(net5514),
    .A(_09267_));
 sg13g2_buf_4 fanout5515 (.X(net5515),
    .A(net5519));
 sg13g2_buf_4 fanout5516 (.X(net5516),
    .A(net5519));
 sg13g2_buf_4 fanout5517 (.X(net5517),
    .A(net5519));
 sg13g2_buf_2 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_8 fanout5519 (.A(_09171_),
    .X(net5519));
 sg13g2_buf_4 fanout5520 (.X(net5520),
    .A(net5522));
 sg13g2_buf_2 fanout5521 (.A(net5522),
    .X(net5521));
 sg13g2_buf_2 fanout5522 (.A(_09171_),
    .X(net5522));
 sg13g2_buf_4 fanout5523 (.X(net5523),
    .A(net5525));
 sg13g2_buf_4 fanout5524 (.X(net5524),
    .A(net5525));
 sg13g2_buf_2 fanout5525 (.A(net5526),
    .X(net5525));
 sg13g2_buf_4 fanout5526 (.X(net5526),
    .A(_09171_));
 sg13g2_buf_4 fanout5527 (.X(net5527),
    .A(net5528));
 sg13g2_buf_2 fanout5528 (.A(net5529),
    .X(net5528));
 sg13g2_buf_4 fanout5529 (.X(net5529),
    .A(_09155_));
 sg13g2_buf_4 fanout5530 (.X(net5530),
    .A(net5531));
 sg13g2_buf_2 fanout5531 (.A(net5532),
    .X(net5531));
 sg13g2_buf_4 fanout5532 (.X(net5532),
    .A(_09154_));
 sg13g2_buf_4 fanout5533 (.X(net5533),
    .A(_09126_));
 sg13g2_buf_2 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_1 fanout5535 (.A(net5536),
    .X(net5535));
 sg13g2_buf_2 fanout5536 (.A(_03024_),
    .X(net5536));
 sg13g2_buf_2 fanout5537 (.A(net5539),
    .X(net5537));
 sg13g2_buf_2 fanout5538 (.A(net5539),
    .X(net5538));
 sg13g2_buf_4 fanout5539 (.X(net5539),
    .A(_10000_));
 sg13g2_buf_2 fanout5540 (.A(net5541),
    .X(net5540));
 sg13g2_buf_4 fanout5541 (.X(net5541),
    .A(_09289_));
 sg13g2_buf_4 fanout5542 (.X(net5542),
    .A(net5543));
 sg13g2_buf_4 fanout5543 (.X(net5543),
    .A(_09260_));
 sg13g2_buf_4 fanout5544 (.X(net5544),
    .A(net5547));
 sg13g2_buf_2 fanout5545 (.A(net5546),
    .X(net5545));
 sg13g2_buf_4 fanout5546 (.X(net5546),
    .A(net5547));
 sg13g2_buf_2 fanout5547 (.A(_09259_),
    .X(net5547));
 sg13g2_buf_8 fanout5548 (.A(_09166_),
    .X(net5548));
 sg13g2_buf_4 fanout5549 (.X(net5549),
    .A(net5551));
 sg13g2_buf_2 fanout5550 (.A(net5551),
    .X(net5550));
 sg13g2_buf_4 fanout5551 (.X(net5551),
    .A(_09166_));
 sg13g2_buf_4 fanout5552 (.X(net5552),
    .A(net5554));
 sg13g2_buf_2 fanout5553 (.A(net5554),
    .X(net5553));
 sg13g2_buf_2 fanout5554 (.A(net5555),
    .X(net5554));
 sg13g2_buf_4 fanout5555 (.X(net5555),
    .A(net5556));
 sg13g2_buf_8 fanout5556 (.A(_09165_),
    .X(net5556));
 sg13g2_buf_4 fanout5557 (.X(net5557),
    .A(net5559));
 sg13g2_buf_2 fanout5558 (.A(net5559),
    .X(net5558));
 sg13g2_buf_2 fanout5559 (.A(net5560),
    .X(net5559));
 sg13g2_buf_4 fanout5560 (.X(net5560),
    .A(_09146_));
 sg13g2_buf_4 fanout5561 (.X(net5561),
    .A(net5562));
 sg13g2_buf_4 fanout5562 (.X(net5562),
    .A(net5563));
 sg13g2_buf_4 fanout5563 (.X(net5563),
    .A(_09145_));
 sg13g2_buf_4 fanout5564 (.X(net5564),
    .A(_09135_));
 sg13g2_buf_2 fanout5565 (.A(net5566),
    .X(net5565));
 sg13g2_buf_2 fanout5566 (.A(net5567),
    .X(net5566));
 sg13g2_buf_2 fanout5567 (.A(_09135_),
    .X(net5567));
 sg13g2_buf_4 fanout5568 (.X(net5568),
    .A(net5569));
 sg13g2_buf_4 fanout5569 (.X(net5569),
    .A(net5570));
 sg13g2_buf_4 fanout5570 (.X(net5570),
    .A(_09104_));
 sg13g2_buf_4 fanout5571 (.X(net5571),
    .A(net5572));
 sg13g2_buf_4 fanout5572 (.X(net5572),
    .A(_09104_));
 sg13g2_buf_2 fanout5573 (.A(_06635_),
    .X(net5573));
 sg13g2_buf_1 fanout5574 (.A(_06635_),
    .X(net5574));
 sg13g2_buf_8 fanout5575 (.A(net5579),
    .X(net5575));
 sg13g2_buf_4 fanout5576 (.X(net5576),
    .A(net5579));
 sg13g2_buf_8 fanout5577 (.A(net5578),
    .X(net5577));
 sg13g2_buf_8 fanout5578 (.A(net5579),
    .X(net5578));
 sg13g2_buf_8 fanout5579 (.A(_03060_),
    .X(net5579));
 sg13g2_buf_8 fanout5580 (.A(net5582),
    .X(net5580));
 sg13g2_buf_8 fanout5581 (.A(net5582),
    .X(net5581));
 sg13g2_buf_4 fanout5582 (.X(net5582),
    .A(_03053_));
 sg13g2_buf_8 fanout5583 (.A(_03053_),
    .X(net5583));
 sg13g2_buf_4 fanout5584 (.X(net5584),
    .A(_03053_));
 sg13g2_buf_4 fanout5585 (.X(net5585),
    .A(net5586));
 sg13g2_buf_4 fanout5586 (.X(net5586),
    .A(net5588));
 sg13g2_buf_4 fanout5587 (.X(net5587),
    .A(net5588));
 sg13g2_buf_1 fanout5588 (.A(net5605),
    .X(net5588));
 sg13g2_buf_4 fanout5589 (.X(net5589),
    .A(net5590));
 sg13g2_buf_4 fanout5590 (.X(net5590),
    .A(net5605));
 sg13g2_buf_4 fanout5591 (.X(net5591),
    .A(net5595));
 sg13g2_buf_2 fanout5592 (.A(net5595),
    .X(net5592));
 sg13g2_buf_4 fanout5593 (.X(net5593),
    .A(net5595));
 sg13g2_buf_2 fanout5594 (.A(net5595),
    .X(net5594));
 sg13g2_buf_2 fanout5595 (.A(net5605),
    .X(net5595));
 sg13g2_buf_4 fanout5596 (.X(net5596),
    .A(net5600));
 sg13g2_buf_2 fanout5597 (.A(net5600),
    .X(net5597));
 sg13g2_buf_4 fanout5598 (.X(net5598),
    .A(net5600));
 sg13g2_buf_2 fanout5599 (.A(net5600),
    .X(net5599));
 sg13g2_buf_2 fanout5600 (.A(net5605),
    .X(net5600));
 sg13g2_buf_4 fanout5601 (.X(net5601),
    .A(net5604));
 sg13g2_buf_4 fanout5602 (.X(net5602),
    .A(net5603));
 sg13g2_buf_4 fanout5603 (.X(net5603),
    .A(net5604));
 sg13g2_buf_2 fanout5604 (.A(net5605),
    .X(net5604));
 sg13g2_buf_8 fanout5605 (.A(_03052_),
    .X(net5605));
 sg13g2_buf_8 fanout5606 (.A(net5607),
    .X(net5606));
 sg13g2_buf_8 fanout5607 (.A(_03045_),
    .X(net5607));
 sg13g2_buf_4 fanout5608 (.X(net5608),
    .A(net5609));
 sg13g2_buf_8 fanout5609 (.A(net5610),
    .X(net5609));
 sg13g2_buf_4 fanout5610 (.X(net5610),
    .A(_03045_));
 sg13g2_buf_8 fanout5611 (.A(net5615),
    .X(net5611));
 sg13g2_buf_8 fanout5612 (.A(net5615),
    .X(net5612));
 sg13g2_buf_4 fanout5613 (.X(net5613),
    .A(net5615));
 sg13g2_buf_8 fanout5614 (.A(net5615),
    .X(net5614));
 sg13g2_buf_8 fanout5615 (.A(_03038_),
    .X(net5615));
 sg13g2_buf_8 fanout5616 (.A(net5621),
    .X(net5616));
 sg13g2_buf_8 fanout5617 (.A(net5620),
    .X(net5617));
 sg13g2_buf_8 fanout5618 (.A(net5620),
    .X(net5618));
 sg13g2_buf_4 fanout5619 (.X(net5619),
    .A(net5620));
 sg13g2_buf_4 fanout5620 (.X(net5620),
    .A(net5621));
 sg13g2_buf_4 fanout5621 (.X(net5621),
    .A(_09191_));
 sg13g2_buf_4 fanout5622 (.X(net5622),
    .A(net5623));
 sg13g2_buf_4 fanout5623 (.X(net5623),
    .A(net5628));
 sg13g2_buf_4 fanout5624 (.X(net5624),
    .A(net5625));
 sg13g2_buf_2 fanout5625 (.A(net5628),
    .X(net5625));
 sg13g2_buf_4 fanout5626 (.X(net5626),
    .A(net5627));
 sg13g2_buf_4 fanout5627 (.X(net5627),
    .A(net5628));
 sg13g2_buf_2 fanout5628 (.A(net5640),
    .X(net5628));
 sg13g2_buf_4 fanout5629 (.X(net5629),
    .A(net5631));
 sg13g2_buf_4 fanout5630 (.X(net5630),
    .A(net5631));
 sg13g2_buf_2 fanout5631 (.A(net5640),
    .X(net5631));
 sg13g2_buf_4 fanout5632 (.X(net5632),
    .A(net5634));
 sg13g2_buf_2 fanout5633 (.A(net5634),
    .X(net5633));
 sg13g2_buf_4 fanout5634 (.X(net5634),
    .A(net5640));
 sg13g2_buf_4 fanout5635 (.X(net5635),
    .A(net5637));
 sg13g2_buf_4 fanout5636 (.X(net5636),
    .A(net5637));
 sg13g2_buf_2 fanout5637 (.A(net5639),
    .X(net5637));
 sg13g2_buf_4 fanout5638 (.X(net5638),
    .A(net5639));
 sg13g2_buf_2 fanout5639 (.A(net5640),
    .X(net5639));
 sg13g2_buf_8 fanout5640 (.A(_03069_),
    .X(net5640));
 sg13g2_buf_8 fanout5641 (.A(net5646),
    .X(net5641));
 sg13g2_buf_8 fanout5642 (.A(net5646),
    .X(net5642));
 sg13g2_buf_8 fanout5643 (.A(net5645),
    .X(net5643));
 sg13g2_buf_8 fanout5644 (.A(net5646),
    .X(net5644));
 sg13g2_buf_4 fanout5645 (.X(net5645),
    .A(net5646));
 sg13g2_buf_4 fanout5646 (.X(net5646),
    .A(_03068_));
 sg13g2_buf_2 fanout5647 (.A(net5648),
    .X(net5647));
 sg13g2_buf_2 fanout5648 (.A(net5649),
    .X(net5648));
 sg13g2_buf_4 fanout5649 (.X(net5649),
    .A(net5651));
 sg13g2_buf_4 fanout5650 (.X(net5650),
    .A(net5651));
 sg13g2_buf_2 fanout5651 (.A(net5665),
    .X(net5651));
 sg13g2_buf_4 fanout5652 (.X(net5652),
    .A(net5656));
 sg13g2_buf_2 fanout5653 (.A(net5654),
    .X(net5653));
 sg13g2_buf_4 fanout5654 (.X(net5654),
    .A(net5656));
 sg13g2_buf_4 fanout5655 (.X(net5655),
    .A(net5656));
 sg13g2_buf_2 fanout5656 (.A(net5665),
    .X(net5656));
 sg13g2_buf_4 fanout5657 (.X(net5657),
    .A(net5659));
 sg13g2_buf_4 fanout5658 (.X(net5658),
    .A(net5659));
 sg13g2_buf_2 fanout5659 (.A(net5660),
    .X(net5659));
 sg13g2_buf_4 fanout5660 (.X(net5660),
    .A(net5665));
 sg13g2_buf_4 fanout5661 (.X(net5661),
    .A(net5662));
 sg13g2_buf_4 fanout5662 (.X(net5662),
    .A(net5664));
 sg13g2_buf_4 fanout5663 (.X(net5663),
    .A(net5664));
 sg13g2_buf_2 fanout5664 (.A(net5665),
    .X(net5664));
 sg13g2_buf_8 fanout5665 (.A(_03061_),
    .X(net5665));
 sg13g2_buf_4 fanout5666 (.X(net5666),
    .A(net5667));
 sg13g2_buf_4 fanout5667 (.X(net5667),
    .A(net5670));
 sg13g2_buf_4 fanout5668 (.X(net5668),
    .A(net5670));
 sg13g2_buf_2 fanout5669 (.A(net5670),
    .X(net5669));
 sg13g2_buf_4 fanout5670 (.X(net5670),
    .A(_03046_));
 sg13g2_buf_4 fanout5671 (.X(net5671),
    .A(net5672));
 sg13g2_buf_4 fanout5672 (.X(net5672),
    .A(net5673));
 sg13g2_buf_2 fanout5673 (.A(net5675),
    .X(net5673));
 sg13g2_buf_4 fanout5674 (.X(net5674),
    .A(net5675));
 sg13g2_buf_4 fanout5675 (.X(net5675),
    .A(_03046_));
 sg13g2_buf_4 fanout5676 (.X(net5676),
    .A(net5678));
 sg13g2_buf_2 fanout5677 (.A(net5678),
    .X(net5677));
 sg13g2_buf_4 fanout5678 (.X(net5678),
    .A(net5679));
 sg13g2_buf_4 fanout5679 (.X(net5679),
    .A(net5685));
 sg13g2_buf_4 fanout5680 (.X(net5680),
    .A(net5682));
 sg13g2_buf_2 fanout5681 (.A(net5682),
    .X(net5681));
 sg13g2_buf_4 fanout5682 (.X(net5682),
    .A(net5685));
 sg13g2_buf_8 fanout5683 (.A(net5685),
    .X(net5683));
 sg13g2_buf_4 fanout5684 (.X(net5684),
    .A(net5685));
 sg13g2_buf_8 fanout5685 (.A(_03046_),
    .X(net5685));
 sg13g2_buf_4 fanout5686 (.X(net5686),
    .A(net5689));
 sg13g2_buf_4 fanout5687 (.X(net5687),
    .A(net5688));
 sg13g2_buf_4 fanout5688 (.X(net5688),
    .A(net5689));
 sg13g2_buf_2 fanout5689 (.A(net5697),
    .X(net5689));
 sg13g2_buf_4 fanout5690 (.X(net5690),
    .A(net5691));
 sg13g2_buf_2 fanout5691 (.A(net5697),
    .X(net5691));
 sg13g2_buf_2 fanout5692 (.A(net5694),
    .X(net5692));
 sg13g2_buf_2 fanout5693 (.A(net5694),
    .X(net5693));
 sg13g2_buf_4 fanout5694 (.X(net5694),
    .A(net5697));
 sg13g2_buf_4 fanout5695 (.X(net5695),
    .A(net5696));
 sg13g2_buf_4 fanout5696 (.X(net5696),
    .A(net5697));
 sg13g2_buf_4 fanout5697 (.X(net5697),
    .A(_03039_));
 sg13g2_buf_4 fanout5698 (.X(net5698),
    .A(net5705));
 sg13g2_buf_2 fanout5699 (.A(net5705),
    .X(net5699));
 sg13g2_buf_4 fanout5700 (.X(net5700),
    .A(net5702));
 sg13g2_buf_2 fanout5701 (.A(net5702),
    .X(net5701));
 sg13g2_buf_4 fanout5702 (.X(net5702),
    .A(net5705));
 sg13g2_buf_8 fanout5703 (.A(net5705),
    .X(net5703));
 sg13g2_buf_2 fanout5704 (.A(net5705),
    .X(net5704));
 sg13g2_buf_4 fanout5705 (.X(net5705),
    .A(_03039_));
 sg13g2_buf_2 fanout5706 (.A(_10075_),
    .X(net5706));
 sg13g2_buf_2 fanout5707 (.A(net5708),
    .X(net5707));
 sg13g2_buf_2 fanout5708 (.A(_10046_),
    .X(net5708));
 sg13g2_buf_4 fanout5709 (.X(net5709),
    .A(net5711));
 sg13g2_buf_4 fanout5710 (.X(net5710),
    .A(net5711));
 sg13g2_buf_2 fanout5711 (.A(net5720),
    .X(net5711));
 sg13g2_buf_4 fanout5712 (.X(net5712),
    .A(net5720));
 sg13g2_buf_2 fanout5713 (.A(net5720),
    .X(net5713));
 sg13g2_buf_4 fanout5714 (.X(net5714),
    .A(net5717));
 sg13g2_buf_4 fanout5715 (.X(net5715),
    .A(net5717));
 sg13g2_buf_2 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_2 fanout5717 (.A(net5720),
    .X(net5717));
 sg13g2_buf_4 fanout5718 (.X(net5718),
    .A(net5719));
 sg13g2_buf_4 fanout5719 (.X(net5719),
    .A(net5720));
 sg13g2_buf_4 fanout5720 (.X(net5720),
    .A(_09192_));
 sg13g2_buf_4 fanout5721 (.X(net5721),
    .A(net5723));
 sg13g2_buf_4 fanout5722 (.X(net5722),
    .A(net5723));
 sg13g2_buf_4 fanout5723 (.X(net5723),
    .A(net5729));
 sg13g2_buf_4 fanout5724 (.X(net5724),
    .A(net5729));
 sg13g2_buf_4 fanout5725 (.X(net5725),
    .A(net5729));
 sg13g2_buf_4 fanout5726 (.X(net5726),
    .A(net5728));
 sg13g2_buf_4 fanout5727 (.X(net5727),
    .A(net5728));
 sg13g2_buf_4 fanout5728 (.X(net5728),
    .A(net5729));
 sg13g2_buf_4 fanout5729 (.X(net5729),
    .A(_09192_));
 sg13g2_buf_2 fanout5730 (.A(_08832_),
    .X(net5730));
 sg13g2_buf_2 fanout5731 (.A(net5732),
    .X(net5731));
 sg13g2_buf_2 fanout5732 (.A(_08762_),
    .X(net5732));
 sg13g2_buf_4 fanout5733 (.X(net5733),
    .A(_08752_));
 sg13g2_buf_1 fanout5734 (.A(_08752_),
    .X(net5734));
 sg13g2_buf_2 fanout5735 (.A(_08751_),
    .X(net5735));
 sg13g2_buf_4 fanout5736 (.X(net5736),
    .A(_08747_));
 sg13g2_buf_2 fanout5737 (.A(net5738),
    .X(net5737));
 sg13g2_buf_2 fanout5738 (.A(_09474_),
    .X(net5738));
 sg13g2_buf_8 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_8 fanout5740 (.A(_09199_),
    .X(net5740));
 sg13g2_buf_8 fanout5741 (.A(net5743),
    .X(net5741));
 sg13g2_buf_4 fanout5742 (.X(net5742),
    .A(net5743));
 sg13g2_buf_8 fanout5743 (.A(_09199_),
    .X(net5743));
 sg13g2_buf_8 fanout5744 (.A(net5745),
    .X(net5744));
 sg13g2_buf_8 fanout5745 (.A(net5749),
    .X(net5745));
 sg13g2_buf_4 fanout5746 (.X(net5746),
    .A(net5748));
 sg13g2_buf_4 fanout5747 (.X(net5747),
    .A(net5748));
 sg13g2_buf_8 fanout5748 (.A(net5749),
    .X(net5748));
 sg13g2_buf_8 fanout5749 (.A(_09184_),
    .X(net5749));
 sg13g2_buf_4 fanout5750 (.X(net5750),
    .A(net5753));
 sg13g2_buf_1 fanout5751 (.A(net5753),
    .X(net5751));
 sg13g2_buf_4 fanout5752 (.X(net5752),
    .A(net5753));
 sg13g2_buf_2 fanout5753 (.A(_09084_),
    .X(net5753));
 sg13g2_buf_2 fanout5754 (.A(_08733_),
    .X(net5754));
 sg13g2_buf_2 fanout5755 (.A(_08726_),
    .X(net5755));
 sg13g2_buf_2 fanout5756 (.A(net5757),
    .X(net5756));
 sg13g2_buf_2 fanout5757 (.A(_06137_),
    .X(net5757));
 sg13g2_buf_4 fanout5758 (.X(net5758),
    .A(_09646_));
 sg13g2_buf_4 fanout5759 (.X(net5759),
    .A(net5760));
 sg13g2_buf_2 fanout5760 (.A(net5761),
    .X(net5760));
 sg13g2_buf_4 fanout5761 (.X(net5761),
    .A(net5763));
 sg13g2_buf_2 fanout5762 (.A(net5763),
    .X(net5762));
 sg13g2_buf_2 fanout5763 (.A(net5779),
    .X(net5763));
 sg13g2_buf_4 fanout5764 (.X(net5764),
    .A(net5767));
 sg13g2_buf_4 fanout5765 (.X(net5765),
    .A(net5767));
 sg13g2_buf_1 fanout5766 (.A(net5767),
    .X(net5766));
 sg13g2_buf_2 fanout5767 (.A(net5779),
    .X(net5767));
 sg13g2_buf_4 fanout5768 (.X(net5768),
    .A(net5769));
 sg13g2_buf_4 fanout5769 (.X(net5769),
    .A(net5779));
 sg13g2_buf_4 fanout5770 (.X(net5770),
    .A(net5773));
 sg13g2_buf_2 fanout5771 (.A(net5773),
    .X(net5771));
 sg13g2_buf_4 fanout5772 (.X(net5772),
    .A(net5773));
 sg13g2_buf_2 fanout5773 (.A(net5778),
    .X(net5773));
 sg13g2_buf_4 fanout5774 (.X(net5774),
    .A(net5778));
 sg13g2_buf_4 fanout5775 (.X(net5775),
    .A(net5778));
 sg13g2_buf_4 fanout5776 (.X(net5776),
    .A(net5778));
 sg13g2_buf_4 fanout5777 (.X(net5777),
    .A(net5778));
 sg13g2_buf_4 fanout5778 (.X(net5778),
    .A(net5779));
 sg13g2_buf_4 fanout5779 (.X(net5779),
    .A(_09200_));
 sg13g2_buf_4 fanout5780 (.X(net5780),
    .A(net5781));
 sg13g2_buf_4 fanout5781 (.X(net5781),
    .A(net5783));
 sg13g2_buf_4 fanout5782 (.X(net5782),
    .A(net5783));
 sg13g2_buf_4 fanout5783 (.X(net5783),
    .A(net5790));
 sg13g2_buf_4 fanout5784 (.X(net5784),
    .A(net5786));
 sg13g2_buf_2 fanout5785 (.A(net5786),
    .X(net5785));
 sg13g2_buf_2 fanout5786 (.A(net5787),
    .X(net5786));
 sg13g2_buf_4 fanout5787 (.X(net5787),
    .A(net5790));
 sg13g2_buf_4 fanout5788 (.X(net5788),
    .A(net5789));
 sg13g2_buf_4 fanout5789 (.X(net5789),
    .A(net5790));
 sg13g2_buf_4 fanout5790 (.X(net5790),
    .A(_09185_));
 sg13g2_buf_4 fanout5791 (.X(net5791),
    .A(net5793));
 sg13g2_buf_4 fanout5792 (.X(net5792),
    .A(net5793));
 sg13g2_buf_2 fanout5793 (.A(net5800),
    .X(net5793));
 sg13g2_buf_4 fanout5794 (.X(net5794),
    .A(net5800));
 sg13g2_buf_2 fanout5795 (.A(net5800),
    .X(net5795));
 sg13g2_buf_4 fanout5796 (.X(net5796),
    .A(net5799));
 sg13g2_buf_4 fanout5797 (.X(net5797),
    .A(net5799));
 sg13g2_buf_4 fanout5798 (.X(net5798),
    .A(net5799));
 sg13g2_buf_2 fanout5799 (.A(net5800),
    .X(net5799));
 sg13g2_buf_4 fanout5800 (.X(net5800),
    .A(_09185_));
 sg13g2_buf_2 fanout5801 (.A(_07474_),
    .X(net5801));
 sg13g2_buf_1 fanout5802 (.A(_07474_),
    .X(net5802));
 sg13g2_buf_2 fanout5803 (.A(net5807),
    .X(net5803));
 sg13g2_buf_2 fanout5804 (.A(net5807),
    .X(net5804));
 sg13g2_buf_2 fanout5805 (.A(net5806),
    .X(net5805));
 sg13g2_buf_2 fanout5806 (.A(net5807),
    .X(net5806));
 sg13g2_buf_1 fanout5807 (.A(net5808),
    .X(net5807));
 sg13g2_buf_8 fanout5808 (.A(_05365_),
    .X(net5808));
 sg13g2_buf_2 fanout5809 (.A(net5810),
    .X(net5809));
 sg13g2_buf_2 fanout5810 (.A(net5811),
    .X(net5810));
 sg13g2_buf_2 fanout5811 (.A(_05358_),
    .X(net5811));
 sg13g2_buf_2 fanout5812 (.A(_05324_),
    .X(net5812));
 sg13g2_buf_4 fanout5813 (.X(net5813),
    .A(net5814));
 sg13g2_buf_2 fanout5814 (.A(net5815),
    .X(net5814));
 sg13g2_buf_2 fanout5815 (.A(_04869_),
    .X(net5815));
 sg13g2_buf_4 fanout5816 (.X(net5816),
    .A(_04023_));
 sg13g2_buf_2 fanout5817 (.A(net5818),
    .X(net5817));
 sg13g2_buf_2 fanout5818 (.A(net5821),
    .X(net5818));
 sg13g2_buf_2 fanout5819 (.A(net5820),
    .X(net5819));
 sg13g2_buf_2 fanout5820 (.A(net5821),
    .X(net5820));
 sg13g2_buf_2 fanout5821 (.A(_08773_),
    .X(net5821));
 sg13g2_buf_2 fanout5822 (.A(net5823),
    .X(net5822));
 sg13g2_buf_4 fanout5823 (.X(net5823),
    .A(_08772_));
 sg13g2_buf_4 fanout5824 (.X(net5824),
    .A(_08772_));
 sg13g2_buf_4 fanout5825 (.X(net5825),
    .A(\atari2600.cpu.DIMUX[6] ));
 sg13g2_buf_4 fanout5826 (.X(net5826),
    .A(\atari2600.cpu.DIMUX[3] ));
 sg13g2_buf_4 fanout5827 (.X(net5827),
    .A(\atari2600.cpu.DIMUX[2] ));
 sg13g2_buf_4 fanout5828 (.X(net5828),
    .A(net5829));
 sg13g2_buf_2 fanout5829 (.A(net5832),
    .X(net5829));
 sg13g2_buf_2 fanout5830 (.A(net5831),
    .X(net5830));
 sg13g2_buf_2 fanout5831 (.A(net5832),
    .X(net5831));
 sg13g2_buf_2 fanout5832 (.A(_08713_),
    .X(net5832));
 sg13g2_buf_2 fanout5833 (.A(net5837),
    .X(net5833));
 sg13g2_buf_2 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_2 fanout5835 (.A(net5836),
    .X(net5835));
 sg13g2_buf_2 fanout5836 (.A(net5837),
    .X(net5836));
 sg13g2_buf_2 fanout5837 (.A(_08713_),
    .X(net5837));
 sg13g2_buf_2 fanout5838 (.A(net5840),
    .X(net5838));
 sg13g2_buf_2 fanout5839 (.A(net5840),
    .X(net5839));
 sg13g2_buf_2 fanout5840 (.A(net5842),
    .X(net5840));
 sg13g2_buf_4 fanout5841 (.X(net5841),
    .A(net5842));
 sg13g2_buf_2 fanout5842 (.A(net5843),
    .X(net5842));
 sg13g2_buf_1 fanout5843 (.A(_05613_),
    .X(net5843));
 sg13g2_buf_2 fanout5844 (.A(_05282_),
    .X(net5844));
 sg13g2_buf_2 fanout5845 (.A(_04104_),
    .X(net5845));
 sg13g2_buf_2 fanout5846 (.A(_04086_),
    .X(net5846));
 sg13g2_buf_4 fanout5847 (.X(net5847),
    .A(_04081_));
 sg13g2_buf_2 fanout5848 (.A(_04056_),
    .X(net5848));
 sg13g2_buf_4 fanout5849 (.X(net5849),
    .A(_04019_));
 sg13g2_buf_2 fanout5850 (.A(net5851),
    .X(net5850));
 sg13g2_buf_2 fanout5851 (.A(net5853),
    .X(net5851));
 sg13g2_buf_2 fanout5852 (.A(net5853),
    .X(net5852));
 sg13g2_buf_4 fanout5853 (.X(net5853),
    .A(_08724_));
 sg13g2_buf_2 fanout5854 (.A(net5855),
    .X(net5854));
 sg13g2_buf_4 fanout5855 (.X(net5855),
    .A(net5857));
 sg13g2_buf_4 fanout5856 (.X(net5856),
    .A(net5857));
 sg13g2_buf_4 fanout5857 (.X(net5857),
    .A(_08723_));
 sg13g2_buf_4 fanout5858 (.X(net5858),
    .A(_08714_));
 sg13g2_buf_2 fanout5859 (.A(_08714_),
    .X(net5859));
 sg13g2_buf_2 fanout5860 (.A(net5861),
    .X(net5860));
 sg13g2_buf_2 fanout5861 (.A(net5862),
    .X(net5861));
 sg13g2_buf_2 fanout5862 (.A(net5867),
    .X(net5862));
 sg13g2_buf_2 fanout5863 (.A(net5865),
    .X(net5863));
 sg13g2_buf_2 fanout5864 (.A(net5865),
    .X(net5864));
 sg13g2_buf_2 fanout5865 (.A(net5867),
    .X(net5865));
 sg13g2_buf_4 fanout5866 (.X(net5866),
    .A(net5867));
 sg13g2_buf_2 fanout5867 (.A(_08714_),
    .X(net5867));
 sg13g2_buf_4 fanout5868 (.X(net5868),
    .A(net5869));
 sg13g2_buf_2 fanout5869 (.A(_08712_),
    .X(net5869));
 sg13g2_buf_2 fanout5870 (.A(_07686_),
    .X(net5870));
 sg13g2_buf_2 fanout5871 (.A(_05669_),
    .X(net5871));
 sg13g2_buf_2 fanout5872 (.A(_05657_),
    .X(net5872));
 sg13g2_buf_2 fanout5873 (.A(net5874),
    .X(net5873));
 sg13g2_buf_1 fanout5874 (.A(_05322_),
    .X(net5874));
 sg13g2_buf_2 fanout5875 (.A(_05265_),
    .X(net5875));
 sg13g2_buf_2 fanout5876 (.A(_04050_),
    .X(net5876));
 sg13g2_buf_4 fanout5877 (.X(net5877),
    .A(_04043_));
 sg13g2_buf_2 fanout5878 (.A(_04043_),
    .X(net5878));
 sg13g2_buf_4 fanout5879 (.X(net5879),
    .A(_04032_));
 sg13g2_buf_2 fanout5880 (.A(net5887),
    .X(net5880));
 sg13g2_buf_1 fanout5881 (.A(net5887),
    .X(net5881));
 sg13g2_buf_2 fanout5882 (.A(net5887),
    .X(net5882));
 sg13g2_buf_2 fanout5883 (.A(net5886),
    .X(net5883));
 sg13g2_buf_1 fanout5884 (.A(net5886),
    .X(net5884));
 sg13g2_buf_2 fanout5885 (.A(net5886),
    .X(net5885));
 sg13g2_buf_1 fanout5886 (.A(net5887),
    .X(net5886));
 sg13g2_buf_1 fanout5887 (.A(_03816_),
    .X(net5887));
 sg13g2_buf_2 fanout5888 (.A(_03815_),
    .X(net5888));
 sg13g2_buf_2 fanout5889 (.A(_03815_),
    .X(net5889));
 sg13g2_buf_2 fanout5890 (.A(net5891),
    .X(net5890));
 sg13g2_buf_2 fanout5891 (.A(net5892),
    .X(net5891));
 sg13g2_buf_2 fanout5892 (.A(_03815_),
    .X(net5892));
 sg13g2_buf_2 fanout5893 (.A(_03721_),
    .X(net5893));
 sg13g2_buf_4 fanout5894 (.X(net5894),
    .A(_03715_));
 sg13g2_buf_1 fanout5895 (.A(_03715_),
    .X(net5895));
 sg13g2_buf_4 fanout5896 (.X(net5896),
    .A(_03714_));
 sg13g2_buf_2 fanout5897 (.A(net5899),
    .X(net5897));
 sg13g2_buf_1 fanout5898 (.A(net5899),
    .X(net5898));
 sg13g2_buf_2 fanout5899 (.A(net5903),
    .X(net5899));
 sg13g2_buf_2 fanout5900 (.A(net5901),
    .X(net5900));
 sg13g2_buf_2 fanout5901 (.A(net5903),
    .X(net5901));
 sg13g2_buf_2 fanout5902 (.A(net5903),
    .X(net5902));
 sg13g2_buf_2 fanout5903 (.A(_03436_),
    .X(net5903));
 sg13g2_buf_2 fanout5904 (.A(net5905),
    .X(net5904));
 sg13g2_buf_4 fanout5905 (.X(net5905),
    .A(net5909));
 sg13g2_buf_2 fanout5906 (.A(net5907),
    .X(net5906));
 sg13g2_buf_2 fanout5907 (.A(net5909),
    .X(net5907));
 sg13g2_buf_2 fanout5908 (.A(net5909),
    .X(net5908));
 sg13g2_buf_2 fanout5909 (.A(_03435_),
    .X(net5909));
 sg13g2_buf_2 fanout5910 (.A(net5912),
    .X(net5910));
 sg13g2_buf_2 fanout5911 (.A(net5912),
    .X(net5911));
 sg13g2_buf_1 fanout5912 (.A(net5913),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(_08711_),
    .X(net5913));
 sg13g2_buf_2 fanout5914 (.A(_05679_),
    .X(net5914));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5916));
 sg13g2_buf_2 fanout5916 (.A(_05247_),
    .X(net5916));
 sg13g2_buf_2 fanout5917 (.A(_05236_),
    .X(net5917));
 sg13g2_buf_4 fanout5918 (.X(net5918),
    .A(_03924_));
 sg13g2_buf_2 fanout5919 (.A(_03712_),
    .X(net5919));
 sg13g2_buf_2 fanout5920 (.A(net5923),
    .X(net5920));
 sg13g2_buf_2 fanout5921 (.A(net5923),
    .X(net5921));
 sg13g2_buf_1 fanout5922 (.A(net5923),
    .X(net5922));
 sg13g2_buf_1 fanout5923 (.A(_03617_),
    .X(net5923));
 sg13g2_buf_2 fanout5924 (.A(net5926),
    .X(net5924));
 sg13g2_buf_2 fanout5925 (.A(net5926),
    .X(net5925));
 sg13g2_buf_2 fanout5926 (.A(_03524_),
    .X(net5926));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(_09077_));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(_09072_));
 sg13g2_buf_2 fanout5929 (.A(_08709_),
    .X(net5929));
 sg13g2_buf_1 fanout5930 (.A(_08709_),
    .X(net5930));
 sg13g2_buf_2 fanout5931 (.A(net5932),
    .X(net5931));
 sg13g2_buf_2 fanout5932 (.A(_07684_),
    .X(net5932));
 sg13g2_buf_2 fanout5933 (.A(net5934),
    .X(net5933));
 sg13g2_buf_2 fanout5934 (.A(_05250_),
    .X(net5934));
 sg13g2_buf_4 fanout5935 (.X(net5935),
    .A(_10009_));
 sg13g2_buf_2 fanout5936 (.A(net5937),
    .X(net5936));
 sg13g2_buf_2 fanout5937 (.A(net5938),
    .X(net5937));
 sg13g2_buf_2 fanout5938 (.A(_09109_),
    .X(net5938));
 sg13g2_buf_2 fanout5939 (.A(_09067_),
    .X(net5939));
 sg13g2_buf_4 fanout5940 (.X(net5940),
    .A(_09045_));
 sg13g2_buf_4 fanout5941 (.X(net5941),
    .A(_08135_));
 sg13g2_buf_2 fanout5942 (.A(_06136_),
    .X(net5942));
 sg13g2_buf_2 fanout5943 (.A(_06136_),
    .X(net5943));
 sg13g2_buf_2 fanout5944 (.A(_05704_),
    .X(net5944));
 sg13g2_buf_2 fanout5945 (.A(_05704_),
    .X(net5945));
 sg13g2_buf_2 fanout5946 (.A(_05545_),
    .X(net5946));
 sg13g2_buf_2 fanout5947 (.A(_05545_),
    .X(net5947));
 sg13g2_buf_2 fanout5948 (.A(_09081_),
    .X(net5948));
 sg13g2_buf_4 fanout5949 (.X(net5949),
    .A(_09065_));
 sg13g2_buf_8 fanout5950 (.A(_08297_),
    .X(net5950));
 sg13g2_buf_8 fanout5951 (.A(_08290_),
    .X(net5951));
 sg13g2_buf_8 fanout5952 (.A(_08283_),
    .X(net5952));
 sg13g2_buf_8 fanout5953 (.A(_08281_),
    .X(net5953));
 sg13g2_buf_4 fanout5954 (.X(net5954),
    .A(_08270_));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(_08265_));
 sg13g2_buf_2 fanout5956 (.A(_08265_),
    .X(net5956));
 sg13g2_buf_4 fanout5957 (.X(net5957),
    .A(_08263_));
 sg13g2_buf_4 fanout5958 (.X(net5958),
    .A(_08259_));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(_08256_));
 sg13g2_buf_4 fanout5960 (.X(net5960),
    .A(_08250_));
 sg13g2_buf_2 fanout5961 (.A(_08250_),
    .X(net5961));
 sg13g2_buf_8 fanout5962 (.A(_08241_),
    .X(net5962));
 sg13g2_buf_4 fanout5963 (.X(net5963),
    .A(net5964));
 sg13g2_buf_4 fanout5964 (.X(net5964),
    .A(_08238_));
 sg13g2_buf_8 fanout5965 (.A(_08232_),
    .X(net5965));
 sg13g2_buf_4 fanout5966 (.X(net5966),
    .A(_08229_));
 sg13g2_buf_2 fanout5967 (.A(_08229_),
    .X(net5967));
 sg13g2_buf_8 fanout5968 (.A(_08228_),
    .X(net5968));
 sg13g2_buf_8 fanout5969 (.A(_06550_),
    .X(net5969));
 sg13g2_buf_2 fanout5970 (.A(_06145_),
    .X(net5970));
 sg13g2_buf_2 fanout5971 (.A(net5972),
    .X(net5971));
 sg13g2_buf_2 fanout5972 (.A(_06134_),
    .X(net5972));
 sg13g2_buf_2 fanout5973 (.A(_06123_),
    .X(net5973));
 sg13g2_buf_2 fanout5974 (.A(_05703_),
    .X(net5974));
 sg13g2_buf_2 fanout5975 (.A(_05663_),
    .X(net5975));
 sg13g2_buf_2 fanout5976 (.A(net5979),
    .X(net5976));
 sg13g2_buf_2 fanout5977 (.A(net5978),
    .X(net5977));
 sg13g2_buf_2 fanout5978 (.A(net5979),
    .X(net5978));
 sg13g2_buf_2 fanout5979 (.A(_05544_),
    .X(net5979));
 sg13g2_buf_2 fanout5980 (.A(net5983),
    .X(net5980));
 sg13g2_buf_2 fanout5981 (.A(net5982),
    .X(net5981));
 sg13g2_buf_4 fanout5982 (.X(net5982),
    .A(net5983));
 sg13g2_buf_2 fanout5983 (.A(_03327_),
    .X(net5983));
 sg13g2_buf_4 fanout5984 (.X(net5984),
    .A(net5985));
 sg13g2_buf_2 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_2 fanout5986 (.A(_03326_),
    .X(net5986));
 sg13g2_buf_4 fanout5987 (.X(net5987),
    .A(_03326_));
 sg13g2_buf_1 fanout5988 (.A(_03326_),
    .X(net5988));
 sg13g2_buf_4 fanout5989 (.X(net5989),
    .A(_09107_));
 sg13g2_buf_4 fanout5990 (.X(net5990),
    .A(_08975_));
 sg13g2_buf_4 fanout5991 (.X(net5991),
    .A(_08919_));
 sg13g2_buf_4 fanout5992 (.X(net5992),
    .A(_08918_));
 sg13g2_buf_2 fanout5993 (.A(net5994),
    .X(net5993));
 sg13g2_buf_2 fanout5994 (.A(net5996),
    .X(net5994));
 sg13g2_buf_4 fanout5995 (.X(net5995),
    .A(net5996));
 sg13g2_buf_2 fanout5996 (.A(_08917_),
    .X(net5996));
 sg13g2_buf_4 fanout5997 (.X(net5997),
    .A(_08854_));
 sg13g2_buf_2 fanout5998 (.A(net5999),
    .X(net5998));
 sg13g2_buf_2 fanout5999 (.A(_08779_),
    .X(net5999));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6001));
 sg13g2_buf_2 fanout6001 (.A(_08243_),
    .X(net6001));
 sg13g2_buf_4 fanout6002 (.X(net6002),
    .A(_07908_));
 sg13g2_buf_1 fanout6003 (.A(_07908_),
    .X(net6003));
 sg13g2_buf_4 fanout6004 (.X(net6004),
    .A(_07834_));
 sg13g2_buf_1 fanout6005 (.A(_07834_),
    .X(net6005));
 sg13g2_buf_2 fanout6006 (.A(_06058_),
    .X(net6006));
 sg13g2_buf_2 fanout6007 (.A(_05752_),
    .X(net6007));
 sg13g2_buf_2 fanout6008 (.A(_05616_),
    .X(net6008));
 sg13g2_buf_2 fanout6009 (.A(_05615_),
    .X(net6009));
 sg13g2_buf_2 fanout6010 (.A(_05615_),
    .X(net6010));
 sg13g2_buf_4 fanout6011 (.X(net6011),
    .A(_03377_));
 sg13g2_buf_2 fanout6012 (.A(_03377_),
    .X(net6012));
 sg13g2_buf_4 fanout6013 (.X(net6013),
    .A(net6015));
 sg13g2_buf_2 fanout6014 (.A(net6015),
    .X(net6014));
 sg13g2_buf_2 fanout6015 (.A(_03330_),
    .X(net6015));
 sg13g2_buf_2 fanout6016 (.A(net6020),
    .X(net6016));
 sg13g2_buf_1 fanout6017 (.A(net6020),
    .X(net6017));
 sg13g2_buf_4 fanout6018 (.X(net6018),
    .A(net6020));
 sg13g2_buf_2 fanout6019 (.A(net6020),
    .X(net6019));
 sg13g2_buf_2 fanout6020 (.A(_03330_),
    .X(net6020));
 sg13g2_buf_2 fanout6021 (.A(net6024),
    .X(net6021));
 sg13g2_buf_2 fanout6022 (.A(net6024),
    .X(net6022));
 sg13g2_buf_2 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_2 fanout6024 (.A(_03201_),
    .X(net6024));
 sg13g2_buf_8 fanout6025 (.A(_03195_),
    .X(net6025));
 sg13g2_buf_4 fanout6026 (.X(net6026),
    .A(_03195_));
 sg13g2_buf_4 fanout6027 (.X(net6027),
    .A(_03127_));
 sg13g2_buf_2 fanout6028 (.A(_03127_),
    .X(net6028));
 sg13g2_buf_8 fanout6029 (.A(_10137_),
    .X(net6029));
 sg13g2_buf_8 fanout6030 (.A(_10137_),
    .X(net6030));
 sg13g2_buf_4 fanout6031 (.X(net6031),
    .A(_08940_));
 sg13g2_buf_2 fanout6032 (.A(net6033),
    .X(net6032));
 sg13g2_buf_2 fanout6033 (.A(_08853_),
    .X(net6033));
 sg13g2_buf_4 fanout6034 (.X(net6034),
    .A(_08770_));
 sg13g2_buf_1 fanout6035 (.A(_08770_),
    .X(net6035));
 sg13g2_buf_2 fanout6036 (.A(_07907_),
    .X(net6036));
 sg13g2_buf_2 fanout6037 (.A(_07907_),
    .X(net6037));
 sg13g2_buf_2 fanout6038 (.A(_07833_),
    .X(net6038));
 sg13g2_buf_1 fanout6039 (.A(_07833_),
    .X(net6039));
 sg13g2_buf_2 fanout6040 (.A(_07374_),
    .X(net6040));
 sg13g2_buf_2 fanout6041 (.A(_07374_),
    .X(net6041));
 sg13g2_buf_4 fanout6042 (.X(net6042),
    .A(_06072_));
 sg13g2_buf_4 fanout6043 (.X(net6043),
    .A(_05653_));
 sg13g2_buf_4 fanout6044 (.X(net6044),
    .A(net6045));
 sg13g2_buf_4 fanout6045 (.X(net6045),
    .A(net6046));
 sg13g2_buf_4 fanout6046 (.X(net6046),
    .A(_03339_));
 sg13g2_buf_4 fanout6047 (.X(net6047),
    .A(net6049));
 sg13g2_buf_4 fanout6048 (.X(net6048),
    .A(net6049));
 sg13g2_buf_8 fanout6049 (.A(net6054),
    .X(net6049));
 sg13g2_buf_4 fanout6050 (.X(net6050),
    .A(net6051));
 sg13g2_buf_4 fanout6051 (.X(net6051),
    .A(net6054));
 sg13g2_buf_4 fanout6052 (.X(net6052),
    .A(net6053));
 sg13g2_buf_4 fanout6053 (.X(net6053),
    .A(net6054));
 sg13g2_buf_4 fanout6054 (.X(net6054),
    .A(_03338_));
 sg13g2_buf_2 fanout6055 (.A(_03202_),
    .X(net6055));
 sg13g2_buf_4 fanout6056 (.X(net6056),
    .A(net6058));
 sg13g2_buf_2 fanout6057 (.A(net6058),
    .X(net6057));
 sg13g2_buf_4 fanout6058 (.X(net6058),
    .A(_03194_));
 sg13g2_buf_4 fanout6059 (.X(net6059),
    .A(net6061));
 sg13g2_buf_4 fanout6060 (.X(net6060),
    .A(net6061));
 sg13g2_buf_4 fanout6061 (.X(net6061),
    .A(_03193_));
 sg13g2_buf_4 fanout6062 (.X(net6062),
    .A(net6063));
 sg13g2_buf_4 fanout6063 (.X(net6063),
    .A(net6066));
 sg13g2_buf_4 fanout6064 (.X(net6064),
    .A(net6065));
 sg13g2_buf_4 fanout6065 (.X(net6065),
    .A(net6066));
 sg13g2_buf_8 fanout6066 (.A(_03193_),
    .X(net6066));
 sg13g2_buf_4 fanout6067 (.X(net6067),
    .A(_10071_));
 sg13g2_buf_2 fanout6068 (.A(net6069),
    .X(net6068));
 sg13g2_buf_1 fanout6069 (.A(net6070),
    .X(net6069));
 sg13g2_buf_1 fanout6070 (.A(net6071),
    .X(net6070));
 sg13g2_buf_2 fanout6071 (.A(_10044_),
    .X(net6071));
 sg13g2_buf_8 fanout6072 (.A(_10019_),
    .X(net6072));
 sg13g2_buf_4 fanout6073 (.X(net6073),
    .A(net6074));
 sg13g2_buf_4 fanout6074 (.X(net6074),
    .A(net6075));
 sg13g2_buf_4 fanout6075 (.X(net6075),
    .A(_09230_));
 sg13g2_buf_4 fanout6076 (.X(net6076),
    .A(net6077));
 sg13g2_buf_4 fanout6077 (.X(net6077),
    .A(net6078));
 sg13g2_buf_4 fanout6078 (.X(net6078),
    .A(_09229_));
 sg13g2_buf_4 fanout6079 (.X(net6079),
    .A(net6084));
 sg13g2_buf_4 fanout6080 (.X(net6080),
    .A(net6083));
 sg13g2_buf_4 fanout6081 (.X(net6081),
    .A(net6083));
 sg13g2_buf_2 fanout6082 (.A(net6083),
    .X(net6082));
 sg13g2_buf_4 fanout6083 (.X(net6083),
    .A(net6084));
 sg13g2_buf_4 fanout6084 (.X(net6084),
    .A(_09229_));
 sg13g2_buf_2 fanout6085 (.A(net6088),
    .X(net6085));
 sg13g2_buf_2 fanout6086 (.A(net6087),
    .X(net6086));
 sg13g2_buf_2 fanout6087 (.A(net6088),
    .X(net6087));
 sg13g2_buf_1 fanout6088 (.A(net6089),
    .X(net6088));
 sg13g2_buf_1 fanout6089 (.A(_09228_),
    .X(net6089));
 sg13g2_buf_2 fanout6090 (.A(net6091),
    .X(net6090));
 sg13g2_buf_4 fanout6091 (.X(net6091),
    .A(net6092));
 sg13g2_buf_8 fanout6092 (.A(_09222_),
    .X(net6092));
 sg13g2_buf_4 fanout6093 (.X(net6093),
    .A(net6094));
 sg13g2_buf_4 fanout6094 (.X(net6094),
    .A(net6101));
 sg13g2_buf_4 fanout6095 (.X(net6095),
    .A(net6100));
 sg13g2_buf_4 fanout6096 (.X(net6096),
    .A(net6100));
 sg13g2_buf_4 fanout6097 (.X(net6097),
    .A(net6100));
 sg13g2_buf_2 fanout6098 (.A(net6099),
    .X(net6098));
 sg13g2_buf_4 fanout6099 (.X(net6099),
    .A(net6100));
 sg13g2_buf_2 fanout6100 (.A(net6101),
    .X(net6100));
 sg13g2_buf_4 fanout6101 (.X(net6101),
    .A(_09221_));
 sg13g2_buf_2 fanout6102 (.A(_08784_),
    .X(net6102));
 sg13g2_buf_2 fanout6103 (.A(_08776_),
    .X(net6103));
 sg13g2_buf_4 fanout6104 (.X(net6104),
    .A(_08775_));
 sg13g2_buf_2 fanout6105 (.A(_08775_),
    .X(net6105));
 sg13g2_buf_2 fanout6106 (.A(net6107),
    .X(net6106));
 sg13g2_buf_4 fanout6107 (.X(net6107),
    .A(_08768_));
 sg13g2_buf_2 fanout6108 (.A(_08767_),
    .X(net6108));
 sg13g2_buf_4 fanout6109 (.X(net6109),
    .A(_08720_));
 sg13g2_buf_2 fanout6110 (.A(_08717_),
    .X(net6110));
 sg13g2_buf_4 fanout6111 (.X(net6111),
    .A(_08716_));
 sg13g2_buf_2 fanout6112 (.A(_08716_),
    .X(net6112));
 sg13g2_buf_4 fanout6113 (.X(net6113),
    .A(_08654_));
 sg13g2_buf_2 fanout6114 (.A(_08654_),
    .X(net6114));
 sg13g2_buf_4 fanout6115 (.X(net6115),
    .A(_08653_));
 sg13g2_buf_4 fanout6116 (.X(net6116),
    .A(_08653_));
 sg13g2_buf_4 fanout6117 (.X(net6117),
    .A(_08653_));
 sg13g2_buf_4 fanout6118 (.X(net6118),
    .A(_08632_));
 sg13g2_buf_4 fanout6119 (.X(net6119),
    .A(_08631_));
 sg13g2_buf_4 fanout6120 (.X(net6120),
    .A(_08631_));
 sg13g2_buf_4 fanout6121 (.X(net6121),
    .A(_08630_));
 sg13g2_buf_4 fanout6122 (.X(net6122),
    .A(_08628_));
 sg13g2_buf_4 fanout6123 (.X(net6123),
    .A(net6124));
 sg13g2_buf_4 fanout6124 (.X(net6124),
    .A(_08627_));
 sg13g2_buf_4 fanout6125 (.X(net6125),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_buf_2 fanout6126 (.A(net6127),
    .X(net6126));
 sg13g2_buf_4 fanout6127 (.X(net6127),
    .A(\hvsync_gen.hpos[8] ));
 sg13g2_buf_4 fanout6128 (.X(net6128),
    .A(net6130));
 sg13g2_buf_1 fanout6129 (.A(net6130),
    .X(net6129));
 sg13g2_buf_4 fanout6130 (.X(net6130),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_4 fanout6131 (.X(net6131),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_4 fanout6132 (.X(net6132),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_2 fanout6133 (.A(\hvsync_gen.hpos[5] ),
    .X(net6133));
 sg13g2_buf_2 fanout6134 (.A(net7564),
    .X(net6134));
 sg13g2_buf_4 fanout6135 (.X(net6135),
    .A(net6137));
 sg13g2_buf_4 fanout6136 (.X(net6136),
    .A(net6137));
 sg13g2_buf_4 fanout6137 (.X(net6137),
    .A(net6147));
 sg13g2_buf_4 fanout6138 (.X(net6138),
    .A(net6140));
 sg13g2_buf_2 fanout6139 (.A(net6140),
    .X(net6139));
 sg13g2_buf_4 fanout6140 (.X(net6140),
    .A(net6147));
 sg13g2_buf_4 fanout6141 (.X(net6141),
    .A(net6143));
 sg13g2_buf_4 fanout6142 (.X(net6142),
    .A(net6143));
 sg13g2_buf_2 fanout6143 (.A(net6147),
    .X(net6143));
 sg13g2_buf_4 fanout6144 (.X(net6144),
    .A(net6146));
 sg13g2_buf_4 fanout6145 (.X(net6145),
    .A(net6146));
 sg13g2_buf_2 fanout6146 (.A(net6147),
    .X(net6146));
 sg13g2_buf_4 fanout6147 (.X(net6147),
    .A(net6185));
 sg13g2_buf_4 fanout6148 (.X(net6148),
    .A(net6150));
 sg13g2_buf_4 fanout6149 (.X(net6149),
    .A(net6150));
 sg13g2_buf_2 fanout6150 (.A(net6155),
    .X(net6150));
 sg13g2_buf_4 fanout6151 (.X(net6151),
    .A(net6152));
 sg13g2_buf_4 fanout6152 (.X(net6152),
    .A(net6155));
 sg13g2_buf_4 fanout6153 (.X(net6153),
    .A(net6155));
 sg13g2_buf_2 fanout6154 (.A(net6155),
    .X(net6154));
 sg13g2_buf_2 fanout6155 (.A(net6185),
    .X(net6155));
 sg13g2_buf_4 fanout6156 (.X(net6156),
    .A(net6159));
 sg13g2_buf_4 fanout6157 (.X(net6157),
    .A(net6159));
 sg13g2_buf_4 fanout6158 (.X(net6158),
    .A(net6159));
 sg13g2_buf_2 fanout6159 (.A(net6170),
    .X(net6159));
 sg13g2_buf_4 fanout6160 (.X(net6160),
    .A(net6163));
 sg13g2_buf_2 fanout6161 (.A(net6163),
    .X(net6161));
 sg13g2_buf_4 fanout6162 (.X(net6162),
    .A(net6163));
 sg13g2_buf_2 fanout6163 (.A(net6170),
    .X(net6163));
 sg13g2_buf_4 fanout6164 (.X(net6164),
    .A(net6166));
 sg13g2_buf_4 fanout6165 (.X(net6165),
    .A(net6166));
 sg13g2_buf_4 fanout6166 (.X(net6166),
    .A(net6170));
 sg13g2_buf_4 fanout6167 (.X(net6167),
    .A(net6169));
 sg13g2_buf_4 fanout6168 (.X(net6168),
    .A(net6169));
 sg13g2_buf_4 fanout6169 (.X(net6169),
    .A(net6170));
 sg13g2_buf_4 fanout6170 (.X(net6170),
    .A(net6185));
 sg13g2_buf_4 fanout6171 (.X(net6171),
    .A(net6184));
 sg13g2_buf_1 fanout6172 (.A(net6173),
    .X(net6172));
 sg13g2_buf_4 fanout6173 (.X(net6173),
    .A(net6184));
 sg13g2_buf_4 fanout6174 (.X(net6174),
    .A(net6177));
 sg13g2_buf_2 fanout6175 (.A(net6177),
    .X(net6175));
 sg13g2_buf_4 fanout6176 (.X(net6176),
    .A(net6177));
 sg13g2_buf_2 fanout6177 (.A(net6184),
    .X(net6177));
 sg13g2_buf_4 fanout6178 (.X(net6178),
    .A(net6180));
 sg13g2_buf_4 fanout6179 (.X(net6179),
    .A(net6180));
 sg13g2_buf_2 fanout6180 (.A(net6184),
    .X(net6180));
 sg13g2_buf_4 fanout6181 (.X(net6181),
    .A(net6183));
 sg13g2_buf_4 fanout6182 (.X(net6182),
    .A(net6183));
 sg13g2_buf_4 fanout6183 (.X(net6183),
    .A(net6184));
 sg13g2_buf_4 fanout6184 (.X(net6184),
    .A(net6185));
 sg13g2_buf_4 fanout6185 (.X(net6185),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_buf_8 fanout6186 (.A(net6189),
    .X(net6186));
 sg13g2_buf_8 fanout6187 (.A(net6189),
    .X(net6187));
 sg13g2_buf_4 fanout6188 (.X(net6188),
    .A(net6189));
 sg13g2_buf_4 fanout6189 (.X(net6189),
    .A(net6202));
 sg13g2_buf_8 fanout6190 (.A(net6192),
    .X(net6190));
 sg13g2_buf_4 fanout6191 (.X(net6191),
    .A(net6192));
 sg13g2_buf_8 fanout6192 (.A(net6202),
    .X(net6192));
 sg13g2_buf_8 fanout6193 (.A(net6197),
    .X(net6193));
 sg13g2_buf_2 fanout6194 (.A(net6197),
    .X(net6194));
 sg13g2_buf_8 fanout6195 (.A(net6197),
    .X(net6195));
 sg13g2_buf_2 fanout6196 (.A(net6197),
    .X(net6196));
 sg13g2_buf_2 fanout6197 (.A(net6202),
    .X(net6197));
 sg13g2_buf_4 fanout6198 (.X(net6198),
    .A(net6201));
 sg13g2_buf_4 fanout6199 (.X(net6199),
    .A(net6201));
 sg13g2_buf_4 fanout6200 (.X(net6200),
    .A(net6201));
 sg13g2_buf_4 fanout6201 (.X(net6201),
    .A(net6202));
 sg13g2_buf_4 fanout6202 (.X(net6202),
    .A(net6210));
 sg13g2_buf_8 fanout6203 (.A(net6205),
    .X(net6203));
 sg13g2_buf_8 fanout6204 (.A(net6205),
    .X(net6204));
 sg13g2_buf_4 fanout6205 (.X(net6205),
    .A(net6210));
 sg13g2_buf_8 fanout6206 (.A(net6207),
    .X(net6206));
 sg13g2_buf_4 fanout6207 (.X(net6207),
    .A(net6210));
 sg13g2_buf_4 fanout6208 (.X(net6208),
    .A(net6209));
 sg13g2_buf_4 fanout6209 (.X(net6209),
    .A(net6210));
 sg13g2_buf_2 fanout6210 (.A(\hvsync_gen.hpos[2] ),
    .X(net6210));
 sg13g2_buf_8 fanout6211 (.A(net6214),
    .X(net6211));
 sg13g2_buf_8 fanout6212 (.A(net6214),
    .X(net6212));
 sg13g2_buf_4 fanout6213 (.X(net6213),
    .A(net6214));
 sg13g2_buf_2 fanout6214 (.A(net6228),
    .X(net6214));
 sg13g2_buf_8 fanout6215 (.A(net6220),
    .X(net6215));
 sg13g2_buf_2 fanout6216 (.A(net6220),
    .X(net6216));
 sg13g2_buf_2 fanout6217 (.A(net6219),
    .X(net6217));
 sg13g2_buf_1 fanout6218 (.A(net6219),
    .X(net6218));
 sg13g2_buf_4 fanout6219 (.X(net6219),
    .A(net6220));
 sg13g2_buf_4 fanout6220 (.X(net6220),
    .A(net6228));
 sg13g2_buf_8 fanout6221 (.A(net6223),
    .X(net6221));
 sg13g2_buf_8 fanout6222 (.A(net6223),
    .X(net6222));
 sg13g2_buf_8 fanout6223 (.A(net6228),
    .X(net6223));
 sg13g2_buf_4 fanout6224 (.X(net6224),
    .A(net6227));
 sg13g2_buf_8 fanout6225 (.A(net6227),
    .X(net6225));
 sg13g2_buf_4 fanout6226 (.X(net6226),
    .A(net6227));
 sg13g2_buf_4 fanout6227 (.X(net6227),
    .A(net6228));
 sg13g2_buf_4 fanout6228 (.X(net6228),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_2 fanout6229 (.A(net6230),
    .X(net6229));
 sg13g2_buf_4 fanout6230 (.X(net6230),
    .A(net6244));
 sg13g2_buf_8 fanout6231 (.A(net6244),
    .X(net6231));
 sg13g2_buf_4 fanout6232 (.X(net6232),
    .A(net6236));
 sg13g2_buf_4 fanout6233 (.X(net6233),
    .A(net6236));
 sg13g2_buf_8 fanout6234 (.A(net6236),
    .X(net6234));
 sg13g2_buf_4 fanout6235 (.X(net6235),
    .A(net6236));
 sg13g2_buf_2 fanout6236 (.A(net6244),
    .X(net6236));
 sg13g2_buf_4 fanout6237 (.X(net6237),
    .A(net6238));
 sg13g2_buf_8 fanout6238 (.A(net6243),
    .X(net6238));
 sg13g2_buf_8 fanout6239 (.A(net6243),
    .X(net6239));
 sg13g2_buf_8 fanout6240 (.A(net6242),
    .X(net6240));
 sg13g2_buf_8 fanout6241 (.A(net6242),
    .X(net6241));
 sg13g2_buf_8 fanout6242 (.A(net6243),
    .X(net6242));
 sg13g2_buf_4 fanout6243 (.X(net6243),
    .A(net6244));
 sg13g2_buf_4 fanout6244 (.X(net6244),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_2 fanout6245 (.A(net2983),
    .X(net6245));
 sg13g2_buf_4 fanout6246 (.X(net6246),
    .A(net7540));
 sg13g2_buf_4 fanout6247 (.X(net6247),
    .A(\atari2600.cpu.ALU.CO ));
 sg13g2_buf_4 fanout6248 (.X(net6248),
    .A(net7554));
 sg13g2_buf_2 fanout6249 (.A(net7541),
    .X(net6249));
 sg13g2_buf_2 fanout6250 (.A(net7552),
    .X(net6250));
 sg13g2_buf_4 fanout6251 (.X(net6251),
    .A(net7534));
 sg13g2_buf_4 fanout6252 (.X(net6252),
    .A(net7504));
 sg13g2_buf_4 fanout6253 (.X(net6253),
    .A(net7580));
 sg13g2_buf_2 fanout6254 (.A(net6255),
    .X(net6254));
 sg13g2_buf_2 fanout6255 (.A(net6256),
    .X(net6255));
 sg13g2_buf_2 fanout6256 (.A(\atari2600.cpu.IRHOLD_valid ),
    .X(net6256));
 sg13g2_buf_2 fanout6257 (.A(net7581),
    .X(net6257));
 sg13g2_buf_2 fanout6258 (.A(net6259),
    .X(net6258));
 sg13g2_buf_2 fanout6259 (.A(_00127_),
    .X(net6259));
 sg13g2_buf_2 fanout6260 (.A(\atari2600.tia.audf0[2] ),
    .X(net6260));
 sg13g2_buf_2 fanout6261 (.A(net7594),
    .X(net6261));
 sg13g2_buf_2 fanout6262 (.A(net7577),
    .X(net6262));
 sg13g2_buf_2 fanout6263 (.A(net7592),
    .X(net6263));
 sg13g2_buf_4 fanout6264 (.X(net6264),
    .A(\atari2600.tia.hmbl[3] ));
 sg13g2_buf_2 fanout6265 (.A(\atari2600.tia.hmm1[3] ),
    .X(net6265));
 sg13g2_buf_4 fanout6266 (.X(net6266),
    .A(\atari2600.tia.hmp1[3] ));
 sg13g2_buf_2 fanout6267 (.A(\atari2600.tia.hmp0[3] ),
    .X(net6267));
 sg13g2_buf_2 fanout6268 (.A(net7582),
    .X(net6268));
 sg13g2_buf_4 fanout6269 (.X(net6269),
    .A(\atari2600.tia.diag[61] ));
 sg13g2_buf_4 fanout6270 (.X(net6270),
    .A(\atari2600.tia.diag[60] ));
 sg13g2_buf_4 fanout6271 (.X(net6271),
    .A(net7565));
 sg13g2_buf_2 fanout6272 (.A(\atari2600.tia.diag[71] ),
    .X(net6272));
 sg13g2_buf_4 fanout6273 (.X(net6273),
    .A(\atari2600.tia.diag[69] ));
 sg13g2_buf_2 fanout6274 (.A(net7587),
    .X(net6274));
 sg13g2_buf_2 fanout6275 (.A(\atari2600.tia.diag[68] ),
    .X(net6275));
 sg13g2_buf_2 fanout6276 (.A(\atari2600.tia.diag[67] ),
    .X(net6276));
 sg13g2_buf_2 fanout6277 (.A(net6287),
    .X(net6277));
 sg13g2_buf_2 fanout6278 (.A(net6287),
    .X(net6278));
 sg13g2_buf_2 fanout6279 (.A(net6281),
    .X(net6279));
 sg13g2_buf_2 fanout6280 (.A(net6281),
    .X(net6280));
 sg13g2_buf_4 fanout6281 (.X(net6281),
    .A(net6287));
 sg13g2_buf_2 fanout6282 (.A(net6286),
    .X(net6282));
 sg13g2_buf_1 fanout6283 (.A(net6286),
    .X(net6283));
 sg13g2_buf_2 fanout6284 (.A(net6285),
    .X(net6284));
 sg13g2_buf_2 fanout6285 (.A(net6286),
    .X(net6285));
 sg13g2_buf_4 fanout6286 (.X(net6286),
    .A(net6287));
 sg13g2_buf_2 fanout6287 (.A(\atari2600.tia.vid_out[6] ),
    .X(net6287));
 sg13g2_buf_2 fanout6288 (.A(net6289),
    .X(net6288));
 sg13g2_buf_2 fanout6289 (.A(net6290),
    .X(net6289));
 sg13g2_buf_4 fanout6290 (.X(net6290),
    .A(net6305));
 sg13g2_buf_4 fanout6291 (.X(net6291),
    .A(net6295));
 sg13g2_buf_1 fanout6292 (.A(net6295),
    .X(net6292));
 sg13g2_buf_2 fanout6293 (.A(net6295),
    .X(net6293));
 sg13g2_buf_4 fanout6294 (.X(net6294),
    .A(net6295));
 sg13g2_buf_2 fanout6295 (.A(net6305),
    .X(net6295));
 sg13g2_buf_2 fanout6296 (.A(net6298),
    .X(net6296));
 sg13g2_buf_1 fanout6297 (.A(net6298),
    .X(net6297));
 sg13g2_buf_4 fanout6298 (.X(net6298),
    .A(net6304));
 sg13g2_buf_2 fanout6299 (.A(net6304),
    .X(net6299));
 sg13g2_buf_1 fanout6300 (.A(net6304),
    .X(net6300));
 sg13g2_buf_4 fanout6301 (.X(net6301),
    .A(net6303));
 sg13g2_buf_1 fanout6302 (.A(net6303),
    .X(net6302));
 sg13g2_buf_2 fanout6303 (.A(net6304),
    .X(net6303));
 sg13g2_buf_4 fanout6304 (.X(net6304),
    .A(net6305));
 sg13g2_buf_4 fanout6305 (.X(net6305),
    .A(\atari2600.tia.vid_out[6] ));
 sg13g2_buf_4 fanout6306 (.X(net6306),
    .A(net6308));
 sg13g2_buf_1 fanout6307 (.A(net6308),
    .X(net6307));
 sg13g2_buf_2 fanout6308 (.A(net6317),
    .X(net6308));
 sg13g2_buf_2 fanout6309 (.A(net6310),
    .X(net6309));
 sg13g2_buf_2 fanout6310 (.A(net6317),
    .X(net6310));
 sg13g2_buf_2 fanout6311 (.A(net6312),
    .X(net6311));
 sg13g2_buf_2 fanout6312 (.A(net6317),
    .X(net6312));
 sg13g2_buf_4 fanout6313 (.X(net6313),
    .A(net6316));
 sg13g2_buf_4 fanout6314 (.X(net6314),
    .A(net6316));
 sg13g2_buf_2 fanout6315 (.A(net6316),
    .X(net6315));
 sg13g2_buf_4 fanout6316 (.X(net6316),
    .A(net6317));
 sg13g2_buf_4 fanout6317 (.X(net6317),
    .A(\atari2600.tia.vid_out[5] ));
 sg13g2_buf_2 fanout6318 (.A(net6321),
    .X(net6318));
 sg13g2_buf_2 fanout6319 (.A(net6321),
    .X(net6319));
 sg13g2_buf_4 fanout6320 (.X(net6320),
    .A(net6321));
 sg13g2_buf_2 fanout6321 (.A(net6334),
    .X(net6321));
 sg13g2_buf_4 fanout6322 (.X(net6322),
    .A(net6323));
 sg13g2_buf_2 fanout6323 (.A(net6325),
    .X(net6323));
 sg13g2_buf_1 fanout6324 (.A(net6325),
    .X(net6324));
 sg13g2_buf_4 fanout6325 (.X(net6325),
    .A(net6334));
 sg13g2_buf_2 fanout6326 (.A(net6328),
    .X(net6326));
 sg13g2_buf_2 fanout6327 (.A(net6333),
    .X(net6327));
 sg13g2_buf_2 fanout6328 (.A(net6333),
    .X(net6328));
 sg13g2_buf_2 fanout6329 (.A(net6333),
    .X(net6329));
 sg13g2_buf_2 fanout6330 (.A(net6333),
    .X(net6330));
 sg13g2_buf_4 fanout6331 (.X(net6331),
    .A(net6332));
 sg13g2_buf_4 fanout6332 (.X(net6332),
    .A(net6333));
 sg13g2_buf_4 fanout6333 (.X(net6333),
    .A(net6334));
 sg13g2_buf_4 fanout6334 (.X(net6334),
    .A(\atari2600.tia.vid_out[5] ));
 sg13g2_buf_4 fanout6335 (.X(net6335),
    .A(net6339));
 sg13g2_buf_2 fanout6336 (.A(net6339),
    .X(net6336));
 sg13g2_buf_4 fanout6337 (.X(net6337),
    .A(net6339));
 sg13g2_buf_2 fanout6338 (.A(net6339),
    .X(net6338));
 sg13g2_buf_2 fanout6339 (.A(net6347),
    .X(net6339));
 sg13g2_buf_2 fanout6340 (.A(net6341),
    .X(net6340));
 sg13g2_buf_4 fanout6341 (.X(net6341),
    .A(net6342));
 sg13g2_buf_2 fanout6342 (.A(net6347),
    .X(net6342));
 sg13g2_buf_4 fanout6343 (.X(net6343),
    .A(net6344));
 sg13g2_buf_2 fanout6344 (.A(net6345),
    .X(net6344));
 sg13g2_buf_2 fanout6345 (.A(net6346),
    .X(net6345));
 sg13g2_buf_4 fanout6346 (.X(net6346),
    .A(net6347));
 sg13g2_buf_2 fanout6347 (.A(\atari2600.tia.vid_out[4] ),
    .X(net6347));
 sg13g2_buf_2 fanout6348 (.A(net6350),
    .X(net6348));
 sg13g2_buf_2 fanout6349 (.A(net6350),
    .X(net6349));
 sg13g2_buf_4 fanout6350 (.X(net6350),
    .A(net6364));
 sg13g2_buf_4 fanout6351 (.X(net6351),
    .A(net6355));
 sg13g2_buf_2 fanout6352 (.A(net6355),
    .X(net6352));
 sg13g2_buf_2 fanout6353 (.A(net6355),
    .X(net6353));
 sg13g2_buf_2 fanout6354 (.A(net6355),
    .X(net6354));
 sg13g2_buf_2 fanout6355 (.A(net6364),
    .X(net6355));
 sg13g2_buf_2 fanout6356 (.A(net6358),
    .X(net6356));
 sg13g2_buf_1 fanout6357 (.A(net6358),
    .X(net6357));
 sg13g2_buf_4 fanout6358 (.X(net6358),
    .A(net6364));
 sg13g2_buf_2 fanout6359 (.A(net6363),
    .X(net6359));
 sg13g2_buf_2 fanout6360 (.A(net6363),
    .X(net6360));
 sg13g2_buf_2 fanout6361 (.A(net6362),
    .X(net6361));
 sg13g2_buf_2 fanout6362 (.A(net6363),
    .X(net6362));
 sg13g2_buf_2 fanout6363 (.A(net6364),
    .X(net6363));
 sg13g2_buf_4 fanout6364 (.X(net6364),
    .A(\atari2600.tia.vid_out[4] ));
 sg13g2_buf_2 fanout6365 (.A(net6367),
    .X(net6365));
 sg13g2_buf_1 fanout6366 (.A(net6367),
    .X(net6366));
 sg13g2_buf_4 fanout6367 (.X(net6367),
    .A(net6393));
 sg13g2_buf_4 fanout6368 (.X(net6368),
    .A(net6372));
 sg13g2_buf_2 fanout6369 (.A(net6372),
    .X(net6369));
 sg13g2_buf_2 fanout6370 (.A(net6372),
    .X(net6370));
 sg13g2_buf_4 fanout6371 (.X(net6371),
    .A(net6372));
 sg13g2_buf_2 fanout6372 (.A(net6393),
    .X(net6372));
 sg13g2_buf_4 fanout6373 (.X(net6373),
    .A(net6374));
 sg13g2_buf_4 fanout6374 (.X(net6374),
    .A(net6376));
 sg13g2_buf_2 fanout6375 (.A(net6376),
    .X(net6375));
 sg13g2_buf_1 fanout6376 (.A(net6393),
    .X(net6376));
 sg13g2_buf_2 fanout6377 (.A(net6380),
    .X(net6377));
 sg13g2_buf_2 fanout6378 (.A(net6380),
    .X(net6378));
 sg13g2_buf_2 fanout6379 (.A(net6380),
    .X(net6379));
 sg13g2_buf_2 fanout6380 (.A(net6393),
    .X(net6380));
 sg13g2_buf_4 fanout6381 (.X(net6381),
    .A(net6384));
 sg13g2_buf_4 fanout6382 (.X(net6382),
    .A(net6384));
 sg13g2_buf_2 fanout6383 (.A(net6384),
    .X(net6383));
 sg13g2_buf_4 fanout6384 (.X(net6384),
    .A(net6393));
 sg13g2_buf_2 fanout6385 (.A(net6392),
    .X(net6385));
 sg13g2_buf_2 fanout6386 (.A(net6392),
    .X(net6386));
 sg13g2_buf_2 fanout6387 (.A(net6392),
    .X(net6387));
 sg13g2_buf_4 fanout6388 (.X(net6388),
    .A(net6391));
 sg13g2_buf_4 fanout6389 (.X(net6389),
    .A(net6391));
 sg13g2_buf_1 fanout6390 (.A(net6391),
    .X(net6390));
 sg13g2_buf_4 fanout6391 (.X(net6391),
    .A(net6392));
 sg13g2_buf_2 fanout6392 (.A(net6393),
    .X(net6392));
 sg13g2_buf_8 fanout6393 (.A(\atari2600.tia.vid_out[3] ),
    .X(net6393));
 sg13g2_buf_4 fanout6394 (.X(net6394),
    .A(net6395));
 sg13g2_buf_2 fanout6395 (.A(net6396),
    .X(net6395));
 sg13g2_buf_2 fanout6396 (.A(net6404),
    .X(net6396));
 sg13g2_buf_4 fanout6397 (.X(net6397),
    .A(net6398));
 sg13g2_buf_4 fanout6398 (.X(net6398),
    .A(net6400));
 sg13g2_buf_4 fanout6399 (.X(net6399),
    .A(net6400));
 sg13g2_buf_2 fanout6400 (.A(net6404),
    .X(net6400));
 sg13g2_buf_4 fanout6401 (.X(net6401),
    .A(net6404));
 sg13g2_buf_4 fanout6402 (.X(net6402),
    .A(net6403));
 sg13g2_buf_2 fanout6403 (.A(net6404),
    .X(net6403));
 sg13g2_buf_4 fanout6404 (.X(net6404),
    .A(\atari2600.tia.vid_out[2] ));
 sg13g2_buf_4 fanout6405 (.X(net6405),
    .A(net6407));
 sg13g2_buf_1 fanout6406 (.A(net6407),
    .X(net6406));
 sg13g2_buf_4 fanout6407 (.X(net6407),
    .A(net6413));
 sg13g2_buf_4 fanout6408 (.X(net6408),
    .A(net6412));
 sg13g2_buf_2 fanout6409 (.A(net6410),
    .X(net6409));
 sg13g2_buf_2 fanout6410 (.A(net6411),
    .X(net6410));
 sg13g2_buf_2 fanout6411 (.A(net6412),
    .X(net6411));
 sg13g2_buf_2 fanout6412 (.A(net6413),
    .X(net6412));
 sg13g2_buf_4 fanout6413 (.X(net6413),
    .A(\atari2600.tia.vid_out[2] ));
 sg13g2_buf_4 fanout6414 (.X(net6414),
    .A(net6416));
 sg13g2_buf_4 fanout6415 (.X(net6415),
    .A(net6416));
 sg13g2_buf_2 fanout6416 (.A(net6422),
    .X(net6416));
 sg13g2_buf_2 fanout6417 (.A(net6422),
    .X(net6417));
 sg13g2_buf_1 fanout6418 (.A(net6422),
    .X(net6418));
 sg13g2_buf_4 fanout6419 (.X(net6419),
    .A(net6421));
 sg13g2_buf_2 fanout6420 (.A(net6421),
    .X(net6420));
 sg13g2_buf_2 fanout6421 (.A(net6422),
    .X(net6421));
 sg13g2_buf_4 fanout6422 (.X(net6422),
    .A(\atari2600.tia.vid_out[2] ));
 sg13g2_buf_2 fanout6423 (.A(net6430),
    .X(net6423));
 sg13g2_buf_1 fanout6424 (.A(net6430),
    .X(net6424));
 sg13g2_buf_2 fanout6425 (.A(net6430),
    .X(net6425));
 sg13g2_buf_4 fanout6426 (.X(net6426),
    .A(net6430));
 sg13g2_buf_2 fanout6427 (.A(net6428),
    .X(net6427));
 sg13g2_buf_2 fanout6428 (.A(net6429),
    .X(net6428));
 sg13g2_buf_2 fanout6429 (.A(net6430),
    .X(net6429));
 sg13g2_buf_4 fanout6430 (.X(net6430),
    .A(\atari2600.tia.vid_out[1] ));
 sg13g2_buf_2 fanout6431 (.A(net6433),
    .X(net6431));
 sg13g2_buf_1 fanout6432 (.A(net6433),
    .X(net6432));
 sg13g2_buf_4 fanout6433 (.X(net6433),
    .A(\atari2600.tia.vid_out[1] ));
 sg13g2_buf_4 fanout6434 (.X(net6434),
    .A(net6437));
 sg13g2_buf_2 fanout6435 (.A(net6436),
    .X(net6435));
 sg13g2_buf_2 fanout6436 (.A(net6437),
    .X(net6436));
 sg13g2_buf_4 fanout6437 (.X(net6437),
    .A(net6451));
 sg13g2_buf_4 fanout6438 (.X(net6438),
    .A(net6442));
 sg13g2_buf_1 fanout6439 (.A(net6442),
    .X(net6439));
 sg13g2_buf_2 fanout6440 (.A(net6442),
    .X(net6440));
 sg13g2_buf_2 fanout6441 (.A(net6442),
    .X(net6441));
 sg13g2_buf_2 fanout6442 (.A(net6451),
    .X(net6442));
 sg13g2_buf_4 fanout6443 (.X(net6443),
    .A(net6445));
 sg13g2_buf_2 fanout6444 (.A(net6445),
    .X(net6444));
 sg13g2_buf_4 fanout6445 (.X(net6445),
    .A(net6451));
 sg13g2_buf_4 fanout6446 (.X(net6446),
    .A(net6448));
 sg13g2_buf_4 fanout6447 (.X(net6447),
    .A(net6450));
 sg13g2_buf_2 fanout6448 (.A(net6450),
    .X(net6448));
 sg13g2_buf_2 fanout6449 (.A(net6450),
    .X(net6449));
 sg13g2_buf_2 fanout6450 (.A(net6451),
    .X(net6450));
 sg13g2_buf_4 fanout6451 (.X(net6451),
    .A(\atari2600.tia.vid_out[1] ));
 sg13g2_buf_2 fanout6452 (.A(net6453),
    .X(net6452));
 sg13g2_buf_2 fanout6453 (.A(net6462),
    .X(net6453));
 sg13g2_buf_2 fanout6454 (.A(net6462),
    .X(net6454));
 sg13g2_buf_4 fanout6455 (.X(net6455),
    .A(net6456));
 sg13g2_buf_2 fanout6456 (.A(net6458),
    .X(net6456));
 sg13g2_buf_4 fanout6457 (.X(net6457),
    .A(net6458));
 sg13g2_buf_4 fanout6458 (.X(net6458),
    .A(net6462));
 sg13g2_buf_4 fanout6459 (.X(net6459),
    .A(net6461));
 sg13g2_buf_1 fanout6460 (.A(net6461),
    .X(net6460));
 sg13g2_buf_4 fanout6461 (.X(net6461),
    .A(net6462));
 sg13g2_buf_4 fanout6462 (.X(net6462),
    .A(\atari2600.tia.vid_out[0] ));
 sg13g2_buf_4 fanout6463 (.X(net6463),
    .A(net6466));
 sg13g2_buf_2 fanout6464 (.A(net6465),
    .X(net6464));
 sg13g2_buf_2 fanout6465 (.A(net6466),
    .X(net6465));
 sg13g2_buf_4 fanout6466 (.X(net6466),
    .A(net6478));
 sg13g2_buf_2 fanout6467 (.A(net6468),
    .X(net6467));
 sg13g2_buf_4 fanout6468 (.X(net6468),
    .A(net6471));
 sg13g2_buf_2 fanout6469 (.A(net6470),
    .X(net6469));
 sg13g2_buf_2 fanout6470 (.A(net6471),
    .X(net6470));
 sg13g2_buf_2 fanout6471 (.A(net6478),
    .X(net6471));
 sg13g2_buf_4 fanout6472 (.X(net6472),
    .A(net6474));
 sg13g2_buf_2 fanout6473 (.A(net6474),
    .X(net6473));
 sg13g2_buf_2 fanout6474 (.A(net6478),
    .X(net6474));
 sg13g2_buf_2 fanout6475 (.A(net6476),
    .X(net6475));
 sg13g2_buf_2 fanout6476 (.A(net6478),
    .X(net6476));
 sg13g2_buf_4 fanout6477 (.X(net6477),
    .A(net6478));
 sg13g2_buf_8 fanout6478 (.A(\atari2600.tia.vid_out[0] ),
    .X(net6478));
 sg13g2_buf_2 fanout6479 (.A(net7593),
    .X(net6479));
 sg13g2_buf_4 fanout6480 (.X(net6480),
    .A(net7591));
 sg13g2_buf_2 fanout6481 (.A(net6482),
    .X(net6481));
 sg13g2_buf_4 fanout6482 (.X(net6482),
    .A(\atari2600.tia.vid_xpos[7] ));
 sg13g2_buf_4 fanout6483 (.X(net6483),
    .A(\atari2600.tia.vid_xpos[7] ));
 sg13g2_buf_4 fanout6484 (.X(net6484),
    .A(net6485));
 sg13g2_buf_4 fanout6485 (.X(net6485),
    .A(net7590));
 sg13g2_buf_4 fanout6486 (.X(net6486),
    .A(net6489));
 sg13g2_buf_2 fanout6487 (.A(net6489),
    .X(net6487));
 sg13g2_buf_2 fanout6488 (.A(net6489),
    .X(net6488));
 sg13g2_buf_4 fanout6489 (.X(net6489),
    .A(\atari2600.tia.vid_xpos[6] ));
 sg13g2_buf_4 fanout6490 (.X(net6490),
    .A(\atari2600.tia.vid_xpos[5] ));
 sg13g2_buf_2 fanout6491 (.A(\atari2600.tia.vid_xpos[5] ),
    .X(net6491));
 sg13g2_buf_4 fanout6492 (.X(net6492),
    .A(\atari2600.tia.vid_xpos[5] ));
 sg13g2_buf_2 fanout6493 (.A(net6494),
    .X(net6493));
 sg13g2_buf_4 fanout6494 (.X(net6494),
    .A(_00145_));
 sg13g2_buf_4 fanout6495 (.X(net6495),
    .A(net6496));
 sg13g2_buf_4 fanout6496 (.X(net6496),
    .A(\atari2600.tia.vid_xpos[4] ));
 sg13g2_buf_4 fanout6497 (.X(net6497),
    .A(_00141_));
 sg13g2_buf_4 fanout6498 (.X(net6498),
    .A(net6499));
 sg13g2_buf_4 fanout6499 (.X(net6499),
    .A(net6501));
 sg13g2_buf_2 fanout6500 (.A(net6501),
    .X(net6500));
 sg13g2_buf_4 fanout6501 (.X(net6501),
    .A(\atari2600.tia.vid_xpos[3] ));
 sg13g2_buf_4 fanout6502 (.X(net6502),
    .A(\atari2600.tia.vid_xpos[2] ));
 sg13g2_buf_4 fanout6503 (.X(net6503),
    .A(\atari2600.tia.vid_xpos[2] ));
 sg13g2_buf_4 fanout6504 (.X(net6504),
    .A(net6505));
 sg13g2_buf_4 fanout6505 (.X(net6505),
    .A(\atari2600.tia.vid_xpos[1] ));
 sg13g2_buf_4 fanout6506 (.X(net6506),
    .A(\atari2600.tia.vid_xpos[0] ));
 sg13g2_buf_4 fanout6507 (.X(net6507),
    .A(\atari2600.tia.vid_xpos[0] ));
 sg13g2_buf_2 fanout6508 (.A(net6509),
    .X(net6508));
 sg13g2_buf_2 fanout6509 (.A(net7559),
    .X(net6509));
 sg13g2_buf_2 fanout6510 (.A(net7526),
    .X(net6510));
 sg13g2_buf_2 fanout6511 (.A(net7533),
    .X(net6511));
 sg13g2_buf_1 fanout6512 (.A(\atari2600.tia.p1_scale[0] ),
    .X(net6512));
 sg13g2_buf_2 fanout6513 (.A(\atari2600.cpu.state[5] ),
    .X(net6513));
 sg13g2_buf_2 fanout6514 (.A(\atari2600.cpu.state[5] ),
    .X(net6514));
 sg13g2_buf_2 fanout6515 (.A(net6516),
    .X(net6515));
 sg13g2_buf_2 fanout6516 (.A(\atari2600.cpu.state[4] ),
    .X(net6516));
 sg13g2_buf_2 fanout6517 (.A(net6518),
    .X(net6517));
 sg13g2_buf_2 fanout6518 (.A(\atari2600.cpu.state[3] ),
    .X(net6518));
 sg13g2_buf_2 fanout6519 (.A(\atari2600.cpu.state[2] ),
    .X(net6519));
 sg13g2_buf_2 fanout6520 (.A(\atari2600.cpu.state[1] ),
    .X(net6520));
 sg13g2_buf_2 fanout6521 (.A(\atari2600.cpu.state[0] ),
    .X(net6521));
 sg13g2_buf_4 fanout6522 (.X(net6522),
    .A(net6523));
 sg13g2_buf_4 fanout6523 (.X(net6523),
    .A(net6524));
 sg13g2_buf_4 fanout6524 (.X(net6524),
    .A(net6542));
 sg13g2_buf_2 fanout6525 (.A(net6526),
    .X(net6525));
 sg13g2_buf_2 fanout6526 (.A(net6527),
    .X(net6526));
 sg13g2_buf_2 fanout6527 (.A(net6542),
    .X(net6527));
 sg13g2_buf_4 fanout6528 (.X(net6528),
    .A(net6532));
 sg13g2_buf_1 fanout6529 (.A(net6532),
    .X(net6529));
 sg13g2_buf_4 fanout6530 (.X(net6530),
    .A(net6531));
 sg13g2_buf_2 fanout6531 (.A(net6532),
    .X(net6531));
 sg13g2_buf_2 fanout6532 (.A(net6542),
    .X(net6532));
 sg13g2_buf_4 fanout6533 (.X(net6533),
    .A(net6535));
 sg13g2_buf_2 fanout6534 (.A(net6535),
    .X(net6534));
 sg13g2_buf_4 fanout6535 (.X(net6535),
    .A(net6542));
 sg13g2_buf_2 fanout6536 (.A(net6538),
    .X(net6536));
 sg13g2_buf_1 fanout6537 (.A(net6538),
    .X(net6537));
 sg13g2_buf_2 fanout6538 (.A(net6539),
    .X(net6538));
 sg13g2_buf_4 fanout6539 (.X(net6539),
    .A(net6540));
 sg13g2_buf_2 fanout6540 (.A(net6541),
    .X(net6540));
 sg13g2_buf_2 fanout6541 (.A(net6542),
    .X(net6541));
 sg13g2_buf_8 fanout6542 (.A(_08617_),
    .X(net6542));
 sg13g2_buf_4 fanout6543 (.X(net6543),
    .A(net6545));
 sg13g2_buf_4 fanout6544 (.X(net6544),
    .A(net6545));
 sg13g2_buf_2 fanout6545 (.A(net6546),
    .X(net6545));
 sg13g2_buf_4 fanout6546 (.X(net6546),
    .A(net6549));
 sg13g2_buf_4 fanout6547 (.X(net6547),
    .A(net6548));
 sg13g2_buf_2 fanout6548 (.A(net6549),
    .X(net6548));
 sg13g2_buf_4 fanout6549 (.X(net6549),
    .A(rst_n));
 sg13g2_buf_2 fanout6550 (.A(net6551),
    .X(net6550));
 sg13g2_buf_2 fanout6551 (.A(net6554),
    .X(net6551));
 sg13g2_buf_2 fanout6552 (.A(net6554),
    .X(net6552));
 sg13g2_buf_2 fanout6553 (.A(net6554),
    .X(net6553));
 sg13g2_buf_2 fanout6554 (.A(net6560),
    .X(net6554));
 sg13g2_buf_2 fanout6555 (.A(net6560),
    .X(net6555));
 sg13g2_buf_2 fanout6556 (.A(net6557),
    .X(net6556));
 sg13g2_buf_2 fanout6557 (.A(net6559),
    .X(net6557));
 sg13g2_buf_4 fanout6558 (.X(net6558),
    .A(net6559));
 sg13g2_buf_2 fanout6559 (.A(net6560),
    .X(net6559));
 sg13g2_buf_2 fanout6560 (.A(net6578),
    .X(net6560));
 sg13g2_buf_4 fanout6561 (.X(net6561),
    .A(net6562));
 sg13g2_buf_2 fanout6562 (.A(net6564),
    .X(net6562));
 sg13g2_buf_4 fanout6563 (.X(net6563),
    .A(net6564));
 sg13g2_buf_2 fanout6564 (.A(net6578),
    .X(net6564));
 sg13g2_buf_4 fanout6565 (.X(net6565),
    .A(net6566));
 sg13g2_buf_2 fanout6566 (.A(net6578),
    .X(net6566));
 sg13g2_buf_2 fanout6567 (.A(net6569),
    .X(net6567));
 sg13g2_buf_2 fanout6568 (.A(net6577),
    .X(net6568));
 sg13g2_buf_1 fanout6569 (.A(net6577),
    .X(net6569));
 sg13g2_buf_2 fanout6570 (.A(net6571),
    .X(net6570));
 sg13g2_buf_2 fanout6571 (.A(net6572),
    .X(net6571));
 sg13g2_buf_4 fanout6572 (.X(net6572),
    .A(net6577));
 sg13g2_buf_2 fanout6573 (.A(net6574),
    .X(net6573));
 sg13g2_buf_2 fanout6574 (.A(net6576),
    .X(net6574));
 sg13g2_buf_2 fanout6575 (.A(net6576),
    .X(net6575));
 sg13g2_buf_4 fanout6576 (.X(net6576),
    .A(net6577));
 sg13g2_buf_2 fanout6577 (.A(net6578),
    .X(net6577));
 sg13g2_buf_4 fanout6578 (.X(net6578),
    .A(rst_n));
 sg13g2_buf_2 fanout6579 (.A(net6581),
    .X(net6579));
 sg13g2_buf_1 fanout6580 (.A(net6581),
    .X(net6580));
 sg13g2_buf_2 fanout6581 (.A(net6582),
    .X(net6581));
 sg13g2_buf_2 fanout6582 (.A(rst_n),
    .X(net6582));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_tiehi _30422__13 (.L_HI(net13));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_leaf_260_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_2 clkbuf_leaf_261_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_2 clkbuf_leaf_262_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_2 clkbuf_leaf_263_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_2 clkbuf_leaf_264_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_2 clkbuf_leaf_265_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_2 clkbuf_leaf_266_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_2 clkbuf_leaf_267_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_2 clkbuf_leaf_268_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_2 clkbuf_leaf_269_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_2 clkbuf_leaf_270_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_2 clkbuf_leaf_271_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_2 clkbuf_leaf_272_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_2 clkbuf_leaf_273_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_2 clkbuf_leaf_274_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_2 clkbuf_leaf_275_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_2 clkbuf_leaf_276_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_2 clkbuf_leaf_277_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_2 clkbuf_leaf_278_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_2 clkbuf_leaf_279_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_2 clkbuf_leaf_280_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_2 clkbuf_leaf_281_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_2 clkbuf_leaf_282_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_2 clkbuf_leaf_283_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_2 clkbuf_leaf_284_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_2 clkbuf_leaf_285_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_2 clkbuf_leaf_286_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_2 clkbuf_leaf_287_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_2 clkbuf_leaf_288_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_2 clkbuf_leaf_289_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_2 clkbuf_leaf_290_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_2 clkbuf_leaf_291_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_2 clkbuf_leaf_292_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_2 clkbuf_leaf_293_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_2 clkbuf_leaf_294_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_2 clkbuf_leaf_295_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_2 clkbuf_leaf_296_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_2 clkbuf_leaf_297_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_2 clkbuf_leaf_298_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_2 clkbuf_leaf_299_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_2 clkbuf_leaf_300_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_2 clkbuf_leaf_301_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_2 clkbuf_leaf_302_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_2 clkbuf_leaf_303_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_2 clkbuf_leaf_304_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_2 clkbuf_leaf_305_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_2 clkbuf_leaf_306_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_2 clkbuf_leaf_307_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_2 clkbuf_leaf_308_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_2 clkbuf_leaf_309_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_2 clkbuf_leaf_310_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_2 clkbuf_leaf_311_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_2 clkbuf_leaf_312_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_2 clkbuf_leaf_313_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_2 clkbuf_leaf_314_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_2 clkbuf_leaf_315_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_2 clkbuf_leaf_316_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_2 clkbuf_leaf_317_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_2 clkbuf_leaf_318_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_2 clkbuf_leaf_319_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_2 clkbuf_leaf_320_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_2 clkbuf_leaf_321_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_2 clkbuf_leaf_322_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_2 clkbuf_leaf_323_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_2 clkbuf_leaf_324_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_2 clkbuf_leaf_325_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_2 clkbuf_leaf_326_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_2 clkbuf_leaf_327_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_327_clk));
 sg13g2_buf_2 clkbuf_leaf_328_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_328_clk));
 sg13g2_buf_2 clkbuf_leaf_329_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_329_clk));
 sg13g2_buf_2 clkbuf_leaf_330_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_330_clk));
 sg13g2_buf_2 clkbuf_leaf_331_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_331_clk));
 sg13g2_buf_2 clkbuf_leaf_332_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_332_clk));
 sg13g2_buf_2 clkbuf_leaf_333_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_333_clk));
 sg13g2_buf_2 clkbuf_leaf_334_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_334_clk));
 sg13g2_buf_2 clkbuf_leaf_335_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_335_clk));
 sg13g2_buf_2 clkbuf_leaf_336_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_336_clk));
 sg13g2_buf_2 clkbuf_leaf_337_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_337_clk));
 sg13g2_buf_2 clkbuf_leaf_338_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_338_clk));
 sg13g2_buf_2 clkbuf_leaf_339_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_339_clk));
 sg13g2_buf_2 clkbuf_leaf_340_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_340_clk));
 sg13g2_buf_2 clkbuf_leaf_341_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_341_clk));
 sg13g2_buf_2 clkbuf_leaf_342_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_342_clk));
 sg13g2_buf_2 clkbuf_leaf_343_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_343_clk));
 sg13g2_buf_2 clkbuf_leaf_344_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_344_clk));
 sg13g2_buf_2 clkbuf_leaf_345_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_345_clk));
 sg13g2_buf_2 clkbuf_leaf_346_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_346_clk));
 sg13g2_buf_2 clkbuf_leaf_347_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_347_clk));
 sg13g2_buf_2 clkbuf_leaf_348_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_348_clk));
 sg13g2_buf_2 clkbuf_leaf_349_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_349_clk));
 sg13g2_buf_2 clkbuf_leaf_350_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_350_clk));
 sg13g2_buf_2 clkbuf_leaf_351_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_351_clk));
 sg13g2_buf_2 clkbuf_leaf_352_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_352_clk));
 sg13g2_buf_2 clkbuf_leaf_353_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_353_clk));
 sg13g2_buf_2 clkbuf_leaf_354_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_354_clk));
 sg13g2_buf_2 clkbuf_leaf_355_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_355_clk));
 sg13g2_buf_2 clkbuf_leaf_356_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_356_clk));
 sg13g2_buf_2 clkbuf_leaf_357_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_357_clk));
 sg13g2_buf_2 clkbuf_leaf_358_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_358_clk));
 sg13g2_buf_2 clkbuf_leaf_359_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_359_clk));
 sg13g2_buf_2 clkbuf_leaf_360_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_360_clk));
 sg13g2_buf_2 clkbuf_leaf_361_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_361_clk));
 sg13g2_buf_2 clkbuf_leaf_362_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_362_clk));
 sg13g2_buf_2 clkbuf_leaf_363_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_363_clk));
 sg13g2_buf_2 clkbuf_leaf_364_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_364_clk));
 sg13g2_buf_2 clkbuf_leaf_365_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_365_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_6_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_2 clkbuf_6_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkbuf_6_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_2 clkbuf_6_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkbuf_6_4__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_2 clkbuf_6_5__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_2 clkbuf_6_6__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_2 clkbuf_6_7__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkbuf_6_8__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_2 clkbuf_6_9__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkbuf_6_10__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_2 clkbuf_6_11__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkbuf_6_12__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_2 clkbuf_6_13__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkbuf_6_14__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_2 clkbuf_6_15__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkbuf_6_16__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_2 clkbuf_6_17__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkbuf_6_18__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_2 clkbuf_6_19__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkbuf_6_20__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_2 clkbuf_6_21__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_2 clkbuf_6_22__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_2 clkbuf_6_23__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkbuf_6_24__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_2 clkbuf_6_25__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_2 clkbuf_6_26__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_2 clkbuf_6_27__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkbuf_6_28__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_2 clkbuf_6_29__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkbuf_6_30__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_2 clkbuf_6_31__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkbuf_6_32__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_2 clkbuf_6_33__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkbuf_6_34__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_2 clkbuf_6_35__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkbuf_6_36__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_2 clkbuf_6_37__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_2 clkbuf_6_38__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_2 clkbuf_6_39__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkbuf_6_40__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_2 clkbuf_6_41__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkbuf_6_42__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_2 clkbuf_6_43__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkbuf_6_44__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_2 clkbuf_6_45__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkbuf_6_46__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_2 clkbuf_6_47__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkbuf_6_48__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_2 clkbuf_6_49__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_2 clkbuf_6_50__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_2 clkbuf_6_51__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkbuf_6_52__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_2 clkbuf_6_53__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_2 clkbuf_6_54__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_2 clkbuf_6_55__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkbuf_6_56__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_2 clkbuf_6_57__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_2 clkbuf_6_58__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_2 clkbuf_6_59__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkbuf_6_60__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_2 clkbuf_6_61__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkbuf_6_62__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_2 clkbuf_6_63__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkload16 (.A(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkload17 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_8 clkload18 (.A(clknet_leaf_364_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_365_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_296_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad_pmod.driver.pmod_latch_sync[1] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00169_),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold4 (.A(\atari2600.tia.vid_vsync ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold5 (.A(\flash_rom.data_ready ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00167_),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00347_),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00168_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold9 (.A(_01508_),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold10 (.A(\gamepad_pmod.driver.pmod_latch_sync[0] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold11 (.A(\gamepad_pmod.driver.pmod_clk_sync[0] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00157_),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold13 (.A(\gamepad_pmod.driver.pmod_data_sync[0] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold14 (.A(\atari2600.clk_counter[2] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold15 (.A(\atari2600.clk_counter[3] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold16 (.A(\atari2600.tia.audio_right_counter[15] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold17 (.A(_01022_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold18 (.A(\atari2600.clk_counter[6] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold19 (.A(\atari2600.cpu.res ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold20 (.A(_01384_),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold21 (.A(\atari2600.clk_counter[7] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold22 (.A(_00158_),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold23 (.A(_00047_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold24 (.A(\atari2600.clk_counter[4] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold25 (.A(\atari2600.tia.audio_left_counter[15] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold26 (.A(_01006_),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold27 (.A(\atari2600.clk_counter[5] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold28 (.A(\gamepad_pmod.driver.pmod_data_sync[1] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold29 (.A(_01476_),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold30 (.A(\atari2600.tia.audio_right_counter[7] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold31 (.A(_01014_),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold32 (.A(\atari2600.tia.cx[14] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold33 (.A(_10062_),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold34 (.A(\flash_rom.addr[2] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold35 (.A(\atari2600.ram[51][7] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00162_),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold37 (.A(_00053_),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold38 (.A(\atari2600.tia.audio_left_counter[14] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold39 (.A(_01005_),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold40 (.A(\atari2600.ram[51][4] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold41 (.A(\atari2600.ram[51][2] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold42 (.A(\atari2600.tia.cx[1] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold43 (.A(_09475_),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold44 (.A(\atari2600.ram[51][5] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold45 (.A(\atari2600.tia.cx[7] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold46 (.A(_00035_),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold47 (.A(\atari2600.tia.audio_right_counter[13] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold48 (.A(_01020_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold49 (.A(\atari2600.ram[51][1] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold50 (.A(\flash_rom.addr[0] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold51 (.A(\flash_rom.addr[3] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold52 (.A(\atari2600.tia.p0_copies[2] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold53 (.A(\atari2600.ram[51][0] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold54 (.A(\atari2600.tia.cx[2] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold55 (.A(_00030_),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold56 (.A(\flash_rom.fsm_state[2] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold57 (.A(_09038_),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold58 (.A(\flash_rom.addr[1] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold59 (.A(\atari2600.tia.audio_left_counter[11] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold60 (.A(_01002_),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold61 (.A(\r_pwm_odd[2] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold62 (.A(\flash_rom.addr[12] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold63 (.A(_00975_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold64 (.A(\g_pwm_odd[2] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold65 (.A(\atari2600.tia.cx[9] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold66 (.A(_00037_),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold67 (.A(\flash_rom.addr_in[16] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00963_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold69 (.A(\atari2600.tia.audio_right_counter[9] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold70 (.A(_01016_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold71 (.A(\atari2600.tia.cx[0] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold72 (.A(\atari2600.tia.cx[13] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold73 (.A(_10061_),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold74 (.A(\atari2600.ram[41][0] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold75 (.A(\atari2600.tia.audio_right_counter[11] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold76 (.A(_01018_),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold77 (.A(\atari2600.ram[29][7] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold78 (.A(\atari2600.ram[77][6] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold79 (.A(\atari2600.ram[84][6] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold80 (.A(\atari2600.cpu.cli ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold81 (.A(_01358_),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold82 (.A(\atari2600.ram[16][0] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold83 (.A(\atari2600.ram[76][6] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold84 (.A(\atari2600.tia.audio_right_counter[14] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold85 (.A(_01021_),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold86 (.A(\atari2600.ram[101][0] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold87 (.A(\atari2600.ram[48][5] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold88 (.A(\atari2600.ram[49][3] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00057_),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold90 (.A(_08210_),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold91 (.A(\atari2600.ram[9][5] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold92 (.A(\atari2600.tia.audio_left_counter[3] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold93 (.A(_00994_),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold94 (.A(\atari2600.ram[80][4] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold95 (.A(\atari2600.ram[53][3] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold96 (.A(\atari2600.ram[40][7] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold97 (.A(\atari2600.ram[81][4] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold98 (.A(\atari2600.ram[5][4] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold99 (.A(\atari2600.ram[5][1] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold100 (.A(\atari2600.tia.audio_right_counter[5] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold101 (.A(_01012_),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold102 (.A(\atari2600.ram[60][1] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold103 (.A(\atari2600.ram[4][2] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold104 (.A(\atari2600.ram[120][3] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold105 (.A(\atari2600.ram[8][5] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold106 (.A(\atari2600.ram[32][4] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold107 (.A(\atari2600.ram[41][5] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold108 (.A(\atari2600.ram[51][3] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold109 (.A(\atari2600.ram[61][3] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold110 (.A(\atari2600.ram[0][0] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold111 (.A(\atari2600.ram[0][7] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold112 (.A(\atari2600.ram[96][0] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold113 (.A(\atari2600.ram[1][4] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold114 (.A(\atari2600.ram[0][2] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold115 (.A(\atari2600.ram[88][0] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold116 (.A(\atari2600.tia.audio_right_counter[8] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold117 (.A(_01015_),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold118 (.A(\atari2600.ram[69][0] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold119 (.A(\atari2600.ram[40][3] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold120 (.A(\atari2600.ram[116][6] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold121 (.A(\atari2600.ram[49][6] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold122 (.A(\flash_rom.addr[14] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold123 (.A(_00977_),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold124 (.A(\atari2600.ram[92][5] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold125 (.A(\atari2600.ram[125][7] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold126 (.A(\atari2600.ram[12][6] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold127 (.A(\atari2600.ram[116][4] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold128 (.A(\atari2600.ram[117][2] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold129 (.A(\atari2600.ram[80][3] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold130 (.A(\atari2600.ram[13][5] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold131 (.A(\atari2600.ram[41][2] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold132 (.A(\atari2600.ram[24][5] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold133 (.A(\atari2600.ram[45][4] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold134 (.A(\atari2600.ram[20][3] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold135 (.A(\atari2600.ram[105][4] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold136 (.A(\atari2600.ram[104][1] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold137 (.A(\atari2600.ram[112][2] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold138 (.A(_00129_),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold139 (.A(_07805_),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold140 (.A(_01450_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold141 (.A(\atari2600.ram[57][6] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold142 (.A(\atari2600.ram[16][2] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold143 (.A(\atari2600.ram[88][3] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold144 (.A(\atari2600.ram[32][3] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold145 (.A(\atari2600.ram[9][1] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold146 (.A(\atari2600.ram[101][7] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold147 (.A(\atari2600.tia.cx[3] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00031_),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold149 (.A(\atari2600.ram[21][5] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold150 (.A(\atari2600.ram[56][2] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold151 (.A(\atari2600.ram[20][0] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold152 (.A(\atari2600.ram[17][0] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold153 (.A(\atari2600.ram[57][5] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold154 (.A(\atari2600.ram[93][5] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold155 (.A(\atari2600.ram[62][7] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold156 (.A(\atari2600.ram[77][0] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold157 (.A(\atari2600.ram[108][3] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold158 (.A(\atari2600.ram[8][1] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold159 (.A(\atari2600.ram[124][0] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold160 (.A(\atari2600.ram[51][6] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold161 (.A(\atari2600.ram[1][0] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold162 (.A(\atari2600.ram[104][6] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold163 (.A(\atari2600.ram[8][7] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold164 (.A(\atari2600.tia.audio_right_counter[3] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold165 (.A(_01010_),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold166 (.A(\atari2600.ram[125][3] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold167 (.A(\atari2600.ram[29][0] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold168 (.A(\atari2600.ram[118][7] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold169 (.A(\atari2600.ram[29][2] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold170 (.A(\atari2600.ram[53][1] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold171 (.A(\atari2600.ram[50][4] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold172 (.A(\atari2600.ram[17][1] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold173 (.A(\atari2600.ram[96][4] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold174 (.A(\atari2600.ram[120][0] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold175 (.A(\atari2600.ram[9][6] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold176 (.A(\atari2600.ram[48][7] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold177 (.A(\atari2600.ram[37][4] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold178 (.A(\atari2600.ram[37][2] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold179 (.A(\atari2600.tia.audio_left_counter[5] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00996_),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold181 (.A(\atari2600.ram[76][7] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold182 (.A(\atari2600.ram[46][6] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold183 (.A(\atari2600.ram[112][0] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold184 (.A(\atari2600.ram[96][1] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold185 (.A(\atari2600.ram[49][0] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold186 (.A(\atari2600.ram[70][2] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold187 (.A(_00159_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00048_),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold189 (.A(\atari2600.ram[81][0] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold190 (.A(\atari2600.ram[0][1] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold191 (.A(\atari2600.tia.audio_left_counter[9] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold192 (.A(_01000_),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold193 (.A(\atari2600.ram[24][2] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold194 (.A(\atari2600.pia.instat[0] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold195 (.A(_01240_),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold196 (.A(\atari2600.ram[65][6] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold197 (.A(\atari2600.ram[41][3] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold198 (.A(\atari2600.ram[34][6] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold199 (.A(\atari2600.ram[30][1] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold200 (.A(\atari2600.ram[29][4] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold201 (.A(\atari2600.ram[93][0] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold202 (.A(\atari2600.ram[125][2] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold203 (.A(\atari2600.ram[76][2] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold204 (.A(\atari2600.ram[81][6] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold205 (.A(\atari2600.ram[41][7] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold206 (.A(\atari2600.ram[100][6] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold207 (.A(\atari2600.ram[108][6] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold208 (.A(\atari2600.ram[109][2] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold209 (.A(\atari2600.ram[101][6] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold210 (.A(\atari2600.tia.audio_left_counter[6] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold211 (.A(_00997_),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold212 (.A(\atari2600.ram[85][3] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold213 (.A(\atari2600.ram[1][2] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold214 (.A(\atari2600.ram[65][7] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold215 (.A(\atari2600.ram[13][1] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold216 (.A(\atari2600.ram[121][6] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold217 (.A(_00058_),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold218 (.A(_08214_),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold219 (.A(\atari2600.ram[72][4] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold220 (.A(\atari2600.ram[109][4] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold221 (.A(\atari2600.ram[105][0] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold222 (.A(\atari2600.ram[33][4] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold223 (.A(\atari2600.ram[68][1] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold224 (.A(\atari2600.ram[8][4] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold225 (.A(\atari2600.ram[72][2] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold226 (.A(\atari2600.ram[12][1] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold227 (.A(\atari2600.cpu.src_reg[1] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold228 (.A(\atari2600.ram[108][4] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold229 (.A(\atari2600.ram[81][1] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold230 (.A(\atari2600.ram[108][0] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold231 (.A(\atari2600.ram[64][4] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold232 (.A(\atari2600.ram[100][4] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold233 (.A(\atari2600.ram[69][1] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold234 (.A(\scanline[102][5] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold235 (.A(\atari2600.ram[120][2] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold236 (.A(\atari2600.ram[57][3] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold237 (.A(\atari2600.ram[57][2] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold238 (.A(\atari2600.ram[94][0] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold239 (.A(\atari2600.cpu.AXYS[3][2] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold240 (.A(\atari2600.ram[80][2] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold241 (.A(\atari2600.ram[89][6] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold242 (.A(\atari2600.ram[112][6] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold243 (.A(\atari2600.ram[121][1] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold244 (.A(\atari2600.ram[126][7] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold245 (.A(\atari2600.ram[69][3] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold246 (.A(\atari2600.ram[12][2] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold247 (.A(\atari2600.ram[3][4] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold248 (.A(\atari2600.tia.audio_right_counter[12] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold249 (.A(_01019_),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold250 (.A(\atari2600.ram[56][5] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold251 (.A(\atari2600.ram[36][1] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold252 (.A(\atari2600.ram[1][3] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold253 (.A(\atari2600.ram[62][1] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold254 (.A(\atari2600.ram[94][7] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold255 (.A(\atari2600.ram[81][3] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold256 (.A(\atari2600.ram[118][4] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold257 (.A(\atari2600.ram[18][0] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold258 (.A(\atari2600.ram[12][4] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold259 (.A(\atari2600.ram[120][4] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold260 (.A(\atari2600.ram[82][1] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold261 (.A(\atari2600.ram[14][4] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold262 (.A(\atari2600.ram[93][2] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold263 (.A(\atari2600.ram[12][5] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold264 (.A(\atari2600.ram[4][0] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold265 (.A(\atari2600.ram[93][4] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold266 (.A(\atari2600.ram[40][0] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold267 (.A(\atari2600.ram[124][4] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold268 (.A(\atari2600.ram[20][7] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold269 (.A(\atari2600.ram[24][4] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold270 (.A(\atari2600.ram[44][7] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold271 (.A(\atari2600.ram[80][0] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold272 (.A(\atari2600.pia.swb_dir[4] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold273 (.A(\atari2600.ram[30][7] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold274 (.A(\atari2600.ram[16][7] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold275 (.A(\atari2600.ram[34][7] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold276 (.A(\atari2600.cpu.ALU.BI7 ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold277 (.A(\atari2600.ram[25][0] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold278 (.A(\atari2600.ram[77][3] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold279 (.A(\atari2600.ram[97][3] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold280 (.A(\atari2600.ram[85][2] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold281 (.A(\atari2600.cpu.sed ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold282 (.A(\atari2600.ram[105][5] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold283 (.A(\atari2600.ram[89][1] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold284 (.A(\atari2600.ram[2][0] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold285 (.A(\atari2600.tia.audio_left_counter[13] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold286 (.A(_01004_),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold287 (.A(\flash_rom.addr[15] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold288 (.A(_00978_),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold289 (.A(\atari2600.ram[28][0] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold290 (.A(\atari2600.ram[122][6] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold291 (.A(\atari2600.ram[16][5] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold292 (.A(\atari2600.ram[66][5] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold293 (.A(\atari2600.ram[65][5] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold294 (.A(\atari2600.ram[82][6] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold295 (.A(\atari2600.ram[8][0] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold296 (.A(\atari2600.ram[38][4] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold297 (.A(\atari2600.ram[89][2] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold298 (.A(\gamepad_pmod.decoder.data_reg[0] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold299 (.A(_01552_),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold300 (.A(\atari2600.ram[29][5] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold301 (.A(\atari2600.ram[21][2] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold302 (.A(\atari2600.ram[36][2] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold303 (.A(\atari2600.pia.swa_dir[6] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold304 (.A(\atari2600.ram[73][5] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold305 (.A(\atari2600.ram[105][2] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold306 (.A(\atari2600.ram[0][5] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold307 (.A(\atari2600.pia.swa_dir[0] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold308 (.A(\atari2600.ram[68][2] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold309 (.A(\atari2600.ram[33][2] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold310 (.A(\atari2600.ram[54][0] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold311 (.A(\atari2600.ram[37][6] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold312 (.A(\atari2600.ram[4][1] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold313 (.A(\atari2600.tia.cx[12] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold314 (.A(\atari2600.ram[69][2] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold315 (.A(\atari2600.ram[34][4] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold316 (.A(\atari2600.cpu.AXYS[2][2] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold317 (.A(\atari2600.ram[61][7] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold318 (.A(\atari2600.ram[50][7] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold319 (.A(\atari2600.cpu.cld ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold320 (.A(\atari2600.ram[57][1] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold321 (.A(\atari2600.ram[20][1] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold322 (.A(\atari2600.ram[70][0] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold323 (.A(\atari2600.ram[78][1] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold324 (.A(\atari2600.ram[21][4] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold325 (.A(\atari2600.tia.cx[6] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold326 (.A(\atari2600.ram[60][3] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold327 (.A(\atari2600.tia.audio_left_counter[4] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold328 (.A(_00995_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold329 (.A(\flash_rom.addr[9] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold330 (.A(_00976_),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold331 (.A(\atari2600.ram[100][5] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold332 (.A(\atari2600.ram[17][5] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold333 (.A(\atari2600.ram[56][6] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold334 (.A(\atari2600.ram[94][5] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold335 (.A(\atari2600.tia.audio_left_counter[7] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00998_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold337 (.A(\atari2600.ram[97][4] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold338 (.A(\atari2600.ram[0][4] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold339 (.A(\atari2600.ram[126][3] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold340 (.A(\atari2600.ram[64][0] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold341 (.A(\atari2600.ram[89][5] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold342 (.A(\atari2600.ram[33][0] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold343 (.A(\atari2600.ram[25][6] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold344 (.A(\atari2600.ram[113][1] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold345 (.A(\atari2600.ram[113][6] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold346 (.A(\atari2600.ram[113][7] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold347 (.A(\atari2600.ram[114][4] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold348 (.A(\atari2600.ram[109][3] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold349 (.A(\atari2600.ram[53][4] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold350 (.A(\atari2600.ram[16][4] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold351 (.A(\atari2600.ram[72][6] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold352 (.A(\atari2600.ram[8][6] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold353 (.A(\atari2600.ram[73][7] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold354 (.A(\atari2600.ram[66][6] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold355 (.A(\atari2600.ram[76][4] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold356 (.A(\atari2600.ram[124][3] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold357 (.A(\atari2600.ram[126][0] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold358 (.A(\atari2600.ram[52][4] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold359 (.A(\atari2600.ram[113][4] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold360 (.A(\atari2600.ram[94][2] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold361 (.A(\atari2600.pia.swa_dir[2] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold362 (.A(\atari2600.ram[102][3] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold363 (.A(\atari2600.ram[70][1] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold364 (.A(\atari2600.ram[58][4] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold365 (.A(\atari2600.ram[45][6] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold366 (.A(\atari2600.ram[29][6] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold367 (.A(\atari2600.ram[29][1] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold368 (.A(\atari2600.ram[97][5] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold369 (.A(\atari2600.ram[45][3] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold370 (.A(\atari2600.ram[57][4] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold371 (.A(\atari2600.ram[28][6] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold372 (.A(\atari2600.ram[53][7] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold373 (.A(\atari2600.ram[86][6] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold374 (.A(\atari2600.ram[6][1] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold375 (.A(\atari2600.ram[24][6] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold376 (.A(\atari2600.tia.cx[10] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold377 (.A(\atari2600.ram[52][0] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold378 (.A(\atari2600.ram[89][7] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold379 (.A(\atari2600.ram[72][0] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold380 (.A(\atari2600.ram[46][2] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold381 (.A(\atari2600.ram[13][3] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold382 (.A(\atari2600.ram[65][2] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold383 (.A(\atari2600.ram[96][3] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold384 (.A(\atari2600.ram[56][1] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold385 (.A(\atari2600.ram[94][4] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold386 (.A(\atari2600.ram[36][3] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold387 (.A(\atari2600.ram[64][3] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold388 (.A(\atari2600.ram[62][0] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold389 (.A(\atari2600.cpu.write_back ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold390 (.A(\atari2600.ram[114][7] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold391 (.A(\atari2600.ram[40][1] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold392 (.A(\atari2600.ram[109][5] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold393 (.A(\atari2600.ram[92][4] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold394 (.A(\atari2600.ram[42][3] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold395 (.A(\atari2600.ram[73][3] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold396 (.A(\atari2600.ram[40][2] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold397 (.A(\atari2600.ram[77][1] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold398 (.A(\atari2600.ram[76][5] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold399 (.A(\atari2600.ram[93][6] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold400 (.A(\atari2600.ram[61][1] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold401 (.A(\atari2600.ram[28][7] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold402 (.A(\atari2600.ram[81][7] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold403 (.A(\atari2600.ram[24][7] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold404 (.A(\atari2600.ram[106][7] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold405 (.A(\atari2600.ram[125][5] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold406 (.A(\atari2600.ram[73][2] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold407 (.A(\atari2600.cpu.AXYS[3][4] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00740_),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold409 (.A(spi_restart),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold410 (.A(\atari2600.cpu.AXYS[1][3] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold411 (.A(\atari2600.cpu.AXYS[3][7] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold412 (.A(\scanline[92][2] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold413 (.A(\atari2600.ram[100][2] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold414 (.A(\atari2600.ram[25][4] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold415 (.A(\atari2600.ram[13][6] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold416 (.A(\atari2600.ram[10][1] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold417 (.A(\atari2600.ram[22][6] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold418 (.A(\atari2600.ram[101][5] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold419 (.A(\atari2600.ram[70][7] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold420 (.A(\atari2600.ram[36][5] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold421 (.A(\atari2600.ram[98][1] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold422 (.A(\atari2600.ram[74][5] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold423 (.A(\atari2600.ram[102][2] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold424 (.A(\atari2600.ram[34][3] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold425 (.A(\atari2600.ram[98][6] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold426 (.A(\atari2600.ram[101][2] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold427 (.A(\atari2600.ram[126][1] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold428 (.A(\atari2600.ram[80][6] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold429 (.A(\external_rom_data[5] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold430 (.A(_01820_),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold431 (.A(\atari2600.tia.cx_clr ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold432 (.A(\atari2600.ram[108][1] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold433 (.A(\atari2600.ram[30][4] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold434 (.A(\atari2600.ram[34][2] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold435 (.A(\atari2600.ram[57][7] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold436 (.A(\atari2600.tia.audio_right_counter[4] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold437 (.A(_01011_),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold438 (.A(\atari2600.ram[104][5] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold439 (.A(\atari2600.ram[114][2] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold440 (.A(\atari2600.ram[60][7] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold441 (.A(\atari2600.ram[28][1] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold442 (.A(\atari2600.ram[94][6] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold443 (.A(\atari2600.ram[17][4] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold444 (.A(\atari2600.ram[105][1] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold445 (.A(\atari2600.ram[38][6] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold446 (.A(\atari2600.ram[98][3] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold447 (.A(\atari2600.ram[117][1] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold448 (.A(\atari2600.ram[116][2] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold449 (.A(\atari2600.ram[98][0] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold450 (.A(\atari2600.ram[40][4] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold451 (.A(\scanline[158][1] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold452 (.A(\atari2600.ram[17][7] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold453 (.A(\atari2600.ram[42][2] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold454 (.A(\atari2600.ram[61][4] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold455 (.A(\atari2600.ram[10][2] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold456 (.A(\atari2600.cpu.AXYS[2][7] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold457 (.A(\atari2600.ram[110][5] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold458 (.A(\atari2600.ram[88][7] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold459 (.A(\atari2600.ram[32][2] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold460 (.A(\atari2600.ram[14][6] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold461 (.A(\atari2600.ram[106][2] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold462 (.A(\atari2600.ram[18][2] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold463 (.A(\atari2600.ram[97][7] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold464 (.A(\atari2600.ram[74][6] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold465 (.A(\atari2600.ram[52][3] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold466 (.A(\atari2600.ram[120][6] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold467 (.A(\atari2600.ram[44][2] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold468 (.A(\atari2600.ram[32][5] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold469 (.A(\atari2600.ram[121][7] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold470 (.A(\atari2600.ram[90][2] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold471 (.A(\atari2600.tia.audio_left_counter[2] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold472 (.A(_00993_),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold473 (.A(\atari2600.ram[46][4] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold474 (.A(\atari2600.ram[16][3] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold475 (.A(\atari2600.ram[24][3] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold476 (.A(\atari2600.ram[85][6] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold477 (.A(\atari2600.ram[54][7] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold478 (.A(\atari2600.ram[85][5] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold479 (.A(\atari2600.ram[85][1] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold480 (.A(\atari2600.ram[112][7] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold481 (.A(\atari2600.ram[44][4] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold482 (.A(\atari2600.ram[2][4] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold483 (.A(\atari2600.ram[118][1] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold484 (.A(\atari2600.ram[116][0] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold485 (.A(\atari2600.ram[98][7] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold486 (.A(\atari2600.ram[121][4] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold487 (.A(\scanline[29][0] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold488 (.A(\atari2600.ram[46][7] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold489 (.A(\atari2600.ram[42][5] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold490 (.A(\scanline[105][0] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold491 (.A(\atari2600.ram[101][4] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold492 (.A(\atari2600.ram[122][3] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold493 (.A(\atari2600.ram[97][1] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold494 (.A(\atari2600.ram[106][4] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold495 (.A(\gamepad_pmod.decoder.data_reg[11] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold496 (.A(_01563_),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold497 (.A(\atari2600.ram[90][4] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold498 (.A(\atari2600.ram[3][6] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold499 (.A(\scanline[150][1] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold500 (.A(\atari2600.ram[44][6] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold501 (.A(\atari2600.ram[106][3] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold502 (.A(\scanline[105][2] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold503 (.A(\atari2600.ram[77][2] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold504 (.A(\atari2600.ram[106][6] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold505 (.A(\atari2600.ram[108][2] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold506 (.A(\atari2600.ram[62][5] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold507 (.A(\atari2600.ram[114][1] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold508 (.A(\atari2600.ram[22][3] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold509 (.A(\atari2600.ram[105][3] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold510 (.A(\atari2600.cpu.AXYS[1][4] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold511 (.A(_01600_),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold512 (.A(\atari2600.tia.p0_copies[1] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold513 (.A(\atari2600.ram[10][0] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold514 (.A(\scanline[158][4] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold515 (.A(\scanline[29][3] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold516 (.A(\scanline[91][1] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold517 (.A(\atari2600.ram[22][5] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold518 (.A(\atari2600.ram[20][5] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold519 (.A(\atari2600.ram[58][6] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold520 (.A(\scanline[125][0] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold521 (.A(\scanline[46][0] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold522 (.A(\atari2600.ram[81][2] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold523 (.A(\atari2600.ram[84][7] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold524 (.A(\atari2600.ram[4][4] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold525 (.A(\atari2600.ram[52][7] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold526 (.A(\atari2600.ram[69][4] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold527 (.A(\scanline[77][2] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold528 (.A(\scanline[45][3] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold529 (.A(_00070_),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold530 (.A(_00051_),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold531 (.A(\scanline[117][2] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold532 (.A(\atari2600.ram[28][3] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold533 (.A(\atari2600.ram[117][4] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold534 (.A(\scanline[54][5] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold535 (.A(\atari2600.ram[122][5] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold536 (.A(\atari2600.ram[44][3] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold537 (.A(\scanline[53][4] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold538 (.A(\atari2600.cpu.AXYS[2][5] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold539 (.A(\atari2600.ram[89][3] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold540 (.A(\scanline[62][6] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold541 (.A(\scanline[78][2] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold542 (.A(\atari2600.cpu.src_reg[0] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold543 (.A(\scanline[94][6] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold544 (.A(\atari2600.ram[52][2] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold545 (.A(\scanline[114][5] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold546 (.A(\atari2600.ram[121][2] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold547 (.A(\atari2600.ram[85][7] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold548 (.A(\atari2600.ram[53][5] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold549 (.A(\scanline[29][1] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold550 (.A(\atari2600.ram[126][4] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold551 (.A(\scanline[117][3] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold552 (.A(\scanline[110][6] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold553 (.A(\atari2600.cpu.AXYS[3][5] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold554 (.A(\scanline[153][5] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold555 (.A(\atari2600.ram[42][6] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold556 (.A(\scanline[127][3] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold557 (.A(\scanline[109][0] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold558 (.A(\atari2600.ram[66][0] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold559 (.A(\atari2600.ram[118][6] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold560 (.A(\atari2600.ram[60][4] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold561 (.A(\external_rom_data[4] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold562 (.A(_01819_),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold563 (.A(\scanline[58][2] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold564 (.A(\atari2600.ram[49][7] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold565 (.A(\scanline[89][6] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold566 (.A(\atari2600.ram[106][5] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold567 (.A(\scanline[77][5] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold568 (.A(\atari2600.ram[69][6] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold569 (.A(\atari2600.ram[10][5] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold570 (.A(\scanline[142][4] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold571 (.A(\scanline[106][1] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold572 (.A(\scanline[51][4] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold573 (.A(\scanline[62][1] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold574 (.A(\scanline[142][3] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold575 (.A(\scanline[107][1] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold576 (.A(\scanline[151][6] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold577 (.A(\scanline[110][4] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold578 (.A(\atari2600.ram[69][5] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold579 (.A(\scanline[94][3] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold580 (.A(\atari2600.ram[90][3] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold581 (.A(\scanline[156][5] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold582 (.A(\scanline[122][2] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold583 (.A(\atari2600.ram[18][7] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold584 (.A(\scanline[102][4] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold585 (.A(\scanline[61][3] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold586 (.A(\scanline[15][6] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold587 (.A(\atari2600.ram[56][0] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold588 (.A(\scanline[108][5] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold589 (.A(\scanline[13][2] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold590 (.A(\scanline[103][4] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold591 (.A(\scanline[60][4] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold592 (.A(\scanline[91][5] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold593 (.A(\scanline[31][6] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold594 (.A(\atari2600.cpu.ABL[7] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold595 (.A(\atari2600.ram[41][6] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold596 (.A(\atari2600.ram[98][4] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold597 (.A(\scanline[54][3] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold598 (.A(\atari2600.ram[10][4] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold599 (.A(\atari2600.ram[32][1] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold600 (.A(\atari2600.ram[80][1] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold601 (.A(\atari2600.ram[72][1] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold602 (.A(\atari2600.ram[70][4] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold603 (.A(\atari2600.ram[82][7] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold604 (.A(\atari2600.ram[116][1] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold605 (.A(\atari2600.ram[24][0] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold606 (.A(\atari2600.tia.old_grp0[6] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold607 (.A(_01098_),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold608 (.A(\atari2600.ram[114][3] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold609 (.A(\atari2600.tia.old_grp0[7] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01099_),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold611 (.A(\atari2600.ram[25][7] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold612 (.A(\scanline[105][4] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold613 (.A(\atari2600.ram[100][3] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold614 (.A(\scanline[123][4] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold615 (.A(\scanline[13][4] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold616 (.A(\atari2600.ram[33][1] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold617 (.A(\atari2600.ram[18][4] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold618 (.A(\atari2600.ram[52][5] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold619 (.A(\atari2600.cpu.sei ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold620 (.A(_01359_),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold621 (.A(\scanline[105][6] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold622 (.A(\atari2600.ram[84][0] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold623 (.A(\scanline[108][0] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold624 (.A(\scanline[111][6] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold625 (.A(\atari2600.ram[38][1] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold626 (.A(\atari2600.ram[26][2] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold627 (.A(\atari2600.ram[38][5] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold628 (.A(\atari2600.ram[20][4] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold629 (.A(\scanline[53][1] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold630 (.A(\atari2600.ram[70][3] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold631 (.A(\atari2600.ram[118][0] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold632 (.A(\scanline[31][1] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold633 (.A(\scanline[46][6] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold634 (.A(\atari2600.ram[44][0] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold635 (.A(\atari2600.ram[124][1] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold636 (.A(\scanline[121][0] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold637 (.A(\atari2600.ram[14][3] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold638 (.A(\atari2600.ram[85][4] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold639 (.A(\scanline[61][5] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold640 (.A(\atari2600.ram[96][2] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold641 (.A(\scanline[31][0] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold642 (.A(\atari2600.ram[9][0] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold643 (.A(\scanline[78][3] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold644 (.A(\atari2600.ram[92][6] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold645 (.A(\atari2600.ram[88][1] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold646 (.A(\atari2600.ram[26][3] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold647 (.A(\atari2600.ram[110][4] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold648 (.A(\atari2600.ram[102][1] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold649 (.A(\scanline[51][6] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold650 (.A(\scanline[79][5] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold651 (.A(\scanline[125][3] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold652 (.A(\scanline[107][3] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold653 (.A(\scanline[141][4] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold654 (.A(\scanline[115][3] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold655 (.A(\atari2600.ram[96][5] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold656 (.A(\atari2600.ram[86][2] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold657 (.A(\scanline[141][5] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold658 (.A(\atari2600.ram[64][1] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold659 (.A(\atari2600.ram[13][4] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold660 (.A(\scanline[124][3] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold661 (.A(\atari2600.ram[88][5] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold662 (.A(\atari2600.ram[94][3] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold663 (.A(\scanline[122][3] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold664 (.A(\scanline[110][3] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold665 (.A(\scanline[57][3] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold666 (.A(\atari2600.ram[56][4] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold667 (.A(\scanline[92][3] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold668 (.A(\scanline[30][5] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold669 (.A(\scanline[109][4] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold670 (.A(\atari2600.ram[56][7] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold671 (.A(\atari2600.ram[93][1] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold672 (.A(\scanline[58][4] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold673 (.A(\atari2600.ram[33][5] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold674 (.A(\scanline[60][0] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold675 (.A(\atari2600.ram[12][3] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold676 (.A(\scanline[109][2] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold677 (.A(\atari2600.ram[36][0] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold678 (.A(\atari2600.tia.audio_left_counter[12] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold679 (.A(_01003_),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold680 (.A(\atari2600.ram[28][2] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold681 (.A(\atari2600.ram[65][4] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold682 (.A(\scanline[90][1] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold683 (.A(\atari2600.ram[88][2] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold684 (.A(\atari2600.ram[108][7] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold685 (.A(\scanline[54][6] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold686 (.A(\atari2600.pia.interval[10] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold687 (.A(\scanline[63][1] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold688 (.A(\atari2600.ram[116][7] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold689 (.A(\scanline[156][1] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold690 (.A(\atari2600.pia.time_counter[22] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold691 (.A(_05461_),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold692 (.A(_00896_),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold693 (.A(\atari2600.ram[50][1] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold694 (.A(\scanline[55][2] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold695 (.A(\scanline[62][5] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold696 (.A(\scanline[79][4] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold697 (.A(\scanline[125][5] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold698 (.A(\scanline[78][4] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold699 (.A(\atari2600.ram[104][4] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold700 (.A(\scanline[154][2] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold701 (.A(\scanline[59][6] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold702 (.A(\atari2600.cpu.AXYS[1][5] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold703 (.A(\atari2600.ram[69][7] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold704 (.A(\scanline[121][6] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold705 (.A(\scanline[87][6] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold706 (.A(\scanline[93][3] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold707 (.A(\atari2600.ram[84][5] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold708 (.A(\scanline[45][5] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold709 (.A(\atari2600.ram[86][3] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold710 (.A(\atari2600.ram[17][3] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold711 (.A(\atari2600.cpu.AXYS[2][3] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold712 (.A(\atari2600.tia.old_grp0[0] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold713 (.A(_01092_),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold714 (.A(\atari2600.ram[22][4] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold715 (.A(\atari2600.cpu.PC[2] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold716 (.A(_01412_),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold717 (.A(\atari2600.ram[49][1] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold718 (.A(\atari2600.ram[78][6] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold719 (.A(\scanline[14][3] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold720 (.A(\atari2600.ram[3][0] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold721 (.A(\scanline[63][5] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold722 (.A(\atari2600.ram[81][5] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold723 (.A(\atari2600.ram[21][7] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold724 (.A(\atari2600.ram[106][0] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold725 (.A(\atari2600.cpu.AXYS[2][6] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold726 (.A(\atari2600.tia.cx[4] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold727 (.A(\atari2600.ram[14][1] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold728 (.A(\atari2600.ram[10][7] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold729 (.A(\atari2600.tia.old_grp0[2] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold730 (.A(_01094_),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold731 (.A(\scanline[45][2] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold732 (.A(\scanline[108][3] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold733 (.A(\atari2600.ram[50][5] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold734 (.A(\scanline[91][2] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold735 (.A(\atari2600.ram[45][5] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold736 (.A(\atari2600.ram[105][7] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold737 (.A(\atari2600.ram[2][5] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold738 (.A(\atari2600.tia.old_grp0[4] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold739 (.A(_01096_),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold740 (.A(\atari2600.ram[82][5] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold741 (.A(\scanline[103][3] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold742 (.A(\atari2600.ram[25][5] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold743 (.A(\scanline[94][2] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold744 (.A(\atari2600.ram[5][3] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold745 (.A(\atari2600.cpu.AXYS[1][0] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold746 (.A(\scanline[106][6] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold747 (.A(\atari2600.ram[96][7] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold748 (.A(\atari2600.ram[3][2] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold749 (.A(\atari2600.ram[4][5] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold750 (.A(\scanline[85][5] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold751 (.A(\scanline[105][1] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold752 (.A(\scanline[108][1] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold753 (.A(\scanline[14][0] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold754 (.A(\scanline[103][2] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold755 (.A(\scanline[158][6] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold756 (.A(\atari2600.ram[98][2] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold757 (.A(\scanline[106][0] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold758 (.A(\scanline[57][6] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold759 (.A(\scanline[113][4] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold760 (.A(\scanline[60][1] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold761 (.A(\atari2600.ram[62][6] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold762 (.A(\atari2600.ram[50][6] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold763 (.A(\scanline[93][4] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold764 (.A(\scanline[85][4] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold765 (.A(\atari2600.ram[70][6] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold766 (.A(\atari2600.ram[50][0] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold767 (.A(\scanline[124][4] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold768 (.A(\atari2600.ram[12][7] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold769 (.A(\atari2600.ram[37][1] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold770 (.A(\scanline[92][4] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold771 (.A(\scanline[92][6] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold772 (.A(\scanline[127][1] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold773 (.A(\scanline[93][0] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold774 (.A(\scanline[107][2] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold775 (.A(\atari2600.ram[0][3] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold776 (.A(\atari2600.ram[12][0] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold777 (.A(\scanline[89][5] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold778 (.A(\atari2600.cpu.AXYS[3][6] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold779 (.A(\atari2600.ram[5][5] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold780 (.A(\scanline[126][4] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold781 (.A(\atari2600.ram[90][7] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold782 (.A(\atari2600.pia.swa_dir[5] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold783 (.A(\scanline[47][2] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold784 (.A(\atari2600.ram[116][3] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold785 (.A(\scanline[89][1] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold786 (.A(\atari2600.ram[17][2] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold787 (.A(\atari2600.ram[73][1] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold788 (.A(\atari2600.ram[117][0] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold789 (.A(\atari2600.cpu.AXYS[2][1] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold790 (.A(\atari2600.ram[37][5] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold791 (.A(\atari2600.ram[37][0] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold792 (.A(\atari2600.ram[82][3] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold793 (.A(\atari2600.ram[45][1] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold794 (.A(\scanline[122][1] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold795 (.A(\atari2600.ram[61][6] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold796 (.A(\atari2600.ram[30][0] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold797 (.A(\atari2600.ram[41][1] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold798 (.A(\scanline[149][4] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold799 (.A(\atari2600.pia.instat[1] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold800 (.A(_00865_),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold801 (.A(\atari2600.ram[44][5] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold802 (.A(\scanline[95][0] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold803 (.A(\scanline[58][1] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold804 (.A(\scanline[14][6] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold805 (.A(\atari2600.ram[9][2] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold806 (.A(\atari2600.ram[80][7] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold807 (.A(\scanline[61][0] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold808 (.A(\scanline[13][3] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold809 (.A(\scanline[101][1] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold810 (.A(\atari2600.ram[8][3] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold811 (.A(\atari2600.ram[92][7] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold812 (.A(\scanline[79][2] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold813 (.A(\scanline[117][1] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold814 (.A(\atari2600.ram[86][7] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold815 (.A(\scanline[63][0] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold816 (.A(\scanline[14][4] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold817 (.A(\atari2600.ram[9][4] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold818 (.A(\atari2600.ram[82][4] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold819 (.A(\flash_rom.addr[23] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold820 (.A(_00982_),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold821 (.A(\scanline[122][0] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold822 (.A(\scanline[95][6] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold823 (.A(\atari2600.ram[113][3] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold824 (.A(\scanline[110][0] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold825 (.A(\atari2600.ram[30][3] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold826 (.A(\atari2600.ram[25][2] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold827 (.A(\atari2600.ram[66][3] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold828 (.A(\scanline[90][2] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold829 (.A(\scanline[126][5] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold830 (.A(\atari2600.ram[109][1] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold831 (.A(\atari2600.ram[58][2] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold832 (.A(\atari2600.ram[117][5] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold833 (.A(\scanline[118][1] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold834 (.A(\atari2600.ram[58][7] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold835 (.A(\atari2600.ram[13][2] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold836 (.A(\scanline[114][2] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold837 (.A(\scanline[94][1] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold838 (.A(\scanline[117][4] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold839 (.A(\scanline[78][0] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold840 (.A(\scanline[127][6] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold841 (.A(\scanline[151][4] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold842 (.A(\atari2600.ram[94][1] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold843 (.A(\atari2600.ram[13][7] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold844 (.A(\atari2600.ram[77][5] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold845 (.A(\scanline[101][5] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold846 (.A(\atari2600.ram[109][6] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold847 (.A(\scanline[124][2] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold848 (.A(\atari2600.ram[5][2] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold849 (.A(\atari2600.ram[1][5] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold850 (.A(\atari2600.tia.audio_left_counter[10] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold851 (.A(_01001_),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold852 (.A(\atari2600.ram[125][1] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold853 (.A(\scanline[123][6] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold854 (.A(\atari2600.ram[104][2] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold855 (.A(\atari2600.ram[61][5] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold856 (.A(\scanline[57][1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold857 (.A(\atari2600.ram[30][6] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold858 (.A(\scanline[123][3] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold859 (.A(\gamepad_pmod.decoder.data_reg[4] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold860 (.A(_01556_),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold861 (.A(\atari2600.ram[120][7] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold862 (.A(\scanline[108][6] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold863 (.A(\scanline[58][3] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold864 (.A(\atari2600.ram[120][5] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold865 (.A(\atari2600.ram[6][2] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold866 (.A(\scanline[111][5] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold867 (.A(\atari2600.ram[53][6] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold868 (.A(\scanline[55][0] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold869 (.A(\scanline[77][1] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold870 (.A(\atari2600.ram[26][0] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold871 (.A(\atari2600.ram[5][6] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold872 (.A(\atari2600.tia.audio_right_counter[6] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold873 (.A(_01013_),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold874 (.A(\scanline[123][0] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold875 (.A(\scanline[30][0] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold876 (.A(\scanline[62][3] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold877 (.A(\scanline[13][5] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold878 (.A(\scanline[153][0] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold879 (.A(\scanline[157][2] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold880 (.A(\atari2600.ram[3][5] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold881 (.A(\scanline[115][2] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold882 (.A(\scanline[89][0] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold883 (.A(\atari2600.ram[29][3] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold884 (.A(\atari2600.ram[84][1] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold885 (.A(\atari2600.tia.old_grp0[3] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold886 (.A(_01095_),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold887 (.A(\atari2600.ram[45][7] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold888 (.A(\scanline[126][3] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold889 (.A(\atari2600.ram[3][7] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold890 (.A(\scanline[101][6] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold891 (.A(\scanline[121][1] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold892 (.A(\atari2600.ram[21][1] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold893 (.A(\scanline[45][6] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold894 (.A(\atari2600.ram[68][4] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold895 (.A(\scanline[90][0] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold896 (.A(\scanline[89][3] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold897 (.A(\scanline[105][5] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold898 (.A(\scanline[59][3] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold899 (.A(\atari2600.ram[46][3] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold900 (.A(\atari2600.cpu.AXYS[1][1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold901 (.A(\atari2600.tia.audio_left_counter[8] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold902 (.A(_00999_),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold903 (.A(\scanline[58][6] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold904 (.A(\scanline[14][2] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold905 (.A(\scanline[108][4] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold906 (.A(\scanline[78][5] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold907 (.A(\atari2600.ram[73][6] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold908 (.A(\atari2600.ram[52][1] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold909 (.A(\scanline[31][4] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold910 (.A(\scanline[92][1] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold911 (.A(\scanline[77][0] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold912 (.A(\scanline[106][4] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold913 (.A(\scanline[150][3] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold914 (.A(\scanline[142][0] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold915 (.A(\atari2600.ram[77][4] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold916 (.A(\atari2600.tia.audio_right_counter[10] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold917 (.A(_01017_),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold918 (.A(\atari2600.ram[28][4] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold919 (.A(\scanline[121][3] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold920 (.A(\scanline[30][1] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold921 (.A(\scanline[79][3] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold922 (.A(\scanline[103][6] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold923 (.A(\scanline[85][3] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold924 (.A(\atari2600.ram[88][6] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold925 (.A(\scanline[111][4] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold926 (.A(\scanline[63][4] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold927 (.A(\atari2600.ram[73][4] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold928 (.A(\scanline[154][5] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold929 (.A(\atari2600.ram[124][6] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold930 (.A(\scanline[154][4] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold931 (.A(\scanline[125][2] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold932 (.A(\scanline[155][0] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold933 (.A(\scanline[159][3] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold934 (.A(\atari2600.ram[106][1] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold935 (.A(\atari2600.ram[117][7] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold936 (.A(\scanline[115][6] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold937 (.A(\atari2600.ram[6][3] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold938 (.A(\scanline[107][6] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold939 (.A(\scanline[151][5] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold940 (.A(\scanline[87][4] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold941 (.A(\atari2600.ram[78][0] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold942 (.A(\atari2600.ram[37][7] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold943 (.A(\atari2600.ram[30][2] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold944 (.A(\atari2600.cpu.AXYS[3][3] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold945 (.A(\atari2600.ram[112][3] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold946 (.A(\atari2600.ram[74][7] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold947 (.A(\scanline[114][1] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold948 (.A(\scanline[47][5] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold949 (.A(\scanline[79][1] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold950 (.A(\scanline[47][1] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold951 (.A(\atari2600.ram[46][5] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold952 (.A(\atari2600.ram[97][2] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold953 (.A(\atari2600.ram[20][6] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold954 (.A(\scanline[111][3] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold955 (.A(\atari2600.ram[121][3] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold956 (.A(\atari2600.ram[68][5] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold957 (.A(\atari2600.ram[76][3] ),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold958 (.A(\atari2600.ram[60][6] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold959 (.A(\scanline[141][3] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold960 (.A(\atari2600.ram[60][2] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold961 (.A(\atari2600.pia.swb_dir[5] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold962 (.A(\scanline[115][0] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold963 (.A(\scanline[121][5] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold964 (.A(\atari2600.ram[122][4] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold965 (.A(\scanline[125][1] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold966 (.A(\scanline[102][6] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold967 (.A(\atari2600.cpu.AXYS[2][4] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold968 (.A(_01592_),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold969 (.A(\atari2600.ram[32][7] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold970 (.A(\scanline[60][6] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold971 (.A(\scanline[103][1] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold972 (.A(\atari2600.ram[121][0] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold973 (.A(\atari2600.ram[126][2] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold974 (.A(\scanline[113][5] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold975 (.A(\atari2600.ram[85][0] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold976 (.A(\atari2600.ram[109][0] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold977 (.A(\atari2600.ram[80][5] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold978 (.A(\atari2600.ram[125][0] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold979 (.A(\atari2600.ram[76][1] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold980 (.A(\scanline[108][2] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold981 (.A(\atari2600.ram[93][7] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold982 (.A(\scanline[51][2] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold983 (.A(\atari2600.ram[93][3] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold984 (.A(\scanline[61][2] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold985 (.A(\atari2600.ram[62][4] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold986 (.A(\scanline[90][4] ),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold987 (.A(\scanline[109][6] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold988 (.A(\scanline[13][1] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold989 (.A(\scanline[55][3] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold990 (.A(\scanline[63][3] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold991 (.A(\atari2600.tia.old_grp0[1] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold992 (.A(_01093_),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold993 (.A(\atari2600.ram[113][2] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold994 (.A(\atari2600.ram[53][0] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold995 (.A(\atari2600.ram[21][3] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold996 (.A(\scanline[111][1] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold997 (.A(\scanline[125][6] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold998 (.A(\scanline[55][1] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold999 (.A(\scanline[111][2] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\scanline[102][1] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\scanline[93][2] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\atari2600.ram[25][1] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\scanline[47][3] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\scanline[143][6] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\scanline[46][3] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\scanline[57][4] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\scanline[154][0] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\scanline[86][5] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\scanline[126][0] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\scanline[77][3] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\atari2600.ram[64][6] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\flash_rom.addr[21] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_00980_),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\atari2600.ram[100][1] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\scanline[154][3] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\atari2600.ram[88][4] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\scanline[127][2] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\scanline[47][0] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\scanline[61][4] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\atari2600.ram[118][5] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\scanline[151][0] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\atari2600.ram[22][1] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\scanline[157][6] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\atari2600.ram[2][2] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\atari2600.ram[22][0] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\scanline[92][5] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\scanline[109][5] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\scanline[109][3] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\atari2600.ram[66][2] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\atari2600.ram[0][6] ),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\atari2600.ram[68][0] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\atari2600.ram[6][5] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\scanline[123][1] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\atari2600.ram[1][1] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\scanline[95][2] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\atari2600.ram[58][1] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\atari2600.cpu.AXYS[1][7] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\atari2600.ram[84][3] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\atari2600.ram[82][2] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\scanline[142][5] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\scanline[93][5] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\scanline[107][4] ),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\scanline[119][4] ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\atari2600.ram[105][6] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\atari2600.ram[104][3] ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\atari2600.ram[56][3] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\scanline[113][2] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\scanline[13][6] ),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\atari2600.ram[77][7] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\scanline[124][6] ),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\atari2600.ram[20][2] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\atari2600.ram[101][3] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\atari2600.ram[17][6] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\scanline[59][1] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\atari2600.ram[5][0] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\scanline[149][2] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\scanline[61][1] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\scanline[157][4] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\scanline[15][5] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\scanline[124][5] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\atari2600.ram[54][3] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\atari2600.ram[50][2] ),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\atari2600.ram[117][6] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\scanline[159][2] ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\atari2600.ram[101][1] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\scanline[149][3] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\scanline[142][1] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\scanline[115][1] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\atari2600.ram[14][2] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\scanline[106][3] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\scanline[87][5] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\scanline[142][2] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\scanline[53][2] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\scanline[60][5] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\atari2600.ram[125][6] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\scanline[119][6] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\scanline[155][6] ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\scanline[86][1] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\scanline[47][6] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\scanline[117][6] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\scanline[92][0] ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\atari2600.ram[58][5] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\atari2600.ram[124][7] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\scanline[93][6] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\atari2600.ram[78][5] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\scanline[78][6] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\atari2600.ram[72][3] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\atari2600.ram[109][7] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\scanline[113][3] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\scanline[124][1] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\scanline[85][1] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\scanline[46][1] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\scanline[113][0] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\scanline[14][1] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\scanline[118][6] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\scanline[157][0] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\scanline[153][6] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\scanline[105][3] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\scanline[107][0] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\atari2600.ram[14][7] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\scanline[123][2] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\atari2600.ram[65][3] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\atari2600.ram[33][7] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\atari2600.ram[57][0] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\atari2600.ram[42][1] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\scanline[127][4] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\scanline[143][2] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\scanline[62][0] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\scanline[55][5] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\scanline[15][0] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\atari2600.ram[65][0] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\scanline[153][2] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\scanline[61][6] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\atari2600.ram[4][3] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\scanline[107][5] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\scanline[90][6] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\scanline[78][1] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\scanline[122][6] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\scanline[121][4] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\scanline[95][4] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\atari2600.ram[40][6] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\atari2600.ram[38][7] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\scanline[86][6] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\scanline[94][0] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\scanline[53][5] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\scanline[106][2] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\scanline[118][4] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\scanline[93][1] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\scanline[125][4] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\scanline[103][0] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\scanline[57][2] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\atari2600.ram[110][2] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\atari2600.ram[16][6] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\atari2600.ram[86][0] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\atari2600.ram[113][0] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\scanline[29][6] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\atari2600.ram[110][3] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\atari2600.ram[62][2] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\scanline[151][2] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\scanline[51][0] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\scanline[53][6] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\atari2600.ram[90][0] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\atari2600.ram[112][4] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\atari2600.ram[26][7] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\atari2600.ram[92][1] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\atari2600.ram[52][6] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\scanline[94][4] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\atari2600.ram[26][1] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\scanline[79][0] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\scanline[90][3] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\atari2600.ram[8][2] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\scanline[59][4] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\scanline[124][0] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\atari2600.ram[46][1] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\scanline[57][0] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\atari2600.ram[102][6] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\scanline[109][1] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\scanline[150][6] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\scanline[111][0] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\scanline[89][4] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\scanline[30][4] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\atari2600.pia.swa_dir[4] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\atari2600.ram[48][3] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\atari2600.ram[37][3] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\scanline[94][5] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\scanline[114][3] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\scanline[54][0] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\atari2600.cpu.AXYS[3][0] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\scanline[51][3] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\scanline[77][4] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\atari2600.ram[48][4] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\scanline[106][5] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\scanline[118][3] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\atari2600.ram[62][3] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\scanline[143][5] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\gamepad_pmod.decoder.data_reg[6] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1177 (.A(_01558_),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\atari2600.tia.cx[5] ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\scanline[142][6] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\scanline[14][5] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\atari2600.ram[64][2] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\atari2600.ram[61][2] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\atari2600.ram[90][5] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\scanline[154][6] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\scanline[159][5] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\scanline[143][1] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\atari2600.ram[84][2] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\scanline[46][4] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\atari2600.ram[61][0] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\scanline[153][4] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\scanline[126][6] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\atari2600.ram[102][0] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\scanline[87][1] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\atari2600.ram[98][5] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\atari2600.ram[124][5] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\scanline[158][2] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\scanline[121][2] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\scanline[110][2] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\scanline[157][3] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\scanline[110][1] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\scanline[150][2] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\scanline[15][3] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\scanline[118][2] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\atari2600.ram[2][1] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\scanline[95][3] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\atari2600.ram[76][0] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\scanline[86][2] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\atari2600.ram[72][5] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\scanline[151][1] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\scanline[158][0] ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\scanline[63][6] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\scanline[156][4] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\scanline[101][3] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\atari2600.ram[34][1] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\atari2600.tia.cx[11] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\scanline[101][4] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\scanline[103][5] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\scanline[45][4] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\atari2600.ram[54][1] ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\scanline[51][1] ),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\scanline[102][0] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\scanline[102][2] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\scanline[46][5] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\atari2600.pia.time_counter[5] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1225 (.A(_05418_),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\scanline[60][2] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\atari2600.ram[6][7] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_00132_),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_01812_),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\scanline[91][3] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\atari2600.ram[97][0] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\scanline[115][5] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\scanline[158][5] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\atari2600.ram[60][5] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\scanline[87][0] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\scanline[31][2] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\atari2600.ram[120][1] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\external_rom_data[6] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_01821_),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\scanline[101][0] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\atari2600.ram[65][1] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\scanline[86][0] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\scanline[155][3] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\scanline[155][4] ),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\scanline[151][3] ),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\atari2600.ram[90][1] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\scanline[59][0] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\atari2600.ram[66][7] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\atari2600.cpu.N ),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\scanline[15][2] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\scanline[55][6] ),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\scanline[126][1] ),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\scanline[57][5] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\atari2600.ram[110][0] ),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\scanline[114][4] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\scanline[114][0] ),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\atari2600.ram[74][1] ),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\atari2600.ram[22][7] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\atari2600.ram[122][0] ),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\atari2600.ram[9][7] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\atari2600.ram[114][5] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\atari2600.tia.old_grp0[5] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1263 (.A(_01097_),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\atari2600.pia.swb_dir[2] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\atari2600.ram[26][5] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\scanline[55][4] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\scanline[143][4] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\atari2600.ram[113][5] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\atari2600.ram[38][0] ),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\atari2600.ram[86][1] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\atari2600.ram[49][2] ),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\atari2600.ram[48][2] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\atari2600.ram[66][1] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\scanline[95][1] ),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\scanline[102][3] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\scanline[141][6] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\scanline[86][3] ),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\scanline[115][4] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\scanline[91][4] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\scanline[153][3] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\atari2600.ram[125][4] ),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\atari2600.ram[126][5] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\atari2600.tia.audio_right_counter[2] ),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_01009_),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\atari2600.ram[6][6] ),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\scanline[150][4] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\atari2600.ram[74][0] ),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\atari2600.ram[86][4] ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\atari2600.ram[114][0] ),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\atari2600.ram[42][4] ),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\atari2600.ram[100][0] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\atari2600.ram[78][7] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\atari2600.ram[84][4] ),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\scanline[118][0] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\scanline[113][6] ),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\scanline[13][0] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\atari2600.ram[68][7] ),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\scanline[46][2] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\scanline[60][3] ),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\atari2600.ram[54][4] ),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\atari2600.cpu.AXYS[1][2] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\scanline[156][2] ),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\atari2600.ram[64][5] ),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\scanline[91][6] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\scanline[90][5] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\scanline[119][2] ),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\atari2600.ram[18][6] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\scanline[127][0] ),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\atari2600.ram[26][4] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\atari2600.ram[48][0] ),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\atari2600.ram[110][7] ),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\scanline[114][6] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\scanline[87][3] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\scanline[126][2] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\atari2600.ram[6][0] ),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\scanline[53][0] ),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\frame_counter[2] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1318 (.A(_00348_),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\scanline[29][4] ),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\scanline[31][5] ),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\scanline[85][6] ),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\atari2600.pia.swa_dir[3] ),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\atari2600.ram[45][2] ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\atari2600.ram[78][2] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\atari2600.ram[112][5] ),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\atari2600.ram[104][0] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\atari2600.ram[100][7] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\atari2600.ram[38][2] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\atari2600.ram[86][5] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\scanline[29][5] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\scanline[53][3] ),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\atari2600.ram[34][0] ),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\scanline[143][3] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\scanline[159][1] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\scanline[119][5] ),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\atari2600.ram[10][6] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\scanline[158][3] ),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\scanline[159][6] ),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\scanline[86][4] ),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\scanline[63][2] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\scanline[45][0] ),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\scanline[123][5] ),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\scanline[30][2] ),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\scanline[15][4] ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\scanline[156][0] ),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\atari2600.ram[74][2] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\scanline[79][6] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\g_pwm_even[1] ),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_04607_),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_00338_),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\atari2600.ram[92][3] ),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\atari2600.ram[122][1] ),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\scanline[155][5] ),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\scanline[156][3] ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\atari2600.ram[68][6] ),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\atari2600.ram[92][2] ),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\atari2600.ram[118][3] ),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\atari2600.ram[14][5] ),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\scanline[122][5] ),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\atari2600.ram[74][3] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\atari2600.ram[102][5] ),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\atari2600.ram[78][4] ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\atari2600.ram[49][4] ),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\scanline[119][0] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\atari2600.ram[36][7] ),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\atari2600.tia.p1_copies[2] ),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\atari2600.ram[110][1] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\atari2600.ram[32][0] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\atari2600.ram[74][4] ),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\scanline[149][1] ),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\atari2600.ram[30][5] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\atari2600.ram[60][0] ),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\atari2600.ram[4][6] ),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\atari2600.ram[122][7] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\atari2600.ram[3][3] ),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\atari2600.tia.m1_w[3] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\atari2600.ram[33][6] ),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\atari2600.ram[32][6] ),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\atari2600.cpu.AXYS[3][1] ),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\scanline[113][1] ),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\scanline[154][1] ),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\atari2600.ram[2][3] ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\atari2600.ram[126][6] ),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\scanline[59][5] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\atari2600.ram[124][2] ),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\atari2600.ram[54][6] ),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\scanline[54][4] ),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\atari2600.ram[78][3] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\scanline[59][2] ),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\atari2600.ram[50][3] ),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\atari2600.ram[18][3] ),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\atari2600.ram[121][5] ),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\scanline[101][2] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\atari2600.cpu.clc ),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\atari2600.ram[18][1] ),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\atari2600.ram[104][7] ),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\atari2600.pia.time_counter[17] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1398 (.A(_05450_),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\scanline[62][4] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\scanline[30][6] ),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\atari2600.ram[117][3] ),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\atari2600.ram[89][0] ),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\atari2600.ram[26][6] ),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\scanline[85][2] ),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\atari2600.ram[22][2] ),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\scanline[89][2] ),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\scanline[62][2] ),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\atari2600.ram[1][7] ),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\rom_last_read_addr[5] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_00269_),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\atari2600.ram[48][6] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\atari2600.ram[25][3] ),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\atari2600.ram[5][7] ),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\atari2600.tia.dat_o[7] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\atari2600.cpu.AXYS[1][6] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\scanline[141][2] ),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\scanline[122][4] ),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\atari2600.ram[13][0] ),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\atari2600.tia.diag[101] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1420 (.A(_00920_),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\scanline[87][2] ),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\scanline[85][0] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\gamepad_pmod.decoder.data_reg[7] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_01559_),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\atari2600.ram[90][6] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\atari2600.tia.m1_w[0] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\scanline[58][5] ),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\scanline[117][5] ),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\scanline[141][1] ),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\scanline[47][4] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\atari2600.ram[1][6] ),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\scanline[153][1] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\atari2600.ram[97][6] ),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\scanline[149][6] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\atari2600.ram[72][7] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\scanline[110][5] ),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\atari2600.ram[54][2] ),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\scanline[100][5] ),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\atari2600.ram[14][0] ),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\atari2600.ram[66][4] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\atari2600.ram[54][5] ),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\scanline[91][0] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\rom_last_read_addr[10] ),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1444 (.A(_00274_),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\scanline[149][5] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\atari2600.ram[2][6] ),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\scanline[141][0] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\scanline[42][6] ),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\atari2600.ram[10][3] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\scanline[58][0] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\atari2600.ram[122][2] ),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\atari2600.ram[92][0] ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\external_rom_data[7] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1454 (.A(_01822_),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\atari2600.ram[21][0] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\scanline[54][2] ),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\atari2600.ram[82][0] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\scanline[51][5] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\atari2600.cpu.ABH[6] ),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01878_),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\scanline[40][6] ),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\scanline[77][6] ),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\atari2600.ram[53][2] ),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\atari2600.ram[114][6] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\atari2600.ram[4][7] ),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\scanline[30][3] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\scanline[157][1] ),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\atari2600.ram[6][4] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\scanline[15][1] ),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\atari2600.ram[58][0] ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\atari2600.ram[9][3] ),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\scanline[143][0] ),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\atari2600.ram[36][6] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\scanline[150][5] ),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\scanline[149][0] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\atari2600.ram[102][7] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\atari2600.ram[116][5] ),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\scanline[45][1] ),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\scanline[54][1] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\atari2600.ram[110][6] ),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\atari2600.tia.m1_w[2] ),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\atari2600.pia.swa_dir[1] ),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\atari2600.tia.poly9_r.x[8] ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_01230_),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\scanline[150][0] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\atari2600.ram[118][2] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\atari2600.ram[24][1] ),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\atari2600.ram[89][4] ),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\scanline[95][5] ),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\scanline[155][2] ),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\atari2600.tia.m0_w[3] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\atari2600.cpu.AXYS[2][0] ),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\atari2600.ram[42][0] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\gamepad_pmod.decoder.data_reg[2] ),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1495 (.A(_01554_),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\atari2600.tia.dat_o[6] ),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\atari2600.ram[112][1] ),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\flash_rom.addr_in[19] ),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1499 (.A(_00966_),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\scanline[119][3] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\scanline[117][0] ),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\atari2600.tia.p1_copies[1] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\scanline[159][0] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\gamepad_pmod.decoder.data_reg[10] ),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1505 (.A(_01562_),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\flash_rom.addr[22] ),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1507 (.A(_00981_),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\atari2600.tia.poly4_r.x[3] ),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_01216_),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\atari2600.ram[21][6] ),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\atari2600.ram[49][5] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\atari2600.ram[34][5] ),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\atari2600.ram[41][4] ),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\atari2600.tia.poly9_r.x[3] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_01225_),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\atari2600.cpu.PC[1] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_01411_),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\scanline[157][5] ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\scanline[155][1] ),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\scanline[31][3] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\scanline[159][4] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\atari2600.ram[16][1] ),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\gamepad_pmod.decoder.data_reg[5] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_01557_),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\atari2600.cpu.ABH[7] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_01879_),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\atari2600.ram[103][4] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\atari2600.ram[43][1] ),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\atari2600.tia.poly5_l.x[1] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold1530 (.A(_01199_),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\atari2600.ram[43][2] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\atari2600.pia.dat_o[6] ),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold1533 (.A(_00872_),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\atari2600.ram[102][4] ),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\atari2600.ram[70][5] ),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\scanline[118][5] ),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\atari2600.ram[107][5] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\atari2600.ram[108][5] ),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\atari2600.tia.m0_w[0] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\atari2600.pia.reset_timer[7] ),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\scanline[64][3] ),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\atari2600.ram[43][5] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\scanline[29][2] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\atari2600.cpu.IRHOLD[4] ),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\atari2600.ram[73][0] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\scanline[127][5] ),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\atari2600.ram[46][0] ),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\scanline[76][4] ),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\atari2600.pia.time_counter[10] ),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_05434_),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\atari2600.ram[39][7] ),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\atari2600.tia.cx[8] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\atari2600.cpu.PC[10] ),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_01420_),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\atari2600.cpu.ALU.AI7 ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\gamepad_pmod.decoder.data_reg[8] ),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_01560_),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\scanline[80][2] ),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\atari2600.ram[58][3] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\scanline[16][0] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\atari2600.ram[107][2] ),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\scanline[8][1] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\atari2600.ram[33][3] ),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\scanline[88][6] ),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\atari2600.pia.dat_o[1] ),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_00867_),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\atari2600.ram[11][7] ),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\atari2600.tia.m0_w[2] ),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\atari2600.ram[127][2] ),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\atari2600.ram[55][5] ),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\atari2600.cpu.AXYS[0][4] ),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold1572 (.A(_01309_),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\scanline[64][4] ),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\atari2600.ram[48][1] ),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\scanline[76][2] ),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\scanline[128][3] ),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\atari2600.pia.reset_timer[6] ),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\scanline[119][1] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\atari2600.ram[39][4] ),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\scanline[82][5] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\scanline[120][4] ),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\rom_last_read_addr[2] ),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_00266_),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\atari2600.tia.poly9_l.x[8] ),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold1585 (.A(_01211_),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\atari2600.ram[59][7] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\scanline[4][0] ),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\atari2600.ram[75][3] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\scanline[67][3] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\flash_rom.addr_in[17] ),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold1591 (.A(_00964_),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\atari2600.ram[59][4] ),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\scanline[9][6] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\scanline[66][6] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\atari2600.ram[28][5] ),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\atari2600.ram[2][7] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\scanline[66][3] ),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\atari2600.tia.old_grp1[4] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00919_),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\atari2600.ram[123][3] ),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\scanline[88][1] ),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\scanline[82][2] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\atari2600.ram[79][3] ),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\scanline[148][5] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\scanline[148][3] ),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\scanline[5][6] ),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\gamepad_pmod.driver.shift_reg[11] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_01487_),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold1609 (.A(_00161_),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold1610 (.A(_00095_),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_05994_),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold1612 (.A(_00991_),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\scanline[28][6] ),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\scanline[68][5] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\scanline[135][6] ),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\scanline[25][3] ),
    .X(net4543));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\scanline[2][4] ),
    .X(net4544));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\atari2600.ram[39][3] ),
    .X(net4545));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\scanline[20][0] ),
    .X(net4546));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\scanline[97][6] ),
    .X(net4547));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\scanline[0][3] ),
    .X(net4548));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\scanline[69][1] ),
    .X(net4549));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\scanline[33][6] ),
    .X(net4550));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\atari2600.ram[67][4] ),
    .X(net4551));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\scanline[82][3] ),
    .X(net4552));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\atari2600.ram[40][5] ),
    .X(net4553));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\scanline[20][1] ),
    .X(net4554));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\scanline[76][5] ),
    .X(net4555));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\atari2600.ram[36][4] ),
    .X(net4556));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\atari2600.ram[7][3] ),
    .X(net4557));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\scanline[136][3] ),
    .X(net4558));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\scanline[83][3] ),
    .X(net4559));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\scanline[40][4] ),
    .X(net4560));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\scanline[52][1] ),
    .X(net4561));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\scanline[83][1] ),
    .X(net4562));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\atari2600.ram[107][7] ),
    .X(net4563));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\scanline[73][6] ),
    .X(net4564));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\scanline[21][4] ),
    .X(net4565));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\atari2600.ram[35][6] ),
    .X(net4566));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\scanline[76][1] ),
    .X(net4567));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\atari2600.ram[79][5] ),
    .X(net4568));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\atari2600.ram[11][2] ),
    .X(net4569));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\scanline[39][0] ),
    .X(net4570));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\scanline[152][3] ),
    .X(net4571));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\scanline[22][5] ),
    .X(net4572));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\scanline[20][2] ),
    .X(net4573));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\atari2600.tia.diag[103] ),
    .X(net4574));
 sg13g2_dlygate4sd3_1 hold1648 (.A(_00922_),
    .X(net4575));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\atari2600.ram[75][5] ),
    .X(net4576));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\scanline[74][4] ),
    .X(net4577));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\scanline[7][5] ),
    .X(net4578));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\scanline[16][2] ),
    .X(net4579));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\atari2600.ram[35][1] ),
    .X(net4580));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\scanline[69][3] ),
    .X(net4581));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\scanline[42][2] ),
    .X(net4582));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\scanline[71][6] ),
    .X(net4583));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\scanline[112][0] ),
    .X(net4584));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\scanline[88][3] ),
    .X(net4585));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\scanline[19][6] ),
    .X(net4586));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\atari2600.ram[91][1] ),
    .X(net4587));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\scanline[128][4] ),
    .X(net4588));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\scanline[72][2] ),
    .X(net4589));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\atari2600.ram[39][5] ),
    .X(net4590));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\scanline[133][2] ),
    .X(net4591));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\scanline[28][5] ),
    .X(net4592));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\scanline[37][4] ),
    .X(net4593));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\scanline[81][0] ),
    .X(net4594));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\atari2600.ram[39][6] ),
    .X(net4595));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\atari2600.ram[99][1] ),
    .X(net4596));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\scanline[67][1] ),
    .X(net4597));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\scanline[50][4] ),
    .X(net4598));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\scanline[112][3] ),
    .X(net4599));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\atari2600.ram[19][3] ),
    .X(net4600));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\atari2600.ram[71][1] ),
    .X(net4601));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\scanline[28][2] ),
    .X(net4602));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\scanline[128][1] ),
    .X(net4603));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\scanline[83][4] ),
    .X(net4604));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\scanline[6][2] ),
    .X(net4605));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\scanline[129][0] ),
    .X(net4606));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\scanline[147][1] ),
    .X(net4607));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\scanline[97][5] ),
    .X(net4608));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\scanline[50][6] ),
    .X(net4609));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\scanline[28][0] ),
    .X(net4610));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\scanline[10][3] ),
    .X(net4611));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\scanline[80][5] ),
    .X(net4612));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\scanline[131][2] ),
    .X(net4613));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\scanline[134][3] ),
    .X(net4614));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\scanline[7][0] ),
    .X(net4615));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\atari2600.ram[7][1] ),
    .X(net4616));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\scanline[120][3] ),
    .X(net4617));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\scanline[137][3] ),
    .X(net4618));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\atari2600.ram[15][2] ),
    .X(net4619));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\atari2600.ram[15][4] ),
    .X(net4620));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\scanline[6][6] ),
    .X(net4621));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\scanline[84][4] ),
    .X(net4622));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\scanline[69][0] ),
    .X(net4623));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\scanline[133][5] ),
    .X(net4624));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\atari2600.ram[87][2] ),
    .X(net4625));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\scanline[104][3] ),
    .X(net4626));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\atari2600.pia.interval[6] ),
    .X(net4627));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\atari2600.ram[99][3] ),
    .X(net4628));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\atari2600.ram[75][0] ),
    .X(net4629));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\atari2600.ram[91][7] ),
    .X(net4630));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\scanline[128][5] ),
    .X(net4631));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\atari2600.ram[35][3] ),
    .X(net4632));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\scanline[3][4] ),
    .X(net4633));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\scanline[21][6] ),
    .X(net4634));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\atari2600.ram[115][4] ),
    .X(net4635));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\scanline[38][6] ),
    .X(net4636));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\scanline[40][0] ),
    .X(net4637));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\scanline[44][3] ),
    .X(net4638));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\atari2600.cpu.AXYS[0][2] ),
    .X(net4639));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\atari2600.cpu.IRHOLD[0] ),
    .X(net4640));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_01376_),
    .X(net4641));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\scanline[49][1] ),
    .X(net4642));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\atari2600.pia.dat_o[2] ),
    .X(net4643));
 sg13g2_dlygate4sd3_1 hold1717 (.A(_00868_),
    .X(net4644));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\scanline[28][4] ),
    .X(net4645));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\atari2600.ram[107][6] ),
    .X(net4646));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\atari2600.ram[27][7] ),
    .X(net4647));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\scanline[145][2] ),
    .X(net4648));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\atari2600.ram[63][7] ),
    .X(net4649));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\scanline[71][3] ),
    .X(net4650));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\scanline[2][2] ),
    .X(net4651));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\atari2600.ram[103][5] ),
    .X(net4652));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\scanline[11][1] ),
    .X(net4653));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\scanline[12][2] ),
    .X(net4654));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\atari2600.ram[27][0] ),
    .X(net4655));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\atari2600.ram[103][0] ),
    .X(net4656));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\scanline[134][0] ),
    .X(net4657));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\scanline[0][0] ),
    .X(net4658));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\scanline[75][4] ),
    .X(net4659));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\atari2600.ram[59][6] ),
    .X(net4660));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\scanline[7][1] ),
    .X(net4661));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\atari2600.ram[31][2] ),
    .X(net4662));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\atari2600.ram[15][1] ),
    .X(net4663));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\scanline[100][2] ),
    .X(net4664));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\scanline[69][6] ),
    .X(net4665));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\scanline[138][0] ),
    .X(net4666));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\atari2600.ram[95][3] ),
    .X(net4667));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\scanline[36][4] ),
    .X(net4668));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\scanline[140][6] ),
    .X(net4669));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\rom_last_read_addr[3] ),
    .X(net4670));
 sg13g2_dlygate4sd3_1 hold1744 (.A(_00267_),
    .X(net4671));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\scanline[97][4] ),
    .X(net4672));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\atari2600.ram[95][1] ),
    .X(net4673));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\scanline[145][4] ),
    .X(net4674));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\scanline[72][5] ),
    .X(net4675));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\atari2600.ram[35][4] ),
    .X(net4676));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\atari2600.ram[103][7] ),
    .X(net4677));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\atari2600.ram[23][2] ),
    .X(net4678));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\scanline[24][3] ),
    .X(net4679));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\atari2600.ram[47][2] ),
    .X(net4680));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\atari2600.ram[83][5] ),
    .X(net4681));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\atari2600.ram[43][6] ),
    .X(net4682));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\scanline[148][0] ),
    .X(net4683));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\scanline[71][4] ),
    .X(net4684));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\scanline[136][0] ),
    .X(net4685));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\scanline[116][5] ),
    .X(net4686));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\scanline[8][0] ),
    .X(net4687));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\scanline[34][5] ),
    .X(net4688));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\atari2600.ram[96][6] ),
    .X(net4689));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\atari2600.ram[115][0] ),
    .X(net4690));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\scanline[12][3] ),
    .X(net4691));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\scanline[129][5] ),
    .X(net4692));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\scanline[36][2] ),
    .X(net4693));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\scanline[84][6] ),
    .X(net4694));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\scanline[146][5] ),
    .X(net4695));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\atari2600.ram[59][1] ),
    .X(net4696));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\atari2600.ram[19][5] ),
    .X(net4697));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\scanline[112][2] ),
    .X(net4698));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\atari2600.ram[91][0] ),
    .X(net4699));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\scanline[139][1] ),
    .X(net4700));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\atari2600.ram[87][1] ),
    .X(net4701));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\atari2600.ram[23][4] ),
    .X(net4702));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\scanline[135][3] ),
    .X(net4703));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\atari2600.tia.diag[102] ),
    .X(net4704));
 sg13g2_dlygate4sd3_1 hold1778 (.A(_00921_),
    .X(net4705));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\scanline[18][4] ),
    .X(net4706));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\scanline[147][5] ),
    .X(net4707));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\scanline[68][2] ),
    .X(net4708));
 sg13g2_dlygate4sd3_1 hold1782 (.A(_00131_),
    .X(net4709));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\scanline[132][6] ),
    .X(net4710));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\atari2600.ram[115][6] ),
    .X(net4711));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\scanline[116][0] ),
    .X(net4712));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\scanline[25][2] ),
    .X(net4713));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\scanline[75][3] ),
    .X(net4714));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\atari2600.ram[23][0] ),
    .X(net4715));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\atari2600.ram[19][2] ),
    .X(net4716));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\scanline[139][5] ),
    .X(net4717));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\atari2600.ram[63][4] ),
    .X(net4718));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\scanline[81][4] ),
    .X(net4719));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\scanline[50][5] ),
    .X(net4720));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\scanline[65][3] ),
    .X(net4721));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\atari2600.ram[55][4] ),
    .X(net4722));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\atari2600.ram[18][5] ),
    .X(net4723));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\scanline[100][0] ),
    .X(net4724));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\scanline[65][4] ),
    .X(net4725));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\scanline[43][4] ),
    .X(net4726));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\scanline[9][1] ),
    .X(net4727));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\scanline[21][3] ),
    .X(net4728));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\scanline[5][0] ),
    .X(net4729));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\scanline[116][4] ),
    .X(net4730));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\scanline[136][6] ),
    .X(net4731));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\atari2600.cpu.AXYS[0][5] ),
    .X(net4732));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\scanline[132][3] ),
    .X(net4733));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\scanline[152][4] ),
    .X(net4734));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\atari2600.pia.reset_timer[3] ),
    .X(net4735));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\scanline[2][3] ),
    .X(net4736));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\atari2600.ram[95][4] ),
    .X(net4737));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\atari2600.ram[35][7] ),
    .X(net4738));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\scanline[48][5] ),
    .X(net4739));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\scanline[37][3] ),
    .X(net4740));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\atari2600.ram[111][1] ),
    .X(net4741));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\atari2600.ram[38][3] ),
    .X(net4742));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\atari2600.ram[23][3] ),
    .X(net4743));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\scanline[130][4] ),
    .X(net4744));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\scanline[17][5] ),
    .X(net4745));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\scanline[152][2] ),
    .X(net4746));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\scanline[131][3] ),
    .X(net4747));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\atari2600.ram[75][6] ),
    .X(net4748));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\scanline[156][6] ),
    .X(net4749));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\atari2600.ram[19][0] ),
    .X(net4750));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\scanline[67][0] ),
    .X(net4751));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\scanline[0][6] ),
    .X(net4752));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\scanline[2][0] ),
    .X(net4753));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\scanline[11][0] ),
    .X(net4754));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\scanline[76][3] ),
    .X(net4755));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\scanline[129][6] ),
    .X(net4756));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\scanline[129][2] ),
    .X(net4757));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\frame_counter[1] ),
    .X(net4758));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\scanline[40][3] ),
    .X(net4759));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\scanline[98][5] ),
    .X(net4760));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\atari2600.ram[43][0] ),
    .X(net4761));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\atari2600.ram[71][5] ),
    .X(net4762));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\atari2600.ram[23][5] ),
    .X(net4763));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\atari2600.ram[83][0] ),
    .X(net4764));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\scanline[64][1] ),
    .X(net4765));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\scanline[98][3] ),
    .X(net4766));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\scanline[97][1] ),
    .X(net4767));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\scanline[66][2] ),
    .X(net4768));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\scanline[56][6] ),
    .X(net4769));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\atari2600.ram[55][1] ),
    .X(net4770));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\atari2600.ram[42][7] ),
    .X(net4771));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\scanline[4][1] ),
    .X(net4772));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\scanline[97][2] ),
    .X(net4773));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\scanline[70][1] ),
    .X(net4774));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\scanline[148][4] ),
    .X(net4775));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\scanline[56][4] ),
    .X(net4776));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\scanline[42][5] ),
    .X(net4777));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\scanline[41][0] ),
    .X(net4778));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\atari2600.pia.dat_o[7] ),
    .X(net4779));
 sg13g2_dlygate4sd3_1 hold1853 (.A(_00873_),
    .X(net4780));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\scanline[71][2] ),
    .X(net4781));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\scanline[144][2] ),
    .X(net4782));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\scanline[22][0] ),
    .X(net4783));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\atari2600.ram[27][3] ),
    .X(net4784));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\scanline[88][5] ),
    .X(net4785));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\scanline[139][2] ),
    .X(net4786));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\scanline[35][0] ),
    .X(net4787));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\atari2600.ram[87][0] ),
    .X(net4788));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\scanline[120][0] ),
    .X(net4789));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\scanline[129][3] ),
    .X(net4790));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\atari2600.ram[103][3] ),
    .X(net4791));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\scanline[36][0] ),
    .X(net4792));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\external_rom_data[0] ),
    .X(net4793));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\scanline[82][1] ),
    .X(net4794));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\scanline[17][0] ),
    .X(net4795));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\scanline[3][6] ),
    .X(net4796));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\scanline[81][3] ),
    .X(net4797));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\atari2600.ram[7][0] ),
    .X(net4798));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\scanline[132][5] ),
    .X(net4799));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\scanline[44][4] ),
    .X(net4800));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\scanline[148][6] ),
    .X(net4801));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\scanline[33][4] ),
    .X(net4802));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\scanline[68][6] ),
    .X(net4803));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\atari2600.ram[79][0] ),
    .X(net4804));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\scanline[50][2] ),
    .X(net4805));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\scanline[83][2] ),
    .X(net4806));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\gamepad_pmod.decoder.data_reg[3] ),
    .X(net4807));
 sg13g2_dlygate4sd3_1 hold1881 (.A(_01555_),
    .X(net4808));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\scanline[0][2] ),
    .X(net4809));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\scanline[21][2] ),
    .X(net4810));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\atari2600.cpu.AXYS[0][6] ),
    .X(net4811));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\scanline[88][4] ),
    .X(net4812));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\atari2600.ram[95][6] ),
    .X(net4813));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\atari2600.ram[111][5] ),
    .X(net4814));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\scanline[48][1] ),
    .X(net4815));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\scanline[49][4] ),
    .X(net4816));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\atari2600.ram[127][5] ),
    .X(net4817));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\scanline[99][0] ),
    .X(net4818));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\atari2600.ram[59][3] ),
    .X(net4819));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\atari2600.ram[111][3] ),
    .X(net4820));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\scanline[152][6] ),
    .X(net4821));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\scanline[26][4] ),
    .X(net4822));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\scanline[24][0] ),
    .X(net4823));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\scanline[137][0] ),
    .X(net4824));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\atari2600.ram[35][0] ),
    .X(net4825));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\scanline[152][1] ),
    .X(net4826));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\scanline[133][4] ),
    .X(net4827));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\scanline[144][1] ),
    .X(net4828));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\scanline[24][6] ),
    .X(net4829));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\atari2600.ram[19][4] ),
    .X(net4830));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\atari2600.ram[27][1] ),
    .X(net4831));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\atari2600.ram[47][5] ),
    .X(net4832));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\atari2600.ram[63][0] ),
    .X(net4833));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\scanline[35][1] ),
    .X(net4834));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\atari2600.ram[115][5] ),
    .X(net4835));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\scanline[98][2] ),
    .X(net4836));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\atari2600.ram[79][6] ),
    .X(net4837));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\atari2600.ram[39][2] ),
    .X(net4838));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\atari2600.ram[87][7] ),
    .X(net4839));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\scanline[131][0] ),
    .X(net4840));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\atari2600.ram[45][0] ),
    .X(net4841));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\scanline[4][4] ),
    .X(net4842));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\scanline[9][2] ),
    .X(net4843));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\scanline[128][0] ),
    .X(net4844));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\scanline[32][0] ),
    .X(net4845));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\external_rom_data[2] ),
    .X(net4846));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\atari2600.ram[31][3] ),
    .X(net4847));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\scanline[16][3] ),
    .X(net4848));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\scanline[34][3] ),
    .X(net4849));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\atari2600.ram[119][4] ),
    .X(net4850));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\scanline[75][1] ),
    .X(net4851));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\atari2600.ram[15][0] ),
    .X(net4852));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\scanline[144][5] ),
    .X(net4853));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\scanline[10][0] ),
    .X(net4854));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\scanline[49][0] ),
    .X(net4855));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\scanline[49][3] ),
    .X(net4856));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\atari2600.ram[91][4] ),
    .X(net4857));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\scanline[130][2] ),
    .X(net4858));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\atari2600.ram[79][2] ),
    .X(net4859));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\scanline[147][6] ),
    .X(net4860));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\scanline[80][3] ),
    .X(net4861));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\scanline[7][6] ),
    .X(net4862));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\scanline[19][1] ),
    .X(net4863));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\scanline[10][2] ),
    .X(net4864));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\scanline[100][6] ),
    .X(net4865));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\atari2600.tia.poly5_r.x[3] ),
    .X(net4866));
 sg13g2_dlygate4sd3_1 hold1940 (.A(_01219_),
    .X(net4867));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\scanline[32][3] ),
    .X(net4868));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\scanline[16][4] ),
    .X(net4869));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\scanline[69][5] ),
    .X(net4870));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\scanline[35][6] ),
    .X(net4871));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\scanline[33][2] ),
    .X(net4872));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\atari2600.ram[59][0] ),
    .X(net4873));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\scanline[133][1] ),
    .X(net4874));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\atari2600.ram[119][0] ),
    .X(net4875));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\scanline[56][5] ),
    .X(net4876));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\atari2600.ram[107][0] ),
    .X(net4877));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\atari2600.ram[83][4] ),
    .X(net4878));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\atari2600.ram[55][0] ),
    .X(net4879));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\scanline[37][5] ),
    .X(net4880));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\scanline[80][4] ),
    .X(net4881));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\scanline[0][5] ),
    .X(net4882));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\scanline[41][1] ),
    .X(net4883));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\scanline[32][1] ),
    .X(net4884));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\atari2600.ram[127][7] ),
    .X(net4885));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\scanline[12][1] ),
    .X(net4886));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\atari2600.ram[95][2] ),
    .X(net4887));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\scanline[50][1] ),
    .X(net4888));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\scanline[137][2] ),
    .X(net4889));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\scanline[68][3] ),
    .X(net4890));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\scanline[10][1] ),
    .X(net4891));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\scanline[73][4] ),
    .X(net4892));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\atari2600.ram[127][3] ),
    .X(net4893));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\scanline[40][5] ),
    .X(net4894));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\scanline[49][2] ),
    .X(net4895));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\scanline[6][5] ),
    .X(net4896));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\scanline[147][4] ),
    .X(net4897));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\atari2600.ram[63][5] ),
    .X(net4898));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\atari2600.ram[87][4] ),
    .X(net4899));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\atari2600.ram[119][7] ),
    .X(net4900));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\scanline[12][0] ),
    .X(net4901));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\scanline[36][3] ),
    .X(net4902));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\external_rom_data[3] ),
    .X(net4903));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\scanline[8][4] ),
    .X(net4904));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\scanline[99][3] ),
    .X(net4905));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\atari2600.ram[31][6] ),
    .X(net4906));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\atari2600.ram[91][2] ),
    .X(net4907));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\atari2600.ram[59][2] ),
    .X(net4908));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\scanline[99][4] ),
    .X(net4909));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\atari2600.ram[111][0] ),
    .X(net4910));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\atari2600.ram[75][7] ),
    .X(net4911));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\scanline[65][1] ),
    .X(net4912));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\scanline[50][3] ),
    .X(net4913));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\scanline[81][1] ),
    .X(net4914));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\atari2600.ram[83][3] ),
    .X(net4915));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\atari2600.ram[47][4] ),
    .X(net4916));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\atari2600.ram[119][2] ),
    .X(net4917));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\scanline[139][3] ),
    .X(net4918));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\rom_last_read_addr[8] ),
    .X(net4919));
 sg13g2_dlygate4sd3_1 hold1993 (.A(_00272_),
    .X(net4920));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\atari2600.ram[11][6] ),
    .X(net4921));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\scanline[136][1] ),
    .X(net4922));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\scanline[137][4] ),
    .X(net4923));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\scanline[21][5] ),
    .X(net4924));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\scanline[1][6] ),
    .X(net4925));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\scanline[137][5] ),
    .X(net4926));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\scanline[65][0] ),
    .X(net4927));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\scanline[73][1] ),
    .X(net4928));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\atari2600.ram[19][6] ),
    .X(net4929));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\scanline[40][2] ),
    .X(net4930));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\scanline[40][1] ),
    .X(net4931));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\scanline[80][6] ),
    .X(net4932));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\scanline[23][3] ),
    .X(net4933));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\scanline[41][2] ),
    .X(net4934));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\scanline[96][1] ),
    .X(net4935));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\scanline[145][3] ),
    .X(net4936));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\atari2600.cpu.D ),
    .X(net4937));
 sg13g2_dlygate4sd3_1 hold2011 (.A(_00022_),
    .X(net4938));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\scanline[83][5] ),
    .X(net4939));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\atari2600.ram[31][5] ),
    .X(net4940));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\atari2600.tia.old_grp1[3] ),
    .X(net4941));
 sg13g2_dlygate4sd3_1 hold2015 (.A(_00918_),
    .X(net4942));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\scanline[70][5] ),
    .X(net4943));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\atari2600.ram[87][3] ),
    .X(net4944));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\scanline[64][6] ),
    .X(net4945));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\scanline[16][6] ),
    .X(net4946));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\scanline[35][3] ),
    .X(net4947));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\scanline[33][5] ),
    .X(net4948));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\scanline[8][5] ),
    .X(net4949));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\atari2600.ram[68][3] ),
    .X(net4950));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\scanline[66][1] ),
    .X(net4951));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\atari2600.ram[63][3] ),
    .X(net4952));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\scanline[56][0] ),
    .X(net4953));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\atari2600.ram[7][5] ),
    .X(net4954));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\atari2600.ram[119][5] ),
    .X(net4955));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\scanline[33][0] ),
    .X(net4956));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\scanline[67][2] ),
    .X(net4957));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\scanline[8][2] ),
    .X(net4958));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\scanline[39][4] ),
    .X(net4959));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\atari2600.pia.reset_timer[4] ),
    .X(net4960));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\scanline[104][1] ),
    .X(net6583));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\scanline[70][2] ),
    .X(net6584));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\atari2600.ram[27][6] ),
    .X(net6585));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\atari2600.ram[67][0] ),
    .X(net6586));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\scanline[128][6] ),
    .X(net6587));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\scanline[5][3] ),
    .X(net6588));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\atari2600.ram[63][2] ),
    .X(net6589));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\scanline[100][3] ),
    .X(net6590));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\atari2600.ram[71][2] ),
    .X(net6591));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\atari2600.tia.audf1[4] ),
    .X(net6592));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\atari2600.ram[75][1] ),
    .X(net6593));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\scanline[104][2] ),
    .X(net6594));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\scanline[52][2] ),
    .X(net6595));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\atari2600.ram[27][5] ),
    .X(net6596));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\atari2600.pia.time_counter[15] ),
    .X(net6597));
 sg13g2_dlygate4sd3_1 hold2049 (.A(_00889_),
    .X(net6598));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\scanline[44][0] ),
    .X(net6599));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\scanline[44][5] ),
    .X(net6600));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\atari2600.ram[31][7] ),
    .X(net6601));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\scanline[72][3] ),
    .X(net6602));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\scanline[88][0] ),
    .X(net6603));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\scanline[116][3] ),
    .X(net6604));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\scanline[100][1] ),
    .X(net6605));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\scanline[16][5] ),
    .X(net6606));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\atari2600.ram[23][1] ),
    .X(net6607));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\atari2600.ram[67][3] ),
    .X(net6608));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\scanline[67][5] ),
    .X(net6609));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\atari2600.ram[119][6] ),
    .X(net6610));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\scanline[68][4] ),
    .X(net6611));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\atari2600.pia.time_counter[21] ),
    .X(net6612));
 sg13g2_dlygate4sd3_1 hold2064 (.A(_05460_),
    .X(net6613));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\scanline[66][4] ),
    .X(net6614));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\scanline[26][1] ),
    .X(net6615));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\scanline[80][0] ),
    .X(net6616));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\scanline[37][2] ),
    .X(net6617));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\atari2600.ram[7][4] ),
    .X(net6618));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\atari2600.ram[123][4] ),
    .X(net6619));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\scanline[100][4] ),
    .X(net6620));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\scanline[12][4] ),
    .X(net6621));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\scanline[145][1] ),
    .X(net6622));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\scanline[72][6] ),
    .X(net6623));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\scanline[16][1] ),
    .X(net6624));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\scanline[34][4] ),
    .X(net6625));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\rom_last_read_addr[4] ),
    .X(net6626));
 sg13g2_dlygate4sd3_1 hold2078 (.A(_00268_),
    .X(net6627));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\atari2600.ram[35][2] ),
    .X(net6628));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\scanline[0][1] ),
    .X(net6629));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\atari2600.ram[91][6] ),
    .X(net6630));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\atari2600.cpu.AXYS[0][3] ),
    .X(net6631));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\scanline[135][2] ),
    .X(net6632));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\atari2600.ram[15][7] ),
    .X(net6633));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\scanline[134][4] ),
    .X(net6634));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\scanline[23][5] ),
    .X(net6635));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\scanline[11][3] ),
    .X(net6636));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\scanline[137][1] ),
    .X(net6637));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\atari2600.ram[91][3] ),
    .X(net6638));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\scanline[99][6] ),
    .X(net6639));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\atari2600.ram[43][4] ),
    .X(net6640));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\atari2600.ram[39][1] ),
    .X(net6641));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\atari2600.ram[31][0] ),
    .X(net6642));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\atari2600.ram[7][7] ),
    .X(net6643));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\atari2600.ram[115][2] ),
    .X(net6644));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\scanline[12][6] ),
    .X(net6645));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\atari2600.ram[59][5] ),
    .X(net6646));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\scanline[131][1] ),
    .X(net6647));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\scanline[116][2] ),
    .X(net6648));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\scanline[1][1] ),
    .X(net6649));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\scanline[128][2] ),
    .X(net6650));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\atari2600.ram[111][6] ),
    .X(net6651));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\scanline[28][3] ),
    .X(net6652));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\scanline[135][4] ),
    .X(net6653));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\scanline[2][1] ),
    .X(net6654));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\atari2600.ram[55][2] ),
    .X(net6655));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\atari2600.ram[87][6] ),
    .X(net6656));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\scanline[146][1] ),
    .X(net6657));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\scanline[74][1] ),
    .X(net6658));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\scanline[26][3] ),
    .X(net6659));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\scanline[116][6] ),
    .X(net6660));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\atari2600.ram[103][6] ),
    .X(net6661));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\atari2600.ram[123][5] ),
    .X(net6662));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\scanline[1][5] ),
    .X(net6663));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\scanline[140][4] ),
    .X(net6664));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\scanline[84][0] ),
    .X(net6665));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\atari2600.ram[15][5] ),
    .X(net6666));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\scanline[41][5] ),
    .X(net6667));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\atari2600.tia.refp0 ),
    .X(net6668));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\atari2600.ram[127][6] ),
    .X(net6669));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\atari2600.ram[71][3] ),
    .X(net6670));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\atari2600.cpu.AXYS[0][0] ),
    .X(net6671));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\scanline[35][2] ),
    .X(net6672));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\atari2600.ram[67][1] ),
    .X(net6673));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\atari2600.ram[127][0] ),
    .X(net6674));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\scanline[146][0] ),
    .X(net6675));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\atari2600.ram[95][7] ),
    .X(net6676));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\scanline[138][4] ),
    .X(net6677));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\gamepad_pmod.driver.shift_reg[5] ),
    .X(net6678));
 sg13g2_dlygate4sd3_1 hold2130 (.A(_01481_),
    .X(net6679));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\scanline[134][2] ),
    .X(net6680));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\atari2600.ram[127][1] ),
    .X(net6681));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\scanline[26][2] ),
    .X(net6682));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\scanline[70][4] ),
    .X(net6683));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\scanline[144][3] ),
    .X(net6684));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\scanline[2][6] ),
    .X(net6685));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\atari2600.ram[47][0] ),
    .X(net6686));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\scanline[130][5] ),
    .X(net6687));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\scanline[81][5] ),
    .X(net6688));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\scanline[67][6] ),
    .X(net6689));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\scanline[4][3] ),
    .X(net6690));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\atari2600.ram[79][7] ),
    .X(net6691));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\atari2600.ram[111][4] ),
    .X(net6692));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\scanline[3][2] ),
    .X(net6693));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\atari2600.ram[63][6] ),
    .X(net6694));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\atari2600.ram[107][1] ),
    .X(net6695));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\scanline[144][6] ),
    .X(net6696));
 sg13g2_dlygate4sd3_1 hold2148 (.A(\atari2600.ram[15][6] ),
    .X(net6697));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\scanline[120][6] ),
    .X(net6698));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\scanline[147][2] ),
    .X(net6699));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\scanline[39][1] ),
    .X(net6700));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\scanline[17][3] ),
    .X(net6701));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\atari2600.tia.m1_w[1] ),
    .X(net6702));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\scanline[70][3] ),
    .X(net6703));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\scanline[38][3] ),
    .X(net6704));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\scanline[11][2] ),
    .X(net6705));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\scanline[144][0] ),
    .X(net6706));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\scanline[140][1] ),
    .X(net6707));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\atari2600.ram[47][7] ),
    .X(net6708));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\gamepad_pmod.driver.shift_reg[4] ),
    .X(net6709));
 sg13g2_dlygate4sd3_1 hold2161 (.A(_01480_),
    .X(net6710));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\scanline[84][2] ),
    .X(net6711));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\atari2600.ram[55][7] ),
    .X(net6712));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\scanline[97][3] ),
    .X(net6713));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\scanline[6][3] ),
    .X(net6714));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\atari2600.ram[67][7] ),
    .X(net6715));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\gamepad_pmod.driver.shift_reg[6] ),
    .X(net6716));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\scanline[132][2] ),
    .X(net6717));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\scanline[23][1] ),
    .X(net6718));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\scanline[65][2] ),
    .X(net6719));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\scanline[75][2] ),
    .X(net6720));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\scanline[17][1] ),
    .X(net6721));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\scanline[72][4] ),
    .X(net6722));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\scanline[6][1] ),
    .X(net6723));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\scanline[44][6] ),
    .X(net6724));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\atari2600.ram[99][4] ),
    .X(net6725));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\scanline[139][0] ),
    .X(net6726));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\scanline[25][4] ),
    .X(net6727));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\scanline[25][1] ),
    .X(net6728));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\scanline[23][0] ),
    .X(net6729));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\scanline[43][0] ),
    .X(net6730));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\scanline[120][5] ),
    .X(net6731));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\scanline[27][4] ),
    .X(net6732));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\scanline[76][6] ),
    .X(net6733));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\scanline[130][0] ),
    .X(net6734));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\atari2600.ram[23][6] ),
    .X(net6735));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\scanline[72][0] ),
    .X(net6736));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\scanline[98][0] ),
    .X(net6737));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\scanline[72][1] ),
    .X(net6738));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\atari2600.ram[83][7] ),
    .X(net6739));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\scanline[134][5] ),
    .X(net6740));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\scanline[99][1] ),
    .X(net6741));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\scanline[75][0] ),
    .X(net6742));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\atari2600.ram[31][4] ),
    .X(net6743));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\scanline[38][0] ),
    .X(net6744));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\scanline[20][3] ),
    .X(net6745));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\scanline[98][6] ),
    .X(net6746));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\scanline[52][5] ),
    .X(net6747));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\scanline[32][4] ),
    .X(net6748));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\atari2600.ram[115][3] ),
    .X(net6749));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\scanline[5][4] ),
    .X(net6750));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\scanline[6][0] ),
    .X(net6751));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\scanline[129][1] ),
    .X(net6752));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\scanline[32][2] ),
    .X(net6753));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\atari2600.ram[71][4] ),
    .X(net6754));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\scanline[96][4] ),
    .X(net6755));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\scanline[70][6] ),
    .X(net6756));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\scanline[3][3] ),
    .X(net6757));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\scanline[49][6] ),
    .X(net6758));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\scanline[4][5] ),
    .X(net6759));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\scanline[135][0] ),
    .X(net6760));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\scanline[147][0] ),
    .X(net6761));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\atari2600.ram[99][6] ),
    .X(net6762));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\atari2600.ram[95][0] ),
    .X(net6763));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\atari2600.tia.diag[97] ),
    .X(net6764));
 sg13g2_dlygate4sd3_1 hold2216 (.A(_00916_),
    .X(net6765));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\scanline[7][3] ),
    .X(net6766));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\atari2600.ram[11][1] ),
    .X(net6767));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\scanline[36][5] ),
    .X(net6768));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\scanline[4][6] ),
    .X(net6769));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\scanline[152][0] ),
    .X(net6770));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\scanline[52][6] ),
    .X(net6771));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\scanline[34][0] ),
    .X(net6772));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\scanline[96][0] ),
    .X(net6773));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\atari2600.ram[19][7] ),
    .X(net6774));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\scanline[18][6] ),
    .X(net6775));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\scanline[99][5] ),
    .X(net6776));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\scanline[73][5] ),
    .X(net6777));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\scanline[10][5] ),
    .X(net6778));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\atari2600.ram[43][7] ),
    .X(net6779));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\scanline[21][1] ),
    .X(net6780));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\scanline[146][2] ),
    .X(net6781));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\scanline[130][1] ),
    .X(net6782));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\scanline[7][2] ),
    .X(net6783));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\scanline[140][5] ),
    .X(net6784));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\scanline[138][2] ),
    .X(net6785));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\scanline[24][2] ),
    .X(net6786));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\scanline[74][3] ),
    .X(net6787));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\scanline[120][1] ),
    .X(net6788));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\scanline[97][0] ),
    .X(net6789));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\scanline[52][3] ),
    .X(net6790));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\scanline[22][1] ),
    .X(net6791));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\scanline[133][6] ),
    .X(net6792));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\scanline[9][5] ),
    .X(net6793));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\atari2600.ram[99][0] ),
    .X(net6794));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\scanline[144][4] ),
    .X(net6795));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\atari2600.ram[47][6] ),
    .X(net6796));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\scanline[140][2] ),
    .X(net6797));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\scanline[83][6] ),
    .X(net6798));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\scanline[81][2] ),
    .X(net6799));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\scanline[34][2] ),
    .X(net6800));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\scanline[130][3] ),
    .X(net6801));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\atari2600.ram[127][4] ),
    .X(net6802));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\scanline[43][2] ),
    .X(net6803));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\atari2600.ram[47][1] ),
    .X(net6804));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\scanline[56][2] ),
    .X(net6805));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\scanline[32][5] ),
    .X(net6806));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\atari2600.ram[115][1] ),
    .X(net6807));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\scanline[41][6] ),
    .X(net6808));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\gamepad_pmod.driver.shift_reg[10] ),
    .X(net6809));
 sg13g2_dlygate4sd3_1 hold2261 (.A(_01486_),
    .X(net6810));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\scanline[74][5] ),
    .X(net6811));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\atari2600.ram[47][3] ),
    .X(net6812));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\scanline[104][0] ),
    .X(net6813));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\scanline[21][0] ),
    .X(net6814));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\atari2600.tia.poly5_r.x[1] ),
    .X(net6815));
 sg13g2_dlygate4sd3_1 hold2267 (.A(_01217_),
    .X(net6816));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\scanline[27][2] ),
    .X(net6817));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\scanline[145][6] ),
    .X(net6818));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\scanline[48][2] ),
    .X(net6819));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\scanline[23][4] ),
    .X(net6820));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\atari2600.ram[19][1] ),
    .X(net6821));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\scanline[56][3] ),
    .X(net6822));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\scanline[138][1] ),
    .X(net6823));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\atari2600.cpu.sec ),
    .X(net6824));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\atari2600.ram[11][5] ),
    .X(net6825));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\scanline[120][2] ),
    .X(net6826));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\scanline[80][1] ),
    .X(net6827));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\scanline[71][0] ),
    .X(net6828));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\scanline[52][0] ),
    .X(net6829));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\scanline[42][4] ),
    .X(net6830));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\scanline[147][3] ),
    .X(net6831));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\scanline[12][5] ),
    .X(net6832));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\scanline[82][6] ),
    .X(net6833));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\scanline[24][1] ),
    .X(net6834));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\scanline[28][1] ),
    .X(net6835));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\scanline[67][4] ),
    .X(net6836));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\scanline[10][6] ),
    .X(net6837));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\atari2600.ram[79][4] ),
    .X(net6838));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\scanline[23][6] ),
    .X(net6839));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\scanline[148][1] ),
    .X(net6840));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\scanline[1][3] ),
    .X(net6841));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\scanline[136][4] ),
    .X(net6842));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\scanline[112][5] ),
    .X(net6843));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\scanline[32][6] ),
    .X(net6844));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\gamepad_pmod.decoder.data_reg[9] ),
    .X(net6845));
 sg13g2_dlygate4sd3_1 hold2297 (.A(_01561_),
    .X(net6846));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\scanline[98][1] ),
    .X(net6847));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\scanline[43][3] ),
    .X(net6848));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\scanline[99][2] ),
    .X(net6849));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\scanline[25][0] ),
    .X(net6850));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\atari2600.ram[107][3] ),
    .X(net6851));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\scanline[140][0] ),
    .X(net6852));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\scanline[1][0] ),
    .X(net6853));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\scanline[39][5] ),
    .X(net6854));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\scanline[2][5] ),
    .X(net6855));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\scanline[66][5] ),
    .X(net6856));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\scanline[39][2] ),
    .X(net6857));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\scanline[3][0] ),
    .X(net6858));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\scanline[33][3] ),
    .X(net6859));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\scanline[27][0] ),
    .X(net6860));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\scanline[17][2] ),
    .X(net6861));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\scanline[71][1] ),
    .X(net6862));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\scanline[75][6] ),
    .X(net6863));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\atari2600.cpu.PC[8] ),
    .X(net6864));
 sg13g2_dlygate4sd3_1 hold2316 (.A(_01418_),
    .X(net6865));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\scanline[42][0] ),
    .X(net6866));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\scanline[17][4] ),
    .X(net6867));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\scanline[27][5] ),
    .X(net6868));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\scanline[73][2] ),
    .X(net6869));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\scanline[74][0] ),
    .X(net6870));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\scanline[48][3] ),
    .X(net6871));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\scanline[26][5] ),
    .X(net6872));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\atari2600.tia.poly4_l.x[2] ),
    .X(net6873));
 sg13g2_dlygate4sd3_1 hold2325 (.A(_01196_),
    .X(net6874));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\scanline[73][0] ),
    .X(net6875));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\scanline[104][4] ),
    .X(net6876));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\scanline[18][3] ),
    .X(net6877));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\scanline[10][4] ),
    .X(net6878));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\atari2600.tia.m0_w[1] ),
    .X(net6879));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\scanline[131][4] ),
    .X(net6880));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\scanline[33][1] ),
    .X(net6881));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\scanline[25][5] ),
    .X(net6882));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\scanline[82][4] ),
    .X(net6883));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\scanline[84][1] ),
    .X(net6884));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\scanline[27][3] ),
    .X(net6885));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\scanline[5][5] ),
    .X(net6886));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\scanline[146][6] ),
    .X(net6887));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\scanline[36][6] ),
    .X(net6888));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\atari2600.ram[83][2] ),
    .X(net6889));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\scanline[152][5] ),
    .X(net6890));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\scanline[0][4] ),
    .X(net6891));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\scanline[68][0] ),
    .X(net6892));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\scanline[88][2] ),
    .X(net6893));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\atari2600.ram[63][1] ),
    .X(net6894));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\scanline[43][5] ),
    .X(net6895));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\atari2600.ram[119][3] ),
    .X(net6896));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\scanline[17][6] ),
    .X(net6897));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\scanline[36][1] ),
    .X(net6898));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\scanline[68][1] ),
    .X(net6899));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\atari2600.ram[123][6] ),
    .X(net6900));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\scanline[112][1] ),
    .X(net6901));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\scanline[24][5] ),
    .X(net6902));
 sg13g2_dlygate4sd3_1 hold2354 (.A(\scanline[138][3] ),
    .X(net6903));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\scanline[139][6] ),
    .X(net6904));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\scanline[3][5] ),
    .X(net6905));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\scanline[139][4] ),
    .X(net6906));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\scanline[48][0] ),
    .X(net6907));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\atari2600.ram[3][1] ),
    .X(net6908));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\scanline[27][6] ),
    .X(net6909));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\atari2600.ram[107][4] ),
    .X(net6910));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\atari2600.ram[79][1] ),
    .X(net6911));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\scanline[64][5] ),
    .X(net6912));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\atari2600.ram[83][1] ),
    .X(net6913));
 sg13g2_dlygate4sd3_1 hold2365 (.A(\scanline[41][4] ),
    .X(net6914));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\atari2600.ram[99][2] ),
    .X(net6915));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\atari2600.tia.poly5_l.x[2] ),
    .X(net6916));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\scanline[132][0] ),
    .X(net6917));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\scanline[96][3] ),
    .X(net6918));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\atari2600.ram[99][5] ),
    .X(net6919));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\scanline[133][3] ),
    .X(net6920));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\scanline[138][5] ),
    .X(net6921));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\scanline[64][2] ),
    .X(net6922));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\scanline[41][3] ),
    .X(net6923));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\gamepad_pmod.driver.shift_reg[1] ),
    .X(net6924));
 sg13g2_dlygate4sd3_1 hold2376 (.A(_01477_),
    .X(net6925));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\scanline[43][1] ),
    .X(net6926));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\scanline[37][6] ),
    .X(net6927));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\atari2600.ram[7][2] ),
    .X(net6928));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\scanline[96][6] ),
    .X(net6929));
 sg13g2_dlygate4sd3_1 hold2381 (.A(\atari2600.ram[31][1] ),
    .X(net6930));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\scanline[25][6] ),
    .X(net6931));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\scanline[48][6] ),
    .X(net6932));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\scanline[49][5] ),
    .X(net6933));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\scanline[52][4] ),
    .X(net6934));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\scanline[98][4] ),
    .X(net6935));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\scanline[70][0] ),
    .X(net6936));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\scanline[82][0] ),
    .X(net6937));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\scanline[1][4] ),
    .X(net6938));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\atari2600.ram[7][6] ),
    .X(net6939));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\scanline[39][3] ),
    .X(net6940));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\atari2600.pia.reset_timer[5] ),
    .X(net6941));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\scanline[35][5] ),
    .X(net6942));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\scanline[75][5] ),
    .X(net6943));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\scanline[134][6] ),
    .X(net6944));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\atari2600.tia.poly9_l.x[6] ),
    .X(net6945));
 sg13g2_dlygate4sd3_1 hold2397 (.A(_01209_),
    .X(net6946));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\atari2600.ram[99][7] ),
    .X(net6947));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\scanline[8][3] ),
    .X(net6948));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\scanline[22][3] ),
    .X(net6949));
 sg13g2_dlygate4sd3_1 hold2401 (.A(\atari2600.ram[119][1] ),
    .X(net6950));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\scanline[66][0] ),
    .X(net6951));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\scanline[148][2] ),
    .X(net6952));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\scanline[69][4] ),
    .X(net6953));
 sg13g2_dlygate4sd3_1 hold2405 (.A(\scanline[104][6] ),
    .X(net6954));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\atari2600.ram[71][6] ),
    .X(net6955));
 sg13g2_dlygate4sd3_1 hold2407 (.A(\scanline[11][6] ),
    .X(net6956));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\scanline[37][0] ),
    .X(net6957));
 sg13g2_dlygate4sd3_1 hold2409 (.A(\atari2600.ram[75][4] ),
    .X(net6958));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\scanline[38][2] ),
    .X(net6959));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\scanline[76][0] ),
    .X(net6960));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\scanline[96][2] ),
    .X(net6961));
 sg13g2_dlygate4sd3_1 hold2413 (.A(\atari2600.ram[27][4] ),
    .X(net6962));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\atari2600.ram[11][3] ),
    .X(net6963));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\rom_last_read_addr[11] ),
    .X(net6964));
 sg13g2_dlygate4sd3_1 hold2416 (.A(_00275_),
    .X(net6965));
 sg13g2_dlygate4sd3_1 hold2417 (.A(\scanline[135][5] ),
    .X(net6966));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\scanline[146][4] ),
    .X(net6967));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\scanline[35][4] ),
    .X(net6968));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\scanline[65][6] ),
    .X(net6969));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\atari2600.ram[123][7] ),
    .X(net6970));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\scanline[1][2] ),
    .X(net6971));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\scanline[84][5] ),
    .X(net6972));
 sg13g2_dlygate4sd3_1 hold2424 (.A(\scanline[22][2] ),
    .X(net6973));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\scanline[112][4] ),
    .X(net6974));
 sg13g2_dlygate4sd3_1 hold2426 (.A(\scanline[133][0] ),
    .X(net6975));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\scanline[74][6] ),
    .X(net6976));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\scanline[132][4] ),
    .X(net6977));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\scanline[84][3] ),
    .X(net6978));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\atari2600.tia.poly9_l.x[7] ),
    .X(net6979));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\atari2600.tia.diag[80] ),
    .X(net6980));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\atari2600.ram[67][6] ),
    .X(net6981));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\scanline[34][6] ),
    .X(net6982));
 sg13g2_dlygate4sd3_1 hold2434 (.A(\scanline[18][5] ),
    .X(net6983));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\atari2600.tia.poly5_r.x[4] ),
    .X(net6984));
 sg13g2_dlygate4sd3_1 hold2436 (.A(_01221_),
    .X(net6985));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\scanline[71][5] ),
    .X(net6986));
 sg13g2_dlygate4sd3_1 hold2438 (.A(\atari2600.ram[67][5] ),
    .X(net6987));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\scanline[18][1] ),
    .X(net6988));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\atari2600.pia.swa_dir[7] ),
    .X(net6989));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\scanline[34][1] ),
    .X(net6990));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\scanline[9][4] ),
    .X(net6991));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\scanline[136][5] ),
    .X(net6992));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\scanline[20][4] ),
    .X(net6993));
 sg13g2_dlygate4sd3_1 hold2445 (.A(\scanline[137][6] ),
    .X(net6994));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\scanline[131][6] ),
    .X(net6995));
 sg13g2_dlygate4sd3_1 hold2447 (.A(\scanline[132][1] ),
    .X(net6996));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\scanline[138][6] ),
    .X(net6997));
 sg13g2_dlygate4sd3_1 hold2449 (.A(\scanline[22][4] ),
    .X(net6998));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\atari2600.ram[111][2] ),
    .X(net6999));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\scanline[5][1] ),
    .X(net7000));
 sg13g2_dlygate4sd3_1 hold2452 (.A(\scanline[39][6] ),
    .X(net7001));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\scanline[64][0] ),
    .X(net7002));
 sg13g2_dlygate4sd3_1 hold2454 (.A(\atari2600.cpu.ABL[2] ),
    .X(net7003));
 sg13g2_dlygate4sd3_1 hold2455 (.A(_01393_),
    .X(net7004));
 sg13g2_dlygate4sd3_1 hold2456 (.A(\scanline[27][1] ),
    .X(net7005));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\scanline[38][4] ),
    .X(net7006));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\scanline[134][1] ),
    .X(net7007));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\atari2600.cpu.PC[4] ),
    .X(net7008));
 sg13g2_dlygate4sd3_1 hold2460 (.A(_01414_),
    .X(net7009));
 sg13g2_dlygate4sd3_1 hold2461 (.A(\scanline[42][1] ),
    .X(net7010));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\scanline[3][1] ),
    .X(net7011));
 sg13g2_dlygate4sd3_1 hold2463 (.A(\atari2600.ram[75][2] ),
    .X(net7012));
 sg13g2_dlygate4sd3_1 hold2464 (.A(\atari2600.ram[43][3] ),
    .X(net7013));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\atari2600.ram[103][1] ),
    .X(net7014));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\atari2600.ram[83][6] ),
    .X(net7015));
 sg13g2_dlygate4sd3_1 hold2467 (.A(\atari2600.ram[115][7] ),
    .X(net7016));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\scanline[73][3] ),
    .X(net7017));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\atari2600.pia.time_counter[8] ),
    .X(net7018));
 sg13g2_dlygate4sd3_1 hold2470 (.A(_00882_),
    .X(net7019));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\scanline[81][6] ),
    .X(net7020));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\scanline[23][2] ),
    .X(net7021));
 sg13g2_dlygate4sd3_1 hold2473 (.A(\scanline[22][6] ),
    .X(net7022));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\atari2600.ram[27][2] ),
    .X(net7023));
 sg13g2_dlygate4sd3_1 hold2475 (.A(\atari2600.pia.time_counter[16] ),
    .X(net7024));
 sg13g2_dlygate4sd3_1 hold2476 (.A(_00890_),
    .X(net7025));
 sg13g2_dlygate4sd3_1 hold2477 (.A(\scanline[37][1] ),
    .X(net7026));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\scanline[42][3] ),
    .X(net7027));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\atari2600.pia.interval[0] ),
    .X(net7028));
 sg13g2_dlygate4sd3_1 hold2480 (.A(_01239_),
    .X(net7029));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\atari2600.ram[11][4] ),
    .X(net7030));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\scanline[56][1] ),
    .X(net7031));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\atari2600.tia.diag[88] ),
    .X(net7032));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\atari2600.ram[15][3] ),
    .X(net7033));
 sg13g2_dlygate4sd3_1 hold2485 (.A(\atari2600.ram[23][7] ),
    .X(net7034));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\scanline[130][6] ),
    .X(net7035));
 sg13g2_dlygate4sd3_1 hold2487 (.A(\atari2600.cpu.IRHOLD[5] ),
    .X(net7036));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\scanline[26][0] ),
    .X(net7037));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\atari2600.tia.colubk[0] ),
    .X(net7038));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\atari2600.cpu.AXYS[0][7] ),
    .X(net7039));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\atari2600.tia.old_grp1[0] ),
    .X(net7040));
 sg13g2_dlygate4sd3_1 hold2492 (.A(_00915_),
    .X(net7041));
 sg13g2_dlygate4sd3_1 hold2493 (.A(\scanline[44][2] ),
    .X(net7042));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\atari2600.ram[111][7] ),
    .X(net7043));
 sg13g2_dlygate4sd3_1 hold2495 (.A(\scanline[146][3] ),
    .X(net7044));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\scanline[5][2] ),
    .X(net7045));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\scanline[96][5] ),
    .X(net7046));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\scanline[44][1] ),
    .X(net7047));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\atari2600.ram[71][7] ),
    .X(net7048));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\atari2600.tia.colupf[6] ),
    .X(net7049));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\atari2600.ram[55][3] ),
    .X(net7050));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\scanline[69][2] ),
    .X(net7051));
 sg13g2_dlygate4sd3_1 hold2503 (.A(\scanline[19][5] ),
    .X(net7052));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\scanline[24][4] ),
    .X(net7053));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\scanline[136][2] ),
    .X(net7054));
 sg13g2_dlygate4sd3_1 hold2506 (.A(\scanline[9][0] ),
    .X(net7055));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\scanline[19][0] ),
    .X(net7056));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\atari2600.ram[55][6] ),
    .X(net7057));
 sg13g2_dlygate4sd3_1 hold2509 (.A(\atari2600.ram[64][7] ),
    .X(net7058));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\atari2600.cpu.ABL[3] ),
    .X(net7059));
 sg13g2_dlygate4sd3_1 hold2511 (.A(_01394_),
    .X(net7060));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\scanline[48][4] ),
    .X(net7061));
 sg13g2_dlygate4sd3_1 hold2513 (.A(\scanline[43][6] ),
    .X(net7062));
 sg13g2_dlygate4sd3_1 hold2514 (.A(\scanline[20][5] ),
    .X(net7063));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\atari2600.ram[35][5] ),
    .X(net7064));
 sg13g2_dlygate4sd3_1 hold2516 (.A(\atari2600.cpu.cond_code[0] ),
    .X(net7065));
 sg13g2_dlygate4sd3_1 hold2517 (.A(\scanline[6][4] ),
    .X(net7066));
 sg13g2_dlygate4sd3_1 hold2518 (.A(\scanline[8][6] ),
    .X(net7067));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\atari2600.cpu.PC[0] ),
    .X(net7068));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\scanline[19][3] ),
    .X(net7069));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\atari2600.ram[11][0] ),
    .X(net7070));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\scanline[9][3] ),
    .X(net7071));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\scanline[112][6] ),
    .X(net7072));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\atari2600.ram[39][0] ),
    .X(net7073));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\scanline[11][5] ),
    .X(net7074));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\rom_last_read_addr[1] ),
    .X(net7075));
 sg13g2_dlygate4sd3_1 hold2527 (.A(_00265_),
    .X(net7076));
 sg13g2_dlygate4sd3_1 hold2528 (.A(\scanline[140][3] ),
    .X(net7077));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\scanline[38][1] ),
    .X(net7078));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\scanline[145][5] ),
    .X(net7079));
 sg13g2_dlygate4sd3_1 hold2531 (.A(\scanline[20][6] ),
    .X(net7080));
 sg13g2_dlygate4sd3_1 hold2532 (.A(\atari2600.tia.refp1 ),
    .X(net7081));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\scanline[74][2] ),
    .X(net7082));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\gamepad_pmod.driver.shift_reg[8] ),
    .X(net7083));
 sg13g2_dlygate4sd3_1 hold2535 (.A(_01484_),
    .X(net7084));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\atari2600.ram[123][1] ),
    .X(net7085));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\scanline[50][0] ),
    .X(net7086));
 sg13g2_dlygate4sd3_1 hold2538 (.A(\atari2600.ram[103][2] ),
    .X(net7087));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\atari2600.ram[44][1] ),
    .X(net7088));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\scanline[26][6] ),
    .X(net7089));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\scanline[145][0] ),
    .X(net7090));
 sg13g2_dlygate4sd3_1 hold2542 (.A(\atari2600.tia.diag[83] ),
    .X(net7091));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\scanline[135][1] ),
    .X(net7092));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\atari2600.ram[91][5] ),
    .X(net7093));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\gamepad_pmod.driver.shift_reg[2] ),
    .X(net7094));
 sg13g2_dlygate4sd3_1 hold2546 (.A(_01478_),
    .X(net7095));
 sg13g2_dlygate4sd3_1 hold2547 (.A(\atari2600.cpu.ABL[0] ),
    .X(net7096));
 sg13g2_dlygate4sd3_1 hold2548 (.A(_01391_),
    .X(net7097));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\scanline[38][5] ),
    .X(net7098));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\atari2600.ram[123][2] ),
    .X(net7099));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\scanline[104][5] ),
    .X(net7100));
 sg13g2_dlygate4sd3_1 hold2552 (.A(\scanline[19][4] ),
    .X(net7101));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\atari2600.cpu.index_y ),
    .X(net7102));
 sg13g2_dlygate4sd3_1 hold2554 (.A(\scanline[11][4] ),
    .X(net7103));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\atari2600.pia.time_counter[20] ),
    .X(net7104));
 sg13g2_dlygate4sd3_1 hold2556 (.A(_05456_),
    .X(net7105));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\scanline[83][0] ),
    .X(net7106));
 sg13g2_dlygate4sd3_1 hold2558 (.A(\atari2600.ram[95][5] ),
    .X(net7107));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\atari2600.pia.diag[3] ),
    .X(net7108));
 sg13g2_dlygate4sd3_1 hold2560 (.A(_00860_),
    .X(net7109));
 sg13g2_dlygate4sd3_1 hold2561 (.A(\scanline[18][2] ),
    .X(net7110));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\atari2600.tia.audv0[1] ),
    .X(net7111));
 sg13g2_dlygate4sd3_1 hold2563 (.A(\atari2600.tia.audv0[2] ),
    .X(net7112));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\rom_last_read_addr[7] ),
    .X(net7113));
 sg13g2_dlygate4sd3_1 hold2565 (.A(_00271_),
    .X(net7114));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\atari2600.cpu.ABL[5] ),
    .X(net7115));
 sg13g2_dlygate4sd3_1 hold2567 (.A(\atari2600.cpu.PC[11] ),
    .X(net7116));
 sg13g2_dlygate4sd3_1 hold2568 (.A(_01421_),
    .X(net7117));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\atari2600.tia.hmm0[0] ),
    .X(net7118));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\atari2600.cpu.Z ),
    .X(net7119));
 sg13g2_dlygate4sd3_1 hold2571 (.A(_01388_),
    .X(net7120));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\atari2600.ram[87][5] ),
    .X(net7121));
 sg13g2_dlygate4sd3_1 hold2573 (.A(\atari2600.tia.poly5_l.x[3] ),
    .X(net7122));
 sg13g2_dlygate4sd3_1 hold2574 (.A(\atari2600.cpu.AXYS[0][1] ),
    .X(net7123));
 sg13g2_dlygate4sd3_1 hold2575 (.A(\atari2600.pia.reset_timer[2] ),
    .X(net7124));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\atari2600.cpu.ABH[5] ),
    .X(net7125));
 sg13g2_dlygate4sd3_1 hold2577 (.A(_01877_),
    .X(net7126));
 sg13g2_dlygate4sd3_1 hold2578 (.A(_00160_),
    .X(net7127));
 sg13g2_dlygate4sd3_1 hold2579 (.A(\atari2600.pia.dat_o[3] ),
    .X(net7128));
 sg13g2_dlygate4sd3_1 hold2580 (.A(_00869_),
    .X(net7129));
 sg13g2_dlygate4sd3_1 hold2581 (.A(\atari2600.tia.diag[86] ),
    .X(net7130));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\hvsync_gen.vga.vpos[9] ),
    .X(net7131));
 sg13g2_dlygate4sd3_1 hold2583 (.A(_01517_),
    .X(net7132));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\scanline[18][0] ),
    .X(net7133));
 sg13g2_dlygate4sd3_1 hold2585 (.A(\scanline[7][4] ),
    .X(net7134));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\scanline[65][5] ),
    .X(net7135));
 sg13g2_dlygate4sd3_1 hold2587 (.A(\atari2600.tia.poly4_l.x[3] ),
    .X(net7136));
 sg13g2_dlygate4sd3_1 hold2588 (.A(_01198_),
    .X(net7137));
 sg13g2_dlygate4sd3_1 hold2589 (.A(\atari2600.pia.reset_timer[1] ),
    .X(net7138));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\atari2600.tia.old_grp1[2] ),
    .X(net7139));
 sg13g2_dlygate4sd3_1 hold2591 (.A(_00917_),
    .X(net7140));
 sg13g2_dlygate4sd3_1 hold2592 (.A(\atari2600.tia.poly5_l.x[4] ),
    .X(net7141));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\scanline[131][5] ),
    .X(net7142));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\atari2600.cpu.DI[7] ),
    .X(net7143));
 sg13g2_dlygate4sd3_1 hold2595 (.A(_01390_),
    .X(net7144));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\atari2600.cpu.PC[6] ),
    .X(net7145));
 sg13g2_dlygate4sd3_1 hold2597 (.A(_01416_),
    .X(net7146));
 sg13g2_dlygate4sd3_1 hold2598 (.A(\gamepad_pmod.driver.shift_reg[7] ),
    .X(net7147));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\atari2600.tia.hmm0[1] ),
    .X(net7148));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\atari2600.tia.diag[99] ),
    .X(net7149));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\atari2600.cpu.ABL[4] ),
    .X(net7150));
 sg13g2_dlygate4sd3_1 hold2602 (.A(_01395_),
    .X(net7151));
 sg13g2_dlygate4sd3_1 hold2603 (.A(\atari2600.tia.hmbl[1] ),
    .X(net7152));
 sg13g2_dlygate4sd3_1 hold2604 (.A(\atari2600.tia.poly9_l.x[3] ),
    .X(net7153));
 sg13g2_dlygate4sd3_1 hold2605 (.A(_01206_),
    .X(net7154));
 sg13g2_dlygate4sd3_1 hold2606 (.A(\atari2600.cpu.ALU.HC ),
    .X(net7155));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\atari2600.tia.diag[90] ),
    .X(net7156));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\atari2600.pia.dat_o[5] ),
    .X(net7157));
 sg13g2_dlygate4sd3_1 hold2609 (.A(_00871_),
    .X(net7158));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\atari2600.pia.diag[5] ),
    .X(net7159));
 sg13g2_dlygate4sd3_1 hold2611 (.A(\atari2600.tia.diag[93] ),
    .X(net7160));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\atari2600.cpu.adc_bcd ),
    .X(net7161));
 sg13g2_dlygate4sd3_1 hold2613 (.A(\atari2600.tia.poly9_l.x[5] ),
    .X(net7162));
 sg13g2_dlygate4sd3_1 hold2614 (.A(_01208_),
    .X(net7163));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\atari2600.cpu.bit_ins ),
    .X(net7164));
 sg13g2_dlygate4sd3_1 hold2616 (.A(\rom_next_addr_in_queue[0] ),
    .X(net7165));
 sg13g2_dlygate4sd3_1 hold2617 (.A(_00284_),
    .X(net7166));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\atari2600.pia.dat_o[4] ),
    .X(net7167));
 sg13g2_dlygate4sd3_1 hold2619 (.A(_00870_),
    .X(net7168));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\atari2600.tia.vblank ),
    .X(net7169));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\atari2600.cpu.adc_sbc ),
    .X(net7170));
 sg13g2_dlygate4sd3_1 hold2622 (.A(\atari2600.ram[71][0] ),
    .X(net7171));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\atari2600.tia.colubk[1] ),
    .X(net7172));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\atari2600.tia.diag[91] ),
    .X(net7173));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\atari2600.tia.colupf[1] ),
    .X(net7174));
 sg13g2_dlygate4sd3_1 hold2626 (.A(\atari2600.cpu.PC[12] ),
    .X(net7175));
 sg13g2_dlygate4sd3_1 hold2627 (.A(_01422_),
    .X(net7176));
 sg13g2_dlygate4sd3_1 hold2628 (.A(\scanline[19][2] ),
    .X(net7177));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\hvsync_gen.vga.vpos[5] ),
    .X(net7178));
 sg13g2_dlygate4sd3_1 hold2630 (.A(_07869_),
    .X(net7179));
 sg13g2_dlygate4sd3_1 hold2631 (.A(_01513_),
    .X(net7180));
 sg13g2_dlygate4sd3_1 hold2632 (.A(\atari2600.cpu.IRHOLD[2] ),
    .X(net7181));
 sg13g2_dlygate4sd3_1 hold2633 (.A(_01378_),
    .X(net7182));
 sg13g2_dlygate4sd3_1 hold2634 (.A(\atari2600.cpu.ABL[6] ),
    .X(net7183));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\atari2600.pia.time_counter[3] ),
    .X(net7184));
 sg13g2_dlygate4sd3_1 hold2636 (.A(_05414_),
    .X(net7185));
 sg13g2_dlygate4sd3_1 hold2637 (.A(\scanline[129][4] ),
    .X(net7186));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\atari2600.cpu.IRHOLD[3] ),
    .X(net7187));
 sg13g2_dlygate4sd3_1 hold2639 (.A(_01379_),
    .X(net7188));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\atari2600.ram[67][2] ),
    .X(net7189));
 sg13g2_dlygate4sd3_1 hold2641 (.A(\atari2600.tia.diag[94] ),
    .X(net7190));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\atari2600.cpu.I ),
    .X(net7191));
 sg13g2_dlygate4sd3_1 hold2643 (.A(_01385_),
    .X(net7192));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\atari2600.tia.audf0[4] ),
    .X(net7193));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\flash_rom.addr_in[18] ),
    .X(net7194));
 sg13g2_dlygate4sd3_1 hold2646 (.A(_00965_),
    .X(net7195));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\atari2600.cpu.PC[7] ),
    .X(net7196));
 sg13g2_dlygate4sd3_1 hold2648 (.A(_01417_),
    .X(net7197));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\atari2600.tia.diag[84] ),
    .X(net7198));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\scanline[116][1] ),
    .X(net7199));
 sg13g2_dlygate4sd3_1 hold2651 (.A(\atari2600.input_switches[2] ),
    .X(net7200));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\atari2600.tia.poly5_r.x[2] ),
    .X(net7201));
 sg13g2_dlygate4sd3_1 hold2653 (.A(_01218_),
    .X(net7202));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\atari2600.pia.time_counter[9] ),
    .X(net7203));
 sg13g2_dlygate4sd3_1 hold2655 (.A(\gamepad_pmod.decoder.data_reg[1] ),
    .X(net7204));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\atari2600.tia.poly9_r.x[5] ),
    .X(net7205));
 sg13g2_dlygate4sd3_1 hold2657 (.A(_01226_),
    .X(net7206));
 sg13g2_dlygate4sd3_1 hold2658 (.A(\atari2600.pia.time_counter[12] ),
    .X(net7207));
 sg13g2_dlygate4sd3_1 hold2659 (.A(_05439_),
    .X(net7208));
 sg13g2_dlygate4sd3_1 hold2660 (.A(\atari2600.tia.poly9_l.x[4] ),
    .X(net7209));
 sg13g2_dlygate4sd3_1 hold2661 (.A(\atari2600.tia.colubk[6] ),
    .X(net7210));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\atari2600.tia.diag[81] ),
    .X(net7211));
 sg13g2_dlygate4sd3_1 hold2663 (.A(\atari2600.cpu.clv ),
    .X(net7212));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\atari2600.tia.diag[76] ),
    .X(net7213));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\atari2600.cpu.PC[13] ),
    .X(net7214));
 sg13g2_dlygate4sd3_1 hold2666 (.A(_01423_),
    .X(net7215));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\atari2600.ram[123][0] ),
    .X(net7216));
 sg13g2_dlygate4sd3_1 hold2668 (.A(\atari2600.cpu.IRHOLD[7] ),
    .X(net7217));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\atari2600.cpu.V ),
    .X(net7218));
 sg13g2_dlygate4sd3_1 hold2670 (.A(_01386_),
    .X(net7219));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\atari2600.tia.colupf[2] ),
    .X(net7220));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\atari2600.tia.diag[78] ),
    .X(net7221));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\atari2600.tia.colubk[5] ),
    .X(net7222));
 sg13g2_dlygate4sd3_1 hold2674 (.A(\rom_next_addr_in_queue[1] ),
    .X(net7223));
 sg13g2_dlygate4sd3_1 hold2675 (.A(_00285_),
    .X(net7224));
 sg13g2_dlygate4sd3_1 hold2676 (.A(\atari2600.tia.poly9_l.x[1] ),
    .X(net7225));
 sg13g2_dlygate4sd3_1 hold2677 (.A(_01204_),
    .X(net7226));
 sg13g2_dlygate4sd3_1 hold2678 (.A(\gamepad_pmod.driver.shift_reg[9] ),
    .X(net7227));
 sg13g2_dlygate4sd3_1 hold2679 (.A(_01485_),
    .X(net7228));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\atari2600.tia.diag[89] ),
    .X(net7229));
 sg13g2_dlygate4sd3_1 hold2681 (.A(\scanline[4][2] ),
    .X(net7230));
 sg13g2_dlygate4sd3_1 hold2682 (.A(\gamepad_pmod.driver.shift_reg[3] ),
    .X(net7231));
 sg13g2_dlygate4sd3_1 hold2683 (.A(_01479_),
    .X(net7232));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\rom_last_read_addr[0] ),
    .X(net7233));
 sg13g2_dlygate4sd3_1 hold2685 (.A(\atari2600.input_switches[1] ),
    .X(net7234));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\atari2600.tia.diag[79] ),
    .X(net7235));
 sg13g2_dlygate4sd3_1 hold2687 (.A(\flash_rom.addr[16] ),
    .X(net7236));
 sg13g2_dlygate4sd3_1 hold2688 (.A(_00979_),
    .X(net7237));
 sg13g2_dlygate4sd3_1 hold2689 (.A(\atari2600.cpu.shift_right ),
    .X(net7238));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\hvsync_gen.vga.vpos[8] ),
    .X(net7239));
 sg13g2_dlygate4sd3_1 hold2691 (.A(_07874_),
    .X(net7240));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\atari2600.cpu.PC[5] ),
    .X(net7241));
 sg13g2_dlygate4sd3_1 hold2693 (.A(_01415_),
    .X(net7242));
 sg13g2_dlygate4sd3_1 hold2694 (.A(\atari2600.pia.reset_timer[0] ),
    .X(net7243));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\atari2600.tia.poly4_r.x[2] ),
    .X(net7244));
 sg13g2_dlygate4sd3_1 hold2696 (.A(_01214_),
    .X(net7245));
 sg13g2_dlygate4sd3_1 hold2697 (.A(\rom_last_read_addr[6] ),
    .X(net7246));
 sg13g2_dlygate4sd3_1 hold2698 (.A(_00270_),
    .X(net7247));
 sg13g2_dlygate4sd3_1 hold2699 (.A(\atari2600.cpu.ABL[1] ),
    .X(net7248));
 sg13g2_dlygate4sd3_1 hold2700 (.A(_01392_),
    .X(net7249));
 sg13g2_dlygate4sd3_1 hold2701 (.A(\atari2600.cpu.IRHOLD[6] ),
    .X(net7250));
 sg13g2_dlygate4sd3_1 hold2702 (.A(_01382_),
    .X(net7251));
 sg13g2_dlygate4sd3_1 hold2703 (.A(\atari2600.tia.p9_l ),
    .X(net7252));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\atari2600.cpu.PC[3] ),
    .X(net7253));
 sg13g2_dlygate4sd3_1 hold2705 (.A(_00059_),
    .X(net7254));
 sg13g2_dlygate4sd3_1 hold2706 (.A(_01887_),
    .X(net7255));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\atari2600.tia.diag[82] ),
    .X(net7256));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\atari2600.tia.poly9_r.x[1] ),
    .X(net7257));
 sg13g2_dlygate4sd3_1 hold2709 (.A(_01222_),
    .X(net7258));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\atari2600.ram_data[5] ),
    .X(net7259));
 sg13g2_dlygate4sd3_1 hold2711 (.A(_07402_),
    .X(net7260));
 sg13g2_dlygate4sd3_1 hold2712 (.A(\atari2600.cpu.PC[9] ),
    .X(net7261));
 sg13g2_dlygate4sd3_1 hold2713 (.A(_01419_),
    .X(net7262));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\atari2600.tia.diag[100] ),
    .X(net7263));
 sg13g2_dlygate4sd3_1 hold2715 (.A(\atari2600.tia.colubk[4] ),
    .X(net7264));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\atari2600.tia.diag[92] ),
    .X(net7265));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\atari2600.cpu.IRHOLD[1] ),
    .X(net7266));
 sg13g2_dlygate4sd3_1 hold2718 (.A(\atari2600.cpu.DI[3] ),
    .X(net7267));
 sg13g2_dlygate4sd3_1 hold2719 (.A(\atari2600.cpu.DIMUX[3] ),
    .X(net7268));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\atari2600.ram_data[4] ),
    .X(net7269));
 sg13g2_dlygate4sd3_1 hold2721 (.A(\atari2600.pia.diag[0] ),
    .X(net7270));
 sg13g2_dlygate4sd3_1 hold2722 (.A(_00857_),
    .X(net7271));
 sg13g2_dlygate4sd3_1 hold2723 (.A(\atari2600.tia.poly9_l.x[2] ),
    .X(net7272));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\atari2600.tia.diag[95] ),
    .X(net7273));
 sg13g2_dlygate4sd3_1 hold2725 (.A(\atari2600.pia.diag[4] ),
    .X(net7274));
 sg13g2_dlygate4sd3_1 hold2726 (.A(_00861_),
    .X(net7275));
 sg13g2_dlygate4sd3_1 hold2727 (.A(\atari2600.pia.diag[1] ),
    .X(net7276));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\atari2600.pia.diag[6] ),
    .X(net7277));
 sg13g2_dlygate4sd3_1 hold2729 (.A(_00863_),
    .X(net7278));
 sg13g2_dlygate4sd3_1 hold2730 (.A(\atari2600.tia.audv0[0] ),
    .X(net7279));
 sg13g2_dlygate4sd3_1 hold2731 (.A(\atari2600.cpu.inc ),
    .X(net7280));
 sg13g2_dlygate4sd3_1 hold2732 (.A(\rom_next_addr_in_queue[4] ),
    .X(net7281));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\atari2600.tia.diag[77] ),
    .X(net7282));
 sg13g2_dlygate4sd3_1 hold2734 (.A(\atari2600.pia.diag[7] ),
    .X(net7283));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\atari2600.tia.hmbl[2] ),
    .X(net7284));
 sg13g2_dlygate4sd3_1 hold2736 (.A(\atari2600.input_switches[0] ),
    .X(net7285));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\atari2600.tia.colubk[2] ),
    .X(net7286));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\atari2600.tia.colubk[3] ),
    .X(net7287));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\atari2600.tia.colup1[4] ),
    .X(net7288));
 sg13g2_dlygate4sd3_1 hold2740 (.A(\atari2600.tia.diag[98] ),
    .X(net7289));
 sg13g2_dlygate4sd3_1 hold2741 (.A(\atari2600.cpu.load_only ),
    .X(net7290));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\atari2600.tia.diag[87] ),
    .X(net7291));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\atari2600.cpu.cond_code[2] ),
    .X(net7292));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\atari2600.tia.colup1[0] ),
    .X(net7293));
 sg13g2_dlygate4sd3_1 hold2745 (.A(\atari2600.pia.time_counter[2] ),
    .X(net7294));
 sg13g2_dlygate4sd3_1 hold2746 (.A(\atari2600.tia.hmm0[2] ),
    .X(net7295));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\atari2600.cpu.rotate ),
    .X(net7296));
 sg13g2_dlygate4sd3_1 hold2748 (.A(uio_oe[1]),
    .X(net7297));
 sg13g2_dlygate4sd3_1 hold2749 (.A(_01824_),
    .X(net7298));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\atari2600.cpu.DI[6] ),
    .X(net7299));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\atari2600.cpu.DIMUX[6] ),
    .X(net7300));
 sg13g2_dlygate4sd3_1 hold2752 (.A(\atari2600.tia.diag[110] ),
    .X(net7301));
 sg13g2_dlygate4sd3_1 hold2753 (.A(\atari2600.tia.colupf[0] ),
    .X(net7302));
 sg13g2_dlygate4sd3_1 hold2754 (.A(_00094_),
    .X(net7303));
 sg13g2_dlygate4sd3_1 hold2755 (.A(_11057_),
    .X(net7304));
 sg13g2_dlygate4sd3_1 hold2756 (.A(_01825_),
    .X(net7305));
 sg13g2_dlygate4sd3_1 hold2757 (.A(\atari2600.tia.audio_left_counter[1] ),
    .X(net7306));
 sg13g2_dlygate4sd3_1 hold2758 (.A(_00992_),
    .X(net7307));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\atari2600.pia.time_counter[23] ),
    .X(net7308));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\atari2600.tia.audio_right_counter[1] ),
    .X(net7309));
 sg13g2_dlygate4sd3_1 hold2761 (.A(_01008_),
    .X(net7310));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\atari2600.cpu.DIHOLD[2] ),
    .X(net7311));
 sg13g2_dlygate4sd3_1 hold2763 (.A(\atari2600.cpu.DIMUX[2] ),
    .X(net7312));
 sg13g2_dlygate4sd3_1 hold2764 (.A(\atari2600.pia.diag[2] ),
    .X(net7313));
 sg13g2_dlygate4sd3_1 hold2765 (.A(_00859_),
    .X(net7314));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\atari2600.tia.enabl ),
    .X(net7315));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\rom_next_addr_in_queue[8] ),
    .X(net7316));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\atari2600.tia.diag[85] ),
    .X(net7317));
 sg13g2_dlygate4sd3_1 hold2769 (.A(\atari2600.tia.p0_spacing[6] ),
    .X(net7318));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\atari2600.tia.colupf[5] ),
    .X(net7319));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\atari2600.tia.diag[109] ),
    .X(net7320));
 sg13g2_dlygate4sd3_1 hold2772 (.A(\hvsync_gen.vga.vpos[1] ),
    .X(net7321));
 sg13g2_dlygate4sd3_1 hold2773 (.A(_01509_),
    .X(net7322));
 sg13g2_dlygate4sd3_1 hold2774 (.A(\rom_next_addr_in_queue[10] ),
    .X(net7323));
 sg13g2_dlygate4sd3_1 hold2775 (.A(_00294_),
    .X(net7324));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\atari2600.tia.p4_r ),
    .X(net7325));
 sg13g2_dlygate4sd3_1 hold2777 (.A(_01213_),
    .X(net7326));
 sg13g2_dlygate4sd3_1 hold2778 (.A(\atari2600.pia.dat_o[0] ),
    .X(net7327));
 sg13g2_dlygate4sd3_1 hold2779 (.A(_07378_),
    .X(net7328));
 sg13g2_dlygate4sd3_1 hold2780 (.A(\rom_last_read_addr[9] ),
    .X(net7329));
 sg13g2_dlygate4sd3_1 hold2781 (.A(_00273_),
    .X(net7330));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\atari2600.tia.audv1[0] ),
    .X(net7331));
 sg13g2_dlygate4sd3_1 hold2783 (.A(\atari2600.tia.diag[96] ),
    .X(net7332));
 sg13g2_dlygate4sd3_1 hold2784 (.A(\atari2600.tia.audv0[3] ),
    .X(net7333));
 sg13g2_dlygate4sd3_1 hold2785 (.A(\atari2600.tia.colup1[6] ),
    .X(net7334));
 sg13g2_dlygate4sd3_1 hold2786 (.A(\atari2600.tia.p1_spacing[5] ),
    .X(net7335));
 sg13g2_dlygate4sd3_1 hold2787 (.A(\rom_next_addr_in_queue[5] ),
    .X(net7336));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\atari2600.pia.time_counter[7] ),
    .X(net7337));
 sg13g2_dlygate4sd3_1 hold2789 (.A(_05424_),
    .X(net7338));
 sg13g2_dlygate4sd3_1 hold2790 (.A(_00881_),
    .X(net7339));
 sg13g2_dlygate4sd3_1 hold2791 (.A(\atari2600.ram_data[3] ),
    .X(net7340));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\atari2600.tia.colupf[3] ),
    .X(net7341));
 sg13g2_dlygate4sd3_1 hold2793 (.A(\atari2600.tia.audv1[3] ),
    .X(net7342));
 sg13g2_dlygate4sd3_1 hold2794 (.A(\atari2600.pia.time_counter[6] ),
    .X(net7343));
 sg13g2_dlygate4sd3_1 hold2795 (.A(_05423_),
    .X(net7344));
 sg13g2_dlygate4sd3_1 hold2796 (.A(\atari2600.input_switches[3] ),
    .X(net7345));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\atari2600.ram_data[2] ),
    .X(net7346));
 sg13g2_dlygate4sd3_1 hold2798 (.A(_07387_),
    .X(net7347));
 sg13g2_dlygate4sd3_1 hold2799 (.A(\atari2600.pia.time_counter[1] ),
    .X(net7348));
 sg13g2_dlygate4sd3_1 hold2800 (.A(_05411_),
    .X(net7349));
 sg13g2_dlygate4sd3_1 hold2801 (.A(\rom_next_addr_in_queue[9] ),
    .X(net7350));
 sg13g2_dlygate4sd3_1 hold2802 (.A(_00156_),
    .X(net7351));
 sg13g2_dlygate4sd3_1 hold2803 (.A(_01007_),
    .X(net7352));
 sg13g2_dlygate4sd3_1 hold2804 (.A(\atari2600.pia.time_counter[19] ),
    .X(net7353));
 sg13g2_dlygate4sd3_1 hold2805 (.A(_05455_),
    .X(net7354));
 sg13g2_dlygate4sd3_1 hold2806 (.A(\atari2600.tia.colup1[1] ),
    .X(net7355));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\atari2600.cpu.ABH[4] ),
    .X(net7356));
 sg13g2_dlygate4sd3_1 hold2808 (.A(\r_pwm_odd[1] ),
    .X(net7357));
 sg13g2_dlygate4sd3_1 hold2809 (.A(_04543_),
    .X(net7358));
 sg13g2_dlygate4sd3_1 hold2810 (.A(_00330_),
    .X(net7359));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\atari2600.tia.diag[106] ),
    .X(net7360));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\atari2600.tia.p1_spacing[6] ),
    .X(net7361));
 sg13g2_dlygate4sd3_1 hold2813 (.A(\flash_rom.stall_read ),
    .X(net7362));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\atari2600.tia.colup1[2] ),
    .X(net7363));
 sg13g2_dlygate4sd3_1 hold2815 (.A(\atari2600.tia.diag[104] ),
    .X(net7364));
 sg13g2_dlygate4sd3_1 hold2816 (.A(\rom_next_addr_in_queue[3] ),
    .X(net7365));
 sg13g2_dlygate4sd3_1 hold2817 (.A(\atari2600.ram_data[1] ),
    .X(net7366));
 sg13g2_dlygate4sd3_1 hold2818 (.A(_07382_),
    .X(net7367));
 sg13g2_dlygate4sd3_1 hold2819 (.A(\atari2600.tia.p1_spacing[4] ),
    .X(net7368));
 sg13g2_dlygate4sd3_1 hold2820 (.A(\rom_next_addr_in_queue[2] ),
    .X(net7369));
 sg13g2_dlygate4sd3_1 hold2821 (.A(\atari2600.tia.diag[111] ),
    .X(net7370));
 sg13g2_dlygate4sd3_1 hold2822 (.A(\atari2600.tia.diag[105] ),
    .X(net7371));
 sg13g2_dlygate4sd3_1 hold2823 (.A(\atari2600.tia.poly4_l.x[1] ),
    .X(net7372));
 sg13g2_dlygate4sd3_1 hold2824 (.A(_01195_),
    .X(net7373));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\audio_pwm_accumulator[0] ),
    .X(net7374));
 sg13g2_dlygate4sd3_1 hold2826 (.A(_00296_),
    .X(net7375));
 sg13g2_dlygate4sd3_1 hold2827 (.A(\atari2600.cpu.op[0] ),
    .X(net7376));
 sg13g2_dlygate4sd3_1 hold2828 (.A(\atari2600.tia.hmm1[1] ),
    .X(net7377));
 sg13g2_dlygate4sd3_1 hold2829 (.A(\atari2600.tia.audv1[1] ),
    .X(net7378));
 sg13g2_dlygate4sd3_1 hold2830 (.A(\flash_rom.addr[7] ),
    .X(net7379));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\atari2600.tia.colup1[5] ),
    .X(net7380));
 sg13g2_dlygate4sd3_1 hold2832 (.A(\atari2600.cpu.PC[15] ),
    .X(net7381));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\atari2600.tia.diag[108] ),
    .X(net7382));
 sg13g2_dlygate4sd3_1 hold2834 (.A(\atari2600.tia.hmbl[0] ),
    .X(net7383));
 sg13g2_dlygate4sd3_1 hold2835 (.A(_00130_),
    .X(net7384));
 sg13g2_dlygate4sd3_1 hold2836 (.A(\atari2600.tia.colup0[2] ),
    .X(net7385));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\atari2600.cpu.dst_reg[1] ),
    .X(net7386));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\atari2600.tia.colupf[4] ),
    .X(net7387));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\atari2600.tia.audv1[2] ),
    .X(net7388));
 sg13g2_dlygate4sd3_1 hold2840 (.A(\atari2600.tia.colup0[4] ),
    .X(net7389));
 sg13g2_dlygate4sd3_1 hold2841 (.A(\atari2600.tia.diag[107] ),
    .X(net7390));
 sg13g2_dlygate4sd3_1 hold2842 (.A(\atari2600.pia.time_counter[18] ),
    .X(net7391));
 sg13g2_dlygate4sd3_1 hold2843 (.A(_05453_),
    .X(net7392));
 sg13g2_dlygate4sd3_1 hold2844 (.A(\flash_rom.nibbles_remaining[0] ),
    .X(net7393));
 sg13g2_dlygate4sd3_1 hold2845 (.A(_01809_),
    .X(net7394));
 sg13g2_dlygate4sd3_1 hold2846 (.A(\atari2600.cpu.cond_code[1] ),
    .X(net7395));
 sg13g2_dlygate4sd3_1 hold2847 (.A(\atari2600.tia.hmm1[0] ),
    .X(net7396));
 sg13g2_dlygate4sd3_1 hold2848 (.A(\atari2600.tia.hmp1[0] ),
    .X(net7397));
 sg13g2_dlygate4sd3_1 hold2849 (.A(\atari2600.cpu.ABH[2] ),
    .X(net7398));
 sg13g2_dlygate4sd3_1 hold2850 (.A(\atari2600.cpu.ABH[1] ),
    .X(net7399));
 sg13g2_dlygate4sd3_1 hold2851 (.A(\atari2600.pia.underflow ),
    .X(net7400));
 sg13g2_dlygate4sd3_1 hold2852 (.A(\flash_rom.addr[5] ),
    .X(net7401));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\external_rom_data[1] ),
    .X(net7402));
 sg13g2_dlygate4sd3_1 hold2854 (.A(_01816_),
    .X(net7403));
 sg13g2_dlygate4sd3_1 hold2855 (.A(\atari2600.tia.ball_w[0] ),
    .X(net7404));
 sg13g2_dlygate4sd3_1 hold2856 (.A(\atari2600.pia.time_counter[0] ),
    .X(net7405));
 sg13g2_dlygate4sd3_1 hold2857 (.A(\rom_next_addr_in_queue[11] ),
    .X(net7406));
 sg13g2_dlygate4sd3_1 hold2858 (.A(\atari2600.cpu.dst_reg[0] ),
    .X(net7407));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\atari2600.tia.enam0 ),
    .X(net7408));
 sg13g2_dlygate4sd3_1 hold2860 (.A(\atari2600.tia.ball_w[3] ),
    .X(net7409));
 sg13g2_dlygate4sd3_1 hold2861 (.A(\atari2600.tia.hmp0[0] ),
    .X(net7410));
 sg13g2_dlygate4sd3_1 hold2862 (.A(\atari2600.tia.ball_w[1] ),
    .X(net7411));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\hvsync_gen.vga.vpos[2] ),
    .X(net7412));
 sg13g2_dlygate4sd3_1 hold2864 (.A(\atari2600.cpu.PC[14] ),
    .X(net7413));
 sg13g2_dlygate4sd3_1 hold2865 (.A(\atari2600.pia.time_counter[4] ),
    .X(net7414));
 sg13g2_dlygate4sd3_1 hold2866 (.A(_05417_),
    .X(net7415));
 sg13g2_dlygate4sd3_1 hold2867 (.A(\atari2600.tia.p0_spacing[5] ),
    .X(net7416));
 sg13g2_dlygate4sd3_1 hold2868 (.A(\atari2600.tia.hmp1[1] ),
    .X(net7417));
 sg13g2_dlygate4sd3_1 hold2869 (.A(\flash_rom.addr[4] ),
    .X(net7418));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\atari2600.tia.hmbl[3] ),
    .X(net7419));
 sg13g2_dlygate4sd3_1 hold2871 (.A(\atari2600.cpu.op[1] ),
    .X(net7420));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\atari2600.tia.diag[61] ),
    .X(net7421));
 sg13g2_dlygate4sd3_1 hold2873 (.A(\rom_next_addr_in_queue[7] ),
    .X(net7422));
 sg13g2_dlygate4sd3_1 hold2874 (.A(_00291_),
    .X(net7423));
 sg13g2_dlygate4sd3_1 hold2875 (.A(\flash_rom.addr[6] ),
    .X(net7424));
 sg13g2_dlygate4sd3_1 hold2876 (.A(\atari2600.cpu.ABH[3] ),
    .X(net7425));
 sg13g2_dlygate4sd3_1 hold2877 (.A(\atari2600.tia.audc0[0] ),
    .X(net7426));
 sg13g2_dlygate4sd3_1 hold2878 (.A(\atari2600.tia.hmp0[2] ),
    .X(net7427));
 sg13g2_dlygate4sd3_1 hold2879 (.A(_00112_),
    .X(net7428));
 sg13g2_dlygate4sd3_1 hold2880 (.A(_08136_),
    .X(net7429));
 sg13g2_dlygate4sd3_1 hold2881 (.A(\atari2600.tia.ball_w[2] ),
    .X(net7430));
 sg13g2_dlygate4sd3_1 hold2882 (.A(\atari2600.cpu.ABH[0] ),
    .X(net7431));
 sg13g2_dlygate4sd3_1 hold2883 (.A(\atari2600.tia.hmp0[3] ),
    .X(net7432));
 sg13g2_dlygate4sd3_1 hold2884 (.A(\hvsync_gen.vga.vpos[6] ),
    .X(net7433));
 sg13g2_dlygate4sd3_1 hold2885 (.A(_07871_),
    .X(net7434));
 sg13g2_dlygate4sd3_1 hold2886 (.A(\atari2600.tia.colup0[3] ),
    .X(net7435));
 sg13g2_dlygate4sd3_1 hold2887 (.A(\atari2600.tia.colup1[3] ),
    .X(net7436));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\hvsync_gen.vga.vpos[7] ),
    .X(net7437));
 sg13g2_dlygate4sd3_1 hold2889 (.A(\atari2600.cpu.op[2] ),
    .X(net7438));
 sg13g2_dlygate4sd3_1 hold2890 (.A(\atari2600.tia.colup0[1] ),
    .X(net7439));
 sg13g2_dlygate4sd3_1 hold2891 (.A(\atari2600.tia.p0_spacing[4] ),
    .X(net7440));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\atari2600.tia.hmp1[2] ),
    .X(net7441));
 sg13g2_dlygate4sd3_1 hold2893 (.A(\hvsync_gen.vga.vpos[4] ),
    .X(net7442));
 sg13g2_dlygate4sd3_1 hold2894 (.A(\atari2600.tia.colup0[0] ),
    .X(net7443));
 sg13g2_dlygate4sd3_1 hold2895 (.A(\flash_rom.nibbles_remaining[2] ),
    .X(net7444));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\atari2600.tia.hmm1[2] ),
    .X(net7445));
 sg13g2_dlygate4sd3_1 hold2897 (.A(\atari2600.cpu.compare ),
    .X(net7446));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\atari2600.clk_counter[0] ),
    .X(net7447));
 sg13g2_dlygate4sd3_1 hold2899 (.A(\flash_rom.addr[11] ),
    .X(net7448));
 sg13g2_dlygate4sd3_1 hold2900 (.A(\atari2600.tia.hmp0[1] ),
    .X(net7449));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\r_pwm_even[1] ),
    .X(net7450));
 sg13g2_dlygate4sd3_1 hold2902 (.A(_04542_),
    .X(net7451));
 sg13g2_dlygate4sd3_1 hold2903 (.A(\atari2600.pia.interval[3] ),
    .X(net7452));
 sg13g2_dlygate4sd3_1 hold2904 (.A(\atari2600.tia.colup0[6] ),
    .X(net7453));
 sg13g2_dlygate4sd3_1 hold2905 (.A(\atari2600.cpu.php ),
    .X(net7454));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\atari2600.cpu.op[3] ),
    .X(net7455));
 sg13g2_dlygate4sd3_1 hold2907 (.A(\hvsync_gen.vga.vpos[3] ),
    .X(net7456));
 sg13g2_dlygate4sd3_1 hold2908 (.A(\atari2600.tia.colup0[5] ),
    .X(net7457));
 sg13g2_dlygate4sd3_1 hold2909 (.A(\atari2600.tia.p0_w[4] ),
    .X(net7458));
 sg13g2_dlygate4sd3_1 hold2910 (.A(\atari2600.tia.diag[44] ),
    .X(net7459));
 sg13g2_dlygate4sd3_1 hold2911 (.A(\atari2600.tia.p1_w[4] ),
    .X(net7460));
 sg13g2_dlygate4sd3_1 hold2912 (.A(\atari2600.tia.audio_l ),
    .X(net7461));
 sg13g2_dlygate4sd3_1 hold2913 (.A(_01023_),
    .X(net7462));
 sg13g2_dlygate4sd3_1 hold2914 (.A(\atari2600.tia.audc1[2] ),
    .X(net7463));
 sg13g2_dlygate4sd3_1 hold2915 (.A(\atari2600.cpu.store ),
    .X(net7464));
 sg13g2_dlygate4sd3_1 hold2916 (.A(_01371_),
    .X(net7465));
 sg13g2_dlygate4sd3_1 hold2917 (.A(\atari2600.tia.diag[39] ),
    .X(net7466));
 sg13g2_dlygate4sd3_1 hold2918 (.A(\atari2600.tia.audf0[3] ),
    .X(net7467));
 sg13g2_dlygate4sd3_1 hold2919 (.A(\hvsync_gen.hpos[1] ),
    .X(net7468));
 sg13g2_dlygate4sd3_1 hold2920 (.A(_03200_),
    .X(net7469));
 sg13g2_dlygate4sd3_1 hold2921 (.A(_00263_),
    .X(net7470));
 sg13g2_dlygate4sd3_1 hold2922 (.A(\atari2600.tia.p0_scale[0] ),
    .X(net7471));
 sg13g2_dlygate4sd3_1 hold2923 (.A(\atari2600.tia.audc1[3] ),
    .X(net7472));
 sg13g2_dlygate4sd3_1 hold2924 (.A(\atari2600.ram_data[7] ),
    .X(net7473));
 sg13g2_dlygate4sd3_1 hold2925 (.A(_01348_),
    .X(net7474));
 sg13g2_dlygate4sd3_1 hold2926 (.A(\flash_rom.nibbles_remaining[1] ),
    .X(net7475));
 sg13g2_dlygate4sd3_1 hold2927 (.A(_01810_),
    .X(net7476));
 sg13g2_dlygate4sd3_1 hold2928 (.A(\atari2600.cpu.shift ),
    .X(net7477));
 sg13g2_dlygate4sd3_1 hold2929 (.A(\rom_next_addr_in_queue[6] ),
    .X(net7478));
 sg13g2_dlygate4sd3_1 hold2930 (.A(\atari2600.tia.p0_w[5] ),
    .X(net7479));
 sg13g2_dlygate4sd3_1 hold2931 (.A(\atari2600.cpu.ADD[3] ),
    .X(net7480));
 sg13g2_dlygate4sd3_1 hold2932 (.A(\atari2600.tia.diag[64] ),
    .X(net7481));
 sg13g2_dlygate4sd3_1 hold2933 (.A(_01100_),
    .X(net7482));
 sg13g2_dlygate4sd3_1 hold2934 (.A(\atari2600.tia.enam1 ),
    .X(net7483));
 sg13g2_dlygate4sd3_1 hold2935 (.A(\flash_rom.addr[10] ),
    .X(net7484));
 sg13g2_dlygate4sd3_1 hold2936 (.A(\atari2600.tia.diag[38] ),
    .X(net7485));
 sg13g2_dlygate4sd3_1 hold2937 (.A(\atari2600.tia.poly9_r.x[6] ),
    .X(net7486));
 sg13g2_dlygate4sd3_1 hold2938 (.A(\atari2600.pia.time_counter[11] ),
    .X(net7487));
 sg13g2_dlygate4sd3_1 hold2939 (.A(\atari2600.tia.hmp1[3] ),
    .X(net7488));
 sg13g2_dlygate4sd3_1 hold2940 (.A(\atari2600.tia.p0_scale[1] ),
    .X(net7489));
 sg13g2_dlygate4sd3_1 hold2941 (.A(\atari2600.pia.time_counter[14] ),
    .X(net7490));
 sg13g2_dlygate4sd3_1 hold2942 (.A(_05443_),
    .X(net7491));
 sg13g2_dlygate4sd3_1 hold2943 (.A(\atari2600.tia.diag[47] ),
    .X(net7492));
 sg13g2_dlygate4sd3_1 hold2944 (.A(_01131_),
    .X(net7493));
 sg13g2_dlygate4sd3_1 hold2945 (.A(\atari2600.tia.diag[46] ),
    .X(net7494));
 sg13g2_dlygate4sd3_1 hold2946 (.A(\flash_rom.spi_clk_out ),
    .X(net7495));
 sg13g2_dlygate4sd3_1 hold2947 (.A(\atari2600.tia.poly9_r.x[7] ),
    .X(net7496));
 sg13g2_dlygate4sd3_1 hold2948 (.A(\flash_rom.addr[8] ),
    .X(net7497));
 sg13g2_dlygate4sd3_1 hold2949 (.A(\atari2600.tia.poly9_r.x[2] ),
    .X(net7498));
 sg13g2_dlygate4sd3_1 hold2950 (.A(\atari2600.tia.diag[48] ),
    .X(net7499));
 sg13g2_dlygate4sd3_1 hold2951 (.A(\atari2600.tia.audf1[1] ),
    .X(net7500));
 sg13g2_dlygate4sd3_1 hold2952 (.A(\atari2600.cpu.ADD[7] ),
    .X(net7501));
 sg13g2_dlygate4sd3_1 hold2953 (.A(\atari2600.tia.diag[54] ),
    .X(net7502));
 sg13g2_dlygate4sd3_1 hold2954 (.A(\atari2600.tia.audf0[1] ),
    .X(net7503));
 sg13g2_dlygate4sd3_1 hold2955 (.A(\atari2600.cpu.ADD[1] ),
    .X(net7504));
 sg13g2_dlygate4sd3_1 hold2956 (.A(\atari2600.tia.diag[55] ),
    .X(net7505));
 sg13g2_dlygate4sd3_1 hold2957 (.A(\atari2600.tia.hmm1[3] ),
    .X(net7506));
 sg13g2_dlygate4sd3_1 hold2958 (.A(\atari2600.tia.diag[51] ),
    .X(net7507));
 sg13g2_dlygate4sd3_1 hold2959 (.A(\atari2600.tia.diag[43] ),
    .X(net7508));
 sg13g2_dlygate4sd3_1 hold2960 (.A(\flash_rom.fsm_state[1] ),
    .X(net7509));
 sg13g2_dlygate4sd3_1 hold2961 (.A(\atari2600.tia.diag[52] ),
    .X(net7510));
 sg13g2_dlygate4sd3_1 hold2962 (.A(_01120_),
    .X(net7511));
 sg13g2_dlygate4sd3_1 hold2963 (.A(_00069_),
    .X(net7512));
 sg13g2_dlygate4sd3_1 hold2964 (.A(_04612_),
    .X(net7513));
 sg13g2_dlygate4sd3_1 hold2965 (.A(_04615_),
    .X(net7514));
 sg13g2_dlygate4sd3_1 hold2966 (.A(\atari2600.tia.p1_w[5] ),
    .X(net7515));
 sg13g2_dlygate4sd3_1 hold2967 (.A(_00081_),
    .X(net7516));
 sg13g2_dlygate4sd3_1 hold2968 (.A(_08731_),
    .X(net7517));
 sg13g2_dlygate4sd3_1 hold2969 (.A(_01389_),
    .X(net7518));
 sg13g2_dlygate4sd3_1 hold2970 (.A(\atari2600.tia.diag[34] ),
    .X(net7519));
 sg13g2_dlygate4sd3_1 hold2971 (.A(\atari2600.tia.diag[50] ),
    .X(net7520));
 sg13g2_dlygate4sd3_1 hold2972 (.A(_01118_),
    .X(net7521));
 sg13g2_dlygate4sd3_1 hold2973 (.A(\atari2600.tia.diag[36] ),
    .X(net7522));
 sg13g2_dlygate4sd3_1 hold2974 (.A(\atari2600.cpu.load_reg ),
    .X(net7523));
 sg13g2_dlygate4sd3_1 hold2975 (.A(\atari2600.tia.p0_w[3] ),
    .X(net7524));
 sg13g2_dlygate4sd3_1 hold2976 (.A(\atari2600.tia.audc1[0] ),
    .X(net7525));
 sg13g2_dlygate4sd3_1 hold2977 (.A(\atari2600.tia.p1_scale[1] ),
    .X(net7526));
 sg13g2_dlygate4sd3_1 hold2978 (.A(\atari2600.tia.diag[66] ),
    .X(net7527));
 sg13g2_dlygate4sd3_1 hold2979 (.A(\atari2600.tia.audf1[2] ),
    .X(net7528));
 sg13g2_dlygate4sd3_1 hold2980 (.A(\atari2600.tia.audc1[1] ),
    .X(net7529));
 sg13g2_dlygate4sd3_1 hold2981 (.A(\atari2600.tia.diag[37] ),
    .X(net7530));
 sg13g2_dlygate4sd3_1 hold2982 (.A(\atari2600.tia.diag[32] ),
    .X(net7531));
 sg13g2_dlygate4sd3_1 hold2983 (.A(\atari2600.tia.audc0[1] ),
    .X(net7532));
 sg13g2_dlygate4sd3_1 hold2984 (.A(\atari2600.tia.p1_scale[0] ),
    .X(net7533));
 sg13g2_dlygate4sd3_1 hold2985 (.A(\atari2600.cpu.ADD[2] ),
    .X(net7534));
 sg13g2_dlygate4sd3_1 hold2986 (.A(\atari2600.tia.diag[45] ),
    .X(net7535));
 sg13g2_dlygate4sd3_1 hold2987 (.A(\atari2600.tia.diag[65] ),
    .X(net7536));
 sg13g2_dlygate4sd3_1 hold2988 (.A(_01101_),
    .X(net7537));
 sg13g2_dlygate4sd3_1 hold2989 (.A(\atari2600.tia.diag[35] ),
    .X(net7538));
 sg13g2_dlygate4sd3_1 hold2990 (.A(\atari2600.tia.pf_priority ),
    .X(net7539));
 sg13g2_dlygate4sd3_1 hold2991 (.A(\atari2600.clk_counter[1] ),
    .X(net7540));
 sg13g2_dlygate4sd3_1 hold2992 (.A(\atari2600.cpu.ADD[5] ),
    .X(net7541));
 sg13g2_dlygate4sd3_1 hold2993 (.A(_00153_),
    .X(net7542));
 sg13g2_dlygate4sd3_1 hold2994 (.A(\atari2600.tia.audf1[3] ),
    .X(net7543));
 sg13g2_dlygate4sd3_1 hold2995 (.A(\atari2600.tia.diag[70] ),
    .X(net7544));
 sg13g2_dlygate4sd3_1 hold2996 (.A(\atari2600.tia.diag[42] ),
    .X(net7545));
 sg13g2_dlygate4sd3_1 hold2997 (.A(\atari2600.tia.audf1[0] ),
    .X(net7546));
 sg13g2_dlygate4sd3_1 hold2998 (.A(_00152_),
    .X(net7547));
 sg13g2_dlygate4sd3_1 hold2999 (.A(\atari2600.tia.p1_w[3] ),
    .X(net7548));
 sg13g2_dlygate4sd3_1 hold3000 (.A(\atari2600.pia.time_counter[13] ),
    .X(net7549));
 sg13g2_dlygate4sd3_1 hold3001 (.A(\atari2600.tia.diag[56] ),
    .X(net7550));
 sg13g2_dlygate4sd3_1 hold3002 (.A(\atari2600.tia.diag[40] ),
    .X(net7551));
 sg13g2_dlygate4sd3_1 hold3003 (.A(\atari2600.cpu.ADD[4] ),
    .X(net7552));
 sg13g2_dlygate4sd3_1 hold3004 (.A(\atari2600.tia.vdelp0 ),
    .X(net7553));
 sg13g2_dlygate4sd3_1 hold3005 (.A(\atari2600.cpu.ADD[6] ),
    .X(net7554));
 sg13g2_dlygate4sd3_1 hold3006 (.A(\atari2600.tia.diag[57] ),
    .X(net7555));
 sg13g2_dlygate4sd3_1 hold3007 (.A(\b_pwm_even[1] ),
    .X(net7556));
 sg13g2_dlygate4sd3_1 hold3008 (.A(_04696_),
    .X(net7557));
 sg13g2_dlygate4sd3_1 hold3009 (.A(_04704_),
    .X(net7558));
 sg13g2_dlygate4sd3_1 hold3010 (.A(\atari2600.tia.audio_r ),
    .X(net7559));
 sg13g2_dlygate4sd3_1 hold3011 (.A(\atari2600.tia.diag[49] ),
    .X(net7560));
 sg13g2_dlygate4sd3_1 hold3012 (.A(\hvsync_gen.hpos[0] ),
    .X(net7561));
 sg13g2_dlygate4sd3_1 hold3013 (.A(\flash_rom.fsm_state[0] ),
    .X(net7562));
 sg13g2_dlygate4sd3_1 hold3014 (.A(\r_pwm_odd[3] ),
    .X(net7563));
 sg13g2_dlygate4sd3_1 hold3015 (.A(\hvsync_gen.hpos[4] ),
    .X(net7564));
 sg13g2_dlygate4sd3_1 hold3016 (.A(\atari2600.tia.diag[59] ),
    .X(net7565));
 sg13g2_dlygate4sd3_1 hold3017 (.A(\audio_pwm_accumulator[4] ),
    .X(net7566));
 sg13g2_dlygate4sd3_1 hold3018 (.A(\atari2600.tia.diag[33] ),
    .X(net7567));
 sg13g2_dlygate4sd3_1 hold3019 (.A(_01133_),
    .X(net7568));
 sg13g2_dlygate4sd3_1 hold3020 (.A(_00135_),
    .X(net7569));
 sg13g2_dlygate4sd3_1 hold3021 (.A(\atari2600.tia.diag[62] ),
    .X(net7570));
 sg13g2_dlygate4sd3_1 hold3022 (.A(\atari2600.tia.vdelp1 ),
    .X(net7571));
 sg13g2_dlygate4sd3_1 hold3023 (.A(\atari2600.tia.diag[41] ),
    .X(net7572));
 sg13g2_dlygate4sd3_1 hold3024 (.A(_01125_),
    .X(net7573));
 sg13g2_dlygate4sd3_1 hold3025 (.A(_00080_),
    .X(net7574));
 sg13g2_dlygate4sd3_1 hold3026 (.A(_08735_),
    .X(net7575));
 sg13g2_dlygate4sd3_1 hold3027 (.A(\b_pwm_odd[2] ),
    .X(net7576));
 sg13g2_dlygate4sd3_1 hold3028 (.A(\atari2600.tia.audc0[3] ),
    .X(net7577));
 sg13g2_dlygate4sd3_1 hold3029 (.A(\atari2600.tia.hmm0[3] ),
    .X(net7578));
 sg13g2_dlygate4sd3_1 hold3030 (.A(\atari2600.address_bus_r[0] ),
    .X(net7579));
 sg13g2_dlygate4sd3_1 hold3031 (.A(\atari2600.cpu.ADD[0] ),
    .X(net7580));
 sg13g2_dlygate4sd3_1 hold3032 (.A(\atari2600.cpu.plp ),
    .X(net7581));
 sg13g2_dlygate4sd3_1 hold3033 (.A(\atari2600.tia.diag[53] ),
    .X(net7582));
 sg13g2_dlygate4sd3_1 hold3034 (.A(\atari2600.tia.diag[63] ),
    .X(net7583));
 sg13g2_dlygate4sd3_1 hold3035 (.A(\atari2600.stall_cpu ),
    .X(net7584));
 sg13g2_dlygate4sd3_1 hold3036 (.A(\atari2600.address_bus_r[8] ),
    .X(net7585));
 sg13g2_dlygate4sd3_1 hold3037 (.A(\atari2600.tia.diag[58] ),
    .X(net7586));
 sg13g2_dlygate4sd3_1 hold3038 (.A(\atari2600.tia.diag[68] ),
    .X(net7587));
 sg13g2_dlygate4sd3_1 hold3039 (.A(\atari2600.tia.enam0 ),
    .X(net7588));
 sg13g2_dlygate4sd3_1 hold3040 (.A(\atari2600.tia.refpf ),
    .X(net7589));
 sg13g2_dlygate4sd3_1 hold3041 (.A(_00143_),
    .X(net7590));
 sg13g2_dlygate4sd3_1 hold3042 (.A(_00139_),
    .X(net7591));
 sg13g2_dlygate4sd3_1 hold3043 (.A(\atari2600.tia.audc0[2] ),
    .X(net7592));
 sg13g2_dlygate4sd3_1 hold3044 (.A(\atari2600.tia.scorepf ),
    .X(net7593));
 sg13g2_dlygate4sd3_1 hold3045 (.A(\atari2600.tia.audf0[0] ),
    .X(net7594));
 sg13g2_dlygate4sd3_1 hold3046 (.A(\hvsync_gen.vga.vpos[9] ),
    .X(net7595));
 sg13g2_dlygate4sd3_1 hold3047 (.A(_00021_),
    .X(net7596));
 sg13g2_dlygate4sd3_1 hold3048 (.A(\atari2600.pia.time_counter[2] ),
    .X(net7597));
 sg13g2_dlygate4sd3_1 hold3049 (.A(\atari2600.pia.time_counter[13] ),
    .X(net7598));
 sg13g2_dlygate4sd3_1 hold3050 (.A(\atari2600.pia.time_counter[0] ),
    .X(net7599));
 sg13g2_dlygate4sd3_1 hold3051 (.A(\atari2600.tia.colupf[1] ),
    .X(net7600));
 sg13g2_dlygate4sd3_1 hold3052 (.A(\atari2600.tia.cx_clr ),
    .X(net7601));
 sg13g2_antennanp ANTENNA_1 (.A(_00055_));
 sg13g2_antennanp ANTENNA_2 (.A(_00301_));
 sg13g2_antennanp ANTENNA_3 (.A(_01343_));
 sg13g2_antennanp ANTENNA_4 (.A(_01345_));
 sg13g2_antennanp ANTENNA_5 (.A(_01347_));
 sg13g2_antennanp ANTENNA_6 (.A(_05439_));
 sg13g2_antennanp ANTENNA_7 (.A(_08464_));
 sg13g2_antennanp ANTENNA_8 (.A(_08471_));
 sg13g2_antennanp ANTENNA_9 (.A(clk));
 sg13g2_antennanp ANTENNA_10 (.A(clk));
 sg13g2_antennanp ANTENNA_11 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_12 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_13 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_14 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_15 (.A(rst_n));
 sg13g2_antennanp ANTENNA_16 (.A(rst_n));
 sg13g2_antennanp ANTENNA_17 (.A(rst_n));
 sg13g2_antennanp ANTENNA_18 (.A(rst_n));
 sg13g2_antennanp ANTENNA_19 (.A(rst_n));
 sg13g2_antennanp ANTENNA_20 (.A(rst_n));
 sg13g2_antennanp ANTENNA_21 (.A(net6393));
 sg13g2_antennanp ANTENNA_22 (.A(net6393));
 sg13g2_antennanp ANTENNA_23 (.A(net6393));
 sg13g2_antennanp ANTENNA_24 (.A(net6393));
 sg13g2_antennanp ANTENNA_25 (.A(net6393));
 sg13g2_antennanp ANTENNA_26 (.A(net6393));
 sg13g2_antennanp ANTENNA_27 (.A(net6393));
 sg13g2_antennanp ANTENNA_28 (.A(net6393));
 sg13g2_antennanp ANTENNA_29 (.A(net6393));
 sg13g2_antennanp ANTENNA_30 (.A(net6393));
 sg13g2_antennanp ANTENNA_31 (.A(net6393));
 sg13g2_antennanp ANTENNA_32 (.A(net6393));
 sg13g2_antennanp ANTENNA_33 (.A(_00055_));
 sg13g2_antennanp ANTENNA_34 (.A(_00301_));
 sg13g2_antennanp ANTENNA_35 (.A(_00310_));
 sg13g2_antennanp ANTENNA_36 (.A(_00318_));
 sg13g2_antennanp ANTENNA_37 (.A(_00319_));
 sg13g2_antennanp ANTENNA_38 (.A(_00346_));
 sg13g2_antennanp ANTENNA_39 (.A(_00361_));
 sg13g2_antennanp ANTENNA_40 (.A(_01342_));
 sg13g2_antennanp ANTENNA_41 (.A(_01343_));
 sg13g2_antennanp ANTENNA_42 (.A(_01344_));
 sg13g2_antennanp ANTENNA_43 (.A(_01345_));
 sg13g2_antennanp ANTENNA_44 (.A(_01347_));
 sg13g2_antennanp ANTENNA_45 (.A(_05439_));
 sg13g2_antennanp ANTENNA_46 (.A(_08464_));
 sg13g2_antennanp ANTENNA_47 (.A(clk));
 sg13g2_antennanp ANTENNA_48 (.A(clk));
 sg13g2_antennanp ANTENNA_49 (.A(net5605));
 sg13g2_antennanp ANTENNA_50 (.A(net5605));
 sg13g2_antennanp ANTENNA_51 (.A(net5605));
 sg13g2_antennanp ANTENNA_52 (.A(net5605));
 sg13g2_antennanp ANTENNA_53 (.A(net5605));
 sg13g2_antennanp ANTENNA_54 (.A(net5605));
 sg13g2_antennanp ANTENNA_55 (.A(net5605));
 sg13g2_antennanp ANTENNA_56 (.A(net5605));
 sg13g2_antennanp ANTENNA_57 (.A(net5605));
 sg13g2_antennanp ANTENNA_58 (.A(net5605));
 sg13g2_antennanp ANTENNA_59 (.A(net5605));
 sg13g2_antennanp ANTENNA_60 (.A(net6393));
 sg13g2_antennanp ANTENNA_61 (.A(net6393));
 sg13g2_antennanp ANTENNA_62 (.A(net6393));
 sg13g2_antennanp ANTENNA_63 (.A(net6393));
 sg13g2_antennanp ANTENNA_64 (.A(net6393));
 sg13g2_antennanp ANTENNA_65 (.A(net6393));
 sg13g2_antennanp ANTENNA_66 (.A(net6393));
 sg13g2_antennanp ANTENNA_67 (.A(net6393));
 sg13g2_antennanp ANTENNA_68 (.A(net6393));
 sg13g2_antennanp ANTENNA_69 (.A(net6393));
 sg13g2_antennanp ANTENNA_70 (.A(net6393));
 sg13g2_antennanp ANTENNA_71 (.A(net6393));
 sg13g2_antennanp ANTENNA_72 (.A(_00301_));
 sg13g2_antennanp ANTENNA_73 (.A(_00310_));
 sg13g2_antennanp ANTENNA_74 (.A(_00319_));
 sg13g2_antennanp ANTENNA_75 (.A(_00346_));
 sg13g2_antennanp ANTENNA_76 (.A(_00361_));
 sg13g2_antennanp ANTENNA_77 (.A(_01343_));
 sg13g2_antennanp ANTENNA_78 (.A(_01344_));
 sg13g2_antennanp ANTENNA_79 (.A(_01345_));
 sg13g2_antennanp ANTENNA_80 (.A(_01347_));
 sg13g2_antennanp ANTENNA_81 (.A(_05439_));
 sg13g2_antennanp ANTENNA_82 (.A(_08464_));
 sg13g2_antennanp ANTENNA_83 (.A(clk));
 sg13g2_antennanp ANTENNA_84 (.A(clk));
 sg13g2_antennanp ANTENNA_85 (.A(net5254));
 sg13g2_antennanp ANTENNA_86 (.A(net5254));
 sg13g2_antennanp ANTENNA_87 (.A(net5254));
 sg13g2_antennanp ANTENNA_88 (.A(net5254));
 sg13g2_antennanp ANTENNA_89 (.A(net5254));
 sg13g2_antennanp ANTENNA_90 (.A(net5254));
 sg13g2_antennanp ANTENNA_91 (.A(net5254));
 sg13g2_antennanp ANTENNA_92 (.A(net5254));
 sg13g2_antennanp ANTENNA_93 (.A(net5605));
 sg13g2_antennanp ANTENNA_94 (.A(net5605));
 sg13g2_antennanp ANTENNA_95 (.A(net5605));
 sg13g2_antennanp ANTENNA_96 (.A(net5605));
 sg13g2_antennanp ANTENNA_97 (.A(net5605));
 sg13g2_antennanp ANTENNA_98 (.A(net5605));
 sg13g2_antennanp ANTENNA_99 (.A(net5605));
 sg13g2_antennanp ANTENNA_100 (.A(net5605));
 sg13g2_antennanp ANTENNA_101 (.A(net5605));
 sg13g2_antennanp ANTENNA_102 (.A(net5605));
 sg13g2_antennanp ANTENNA_103 (.A(net5605));
 sg13g2_antennanp ANTENNA_104 (.A(net5605));
 sg13g2_antennanp ANTENNA_105 (.A(net5605));
 sg13g2_antennanp ANTENNA_106 (.A(net6393));
 sg13g2_antennanp ANTENNA_107 (.A(net6393));
 sg13g2_antennanp ANTENNA_108 (.A(net6393));
 sg13g2_antennanp ANTENNA_109 (.A(net6393));
 sg13g2_antennanp ANTENNA_110 (.A(net6393));
 sg13g2_antennanp ANTENNA_111 (.A(net6393));
 sg13g2_antennanp ANTENNA_112 (.A(net6393));
 sg13g2_antennanp ANTENNA_113 (.A(net6393));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_4 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_88 ();
 sg13g2_fill_2 FILLER_0_184 ();
 sg13g2_fill_1 FILLER_0_186 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_2 FILLER_0_237 ();
 sg13g2_fill_2 FILLER_0_305 ();
 sg13g2_fill_1 FILLER_0_307 ();
 sg13g2_fill_2 FILLER_0_317 ();
 sg13g2_fill_2 FILLER_0_345 ();
 sg13g2_fill_1 FILLER_0_347 ();
 sg13g2_fill_1 FILLER_0_382 ();
 sg13g2_fill_2 FILLER_0_400 ();
 sg13g2_fill_1 FILLER_0_402 ();
 sg13g2_fill_2 FILLER_0_412 ();
 sg13g2_fill_1 FILLER_0_414 ();
 sg13g2_fill_1 FILLER_0_485 ();
 sg13g2_fill_1 FILLER_0_513 ();
 sg13g2_fill_2 FILLER_0_578 ();
 sg13g2_fill_1 FILLER_0_589 ();
 sg13g2_fill_2 FILLER_0_650 ();
 sg13g2_fill_2 FILLER_0_699 ();
 sg13g2_fill_1 FILLER_0_701 ();
 sg13g2_fill_2 FILLER_0_728 ();
 sg13g2_fill_1 FILLER_0_730 ();
 sg13g2_fill_1 FILLER_0_761 ();
 sg13g2_fill_2 FILLER_0_771 ();
 sg13g2_fill_1 FILLER_0_799 ();
 sg13g2_fill_2 FILLER_0_845 ();
 sg13g2_fill_2 FILLER_0_865 ();
 sg13g2_fill_2 FILLER_0_923 ();
 sg13g2_fill_1 FILLER_0_925 ();
 sg13g2_fill_1 FILLER_0_931 ();
 sg13g2_fill_2 FILLER_0_986 ();
 sg13g2_fill_1 FILLER_0_1001 ();
 sg13g2_fill_1 FILLER_0_1036 ();
 sg13g2_fill_2 FILLER_0_1071 ();
 sg13g2_fill_1 FILLER_0_1073 ();
 sg13g2_fill_2 FILLER_0_1109 ();
 sg13g2_fill_2 FILLER_0_1123 ();
 sg13g2_fill_1 FILLER_0_1125 ();
 sg13g2_fill_2 FILLER_0_1139 ();
 sg13g2_fill_1 FILLER_0_1141 ();
 sg13g2_fill_1 FILLER_0_1151 ();
 sg13g2_fill_1 FILLER_0_1204 ();
 sg13g2_fill_1 FILLER_0_1210 ();
 sg13g2_fill_1 FILLER_0_1225 ();
 sg13g2_fill_2 FILLER_0_1270 ();
 sg13g2_fill_1 FILLER_0_1272 ();
 sg13g2_fill_2 FILLER_0_1283 ();
 sg13g2_fill_2 FILLER_0_1315 ();
 sg13g2_fill_1 FILLER_0_1354 ();
 sg13g2_fill_2 FILLER_0_1368 ();
 sg13g2_decap_4 FILLER_0_1429 ();
 sg13g2_fill_1 FILLER_0_1433 ();
 sg13g2_fill_2 FILLER_0_1460 ();
 sg13g2_fill_2 FILLER_0_1475 ();
 sg13g2_fill_1 FILLER_0_1477 ();
 sg13g2_fill_2 FILLER_0_1506 ();
 sg13g2_fill_1 FILLER_0_1508 ();
 sg13g2_fill_2 FILLER_0_1535 ();
 sg13g2_fill_2 FILLER_0_1551 ();
 sg13g2_fill_1 FILLER_0_1579 ();
 sg13g2_fill_2 FILLER_0_1610 ();
 sg13g2_fill_1 FILLER_0_1612 ();
 sg13g2_fill_2 FILLER_0_1658 ();
 sg13g2_fill_2 FILLER_0_1700 ();
 sg13g2_fill_1 FILLER_0_1702 ();
 sg13g2_fill_2 FILLER_0_1756 ();
 sg13g2_fill_1 FILLER_0_1758 ();
 sg13g2_fill_1 FILLER_0_1763 ();
 sg13g2_fill_2 FILLER_0_1773 ();
 sg13g2_fill_1 FILLER_0_1775 ();
 sg13g2_fill_1 FILLER_0_1802 ();
 sg13g2_fill_2 FILLER_0_1822 ();
 sg13g2_fill_1 FILLER_0_1855 ();
 sg13g2_fill_2 FILLER_0_1894 ();
 sg13g2_fill_2 FILLER_0_1929 ();
 sg13g2_fill_1 FILLER_0_1931 ();
 sg13g2_fill_2 FILLER_0_1970 ();
 sg13g2_fill_1 FILLER_0_1972 ();
 sg13g2_fill_2 FILLER_0_1986 ();
 sg13g2_decap_4 FILLER_0_2041 ();
 sg13g2_fill_2 FILLER_0_2045 ();
 sg13g2_decap_8 FILLER_0_2056 ();
 sg13g2_decap_8 FILLER_0_2063 ();
 sg13g2_decap_8 FILLER_0_2070 ();
 sg13g2_decap_8 FILLER_0_2077 ();
 sg13g2_fill_2 FILLER_0_2130 ();
 sg13g2_fill_2 FILLER_0_2158 ();
 sg13g2_fill_2 FILLER_0_2195 ();
 sg13g2_fill_2 FILLER_0_2231 ();
 sg13g2_fill_1 FILLER_0_2233 ();
 sg13g2_fill_2 FILLER_0_2248 ();
 sg13g2_fill_1 FILLER_0_2250 ();
 sg13g2_fill_1 FILLER_0_2270 ();
 sg13g2_fill_2 FILLER_0_2289 ();
 sg13g2_fill_1 FILLER_0_2291 ();
 sg13g2_decap_4 FILLER_0_2301 ();
 sg13g2_fill_2 FILLER_0_2305 ();
 sg13g2_decap_4 FILLER_0_2371 ();
 sg13g2_fill_2 FILLER_0_2385 ();
 sg13g2_fill_1 FILLER_0_2387 ();
 sg13g2_fill_1 FILLER_0_2427 ();
 sg13g2_fill_1 FILLER_0_2447 ();
 sg13g2_fill_2 FILLER_0_2488 ();
 sg13g2_fill_1 FILLER_0_2509 ();
 sg13g2_decap_8 FILLER_0_2549 ();
 sg13g2_decap_8 FILLER_0_2556 ();
 sg13g2_decap_8 FILLER_0_2563 ();
 sg13g2_decap_8 FILLER_0_2570 ();
 sg13g2_decap_8 FILLER_0_2577 ();
 sg13g2_decap_8 FILLER_0_2584 ();
 sg13g2_decap_8 FILLER_0_2591 ();
 sg13g2_decap_8 FILLER_0_2598 ();
 sg13g2_decap_8 FILLER_0_2605 ();
 sg13g2_decap_8 FILLER_0_2612 ();
 sg13g2_decap_8 FILLER_0_2619 ();
 sg13g2_decap_8 FILLER_0_2626 ();
 sg13g2_decap_8 FILLER_0_2633 ();
 sg13g2_decap_8 FILLER_0_2640 ();
 sg13g2_decap_8 FILLER_0_2647 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_decap_4 FILLER_0_2668 ();
 sg13g2_fill_2 FILLER_0_2672 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_91 ();
 sg13g2_fill_1 FILLER_1_95 ();
 sg13g2_fill_2 FILLER_1_136 ();
 sg13g2_fill_1 FILLER_1_138 ();
 sg13g2_fill_2 FILLER_1_165 ();
 sg13g2_fill_1 FILLER_1_167 ();
 sg13g2_fill_2 FILLER_1_192 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_fill_1 FILLER_1_262 ();
 sg13g2_fill_2 FILLER_1_272 ();
 sg13g2_fill_1 FILLER_1_274 ();
 sg13g2_fill_2 FILLER_1_289 ();
 sg13g2_fill_2 FILLER_1_317 ();
 sg13g2_fill_2 FILLER_1_333 ();
 sg13g2_fill_2 FILLER_1_457 ();
 sg13g2_fill_1 FILLER_1_459 ();
 sg13g2_fill_2 FILLER_1_465 ();
 sg13g2_fill_1 FILLER_1_537 ();
 sg13g2_fill_2 FILLER_1_558 ();
 sg13g2_fill_1 FILLER_1_632 ();
 sg13g2_fill_1 FILLER_1_664 ();
 sg13g2_fill_1 FILLER_1_715 ();
 sg13g2_fill_2 FILLER_1_721 ();
 sg13g2_fill_1 FILLER_1_744 ();
 sg13g2_fill_2 FILLER_1_771 ();
 sg13g2_fill_2 FILLER_1_801 ();
 sg13g2_fill_1 FILLER_1_803 ();
 sg13g2_fill_1 FILLER_1_900 ();
 sg13g2_fill_2 FILLER_1_957 ();
 sg13g2_fill_2 FILLER_1_1016 ();
 sg13g2_fill_1 FILLER_1_1018 ();
 sg13g2_fill_2 FILLER_1_1038 ();
 sg13g2_fill_1 FILLER_1_1065 ();
 sg13g2_fill_2 FILLER_1_1071 ();
 sg13g2_fill_2 FILLER_1_1160 ();
 sg13g2_fill_2 FILLER_1_1176 ();
 sg13g2_fill_1 FILLER_1_1457 ();
 sg13g2_fill_1 FILLER_1_1533 ();
 sg13g2_fill_2 FILLER_1_1617 ();
 sg13g2_decap_4 FILLER_1_1645 ();
 sg13g2_fill_1 FILLER_1_1649 ();
 sg13g2_fill_1 FILLER_1_1704 ();
 sg13g2_fill_2 FILLER_1_1725 ();
 sg13g2_fill_2 FILLER_1_1833 ();
 sg13g2_fill_1 FILLER_1_1835 ();
 sg13g2_fill_1 FILLER_1_1845 ();
 sg13g2_fill_2 FILLER_1_2000 ();
 sg13g2_decap_8 FILLER_1_2064 ();
 sg13g2_fill_1 FILLER_1_2071 ();
 sg13g2_fill_1 FILLER_1_2143 ();
 sg13g2_fill_1 FILLER_1_2189 ();
 sg13g2_fill_2 FILLER_1_2204 ();
 sg13g2_fill_1 FILLER_1_2414 ();
 sg13g2_fill_2 FILLER_1_2463 ();
 sg13g2_fill_2 FILLER_1_2475 ();
 sg13g2_fill_1 FILLER_1_2477 ();
 sg13g2_decap_8 FILLER_1_2549 ();
 sg13g2_decap_8 FILLER_1_2556 ();
 sg13g2_decap_8 FILLER_1_2563 ();
 sg13g2_decap_8 FILLER_1_2570 ();
 sg13g2_decap_8 FILLER_1_2577 ();
 sg13g2_decap_8 FILLER_1_2584 ();
 sg13g2_decap_8 FILLER_1_2591 ();
 sg13g2_decap_8 FILLER_1_2598 ();
 sg13g2_decap_8 FILLER_1_2605 ();
 sg13g2_decap_8 FILLER_1_2612 ();
 sg13g2_decap_8 FILLER_1_2619 ();
 sg13g2_decap_8 FILLER_1_2626 ();
 sg13g2_decap_8 FILLER_1_2633 ();
 sg13g2_decap_8 FILLER_1_2640 ();
 sg13g2_decap_8 FILLER_1_2647 ();
 sg13g2_decap_8 FILLER_1_2654 ();
 sg13g2_decap_8 FILLER_1_2661 ();
 sg13g2_decap_4 FILLER_1_2668 ();
 sg13g2_fill_2 FILLER_1_2672 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_84 ();
 sg13g2_fill_2 FILLER_2_88 ();
 sg13g2_fill_2 FILLER_2_130 ();
 sg13g2_fill_1 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_195 ();
 sg13g2_fill_1 FILLER_2_222 ();
 sg13g2_fill_2 FILLER_2_232 ();
 sg13g2_fill_1 FILLER_2_234 ();
 sg13g2_fill_2 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_fill_1 FILLER_2_330 ();
 sg13g2_fill_2 FILLER_2_366 ();
 sg13g2_fill_2 FILLER_2_390 ();
 sg13g2_fill_2 FILLER_2_397 ();
 sg13g2_fill_2 FILLER_2_423 ();
 sg13g2_fill_1 FILLER_2_439 ();
 sg13g2_fill_2 FILLER_2_454 ();
 sg13g2_fill_2 FILLER_2_493 ();
 sg13g2_fill_1 FILLER_2_495 ();
 sg13g2_fill_2 FILLER_2_594 ();
 sg13g2_fill_2 FILLER_2_634 ();
 sg13g2_fill_1 FILLER_2_636 ();
 sg13g2_fill_2 FILLER_2_651 ();
 sg13g2_fill_1 FILLER_2_653 ();
 sg13g2_fill_1 FILLER_2_663 ();
 sg13g2_fill_2 FILLER_2_672 ();
 sg13g2_fill_1 FILLER_2_674 ();
 sg13g2_fill_2 FILLER_2_684 ();
 sg13g2_fill_2 FILLER_2_733 ();
 sg13g2_fill_2 FILLER_2_740 ();
 sg13g2_fill_2 FILLER_2_841 ();
 sg13g2_fill_2 FILLER_2_968 ();
 sg13g2_fill_2 FILLER_2_996 ();
 sg13g2_fill_2 FILLER_2_1053 ();
 sg13g2_fill_2 FILLER_2_1087 ();
 sg13g2_fill_1 FILLER_2_1089 ();
 sg13g2_fill_1 FILLER_2_1103 ();
 sg13g2_fill_2 FILLER_2_1119 ();
 sg13g2_fill_1 FILLER_2_1121 ();
 sg13g2_fill_2 FILLER_2_1132 ();
 sg13g2_fill_2 FILLER_2_1139 ();
 sg13g2_fill_2 FILLER_2_1265 ();
 sg13g2_fill_2 FILLER_2_1281 ();
 sg13g2_fill_2 FILLER_2_1306 ();
 sg13g2_fill_1 FILLER_2_1308 ();
 sg13g2_fill_2 FILLER_2_1347 ();
 sg13g2_fill_2 FILLER_2_1354 ();
 sg13g2_decap_8 FILLER_2_1364 ();
 sg13g2_fill_1 FILLER_2_1371 ();
 sg13g2_fill_1 FILLER_2_1390 ();
 sg13g2_decap_8 FILLER_2_1396 ();
 sg13g2_decap_4 FILLER_2_1403 ();
 sg13g2_fill_2 FILLER_2_1442 ();
 sg13g2_fill_1 FILLER_2_1444 ();
 sg13g2_fill_2 FILLER_2_1475 ();
 sg13g2_fill_1 FILLER_2_1482 ();
 sg13g2_fill_1 FILLER_2_1492 ();
 sg13g2_decap_4 FILLER_2_1620 ();
 sg13g2_fill_2 FILLER_2_1624 ();
 sg13g2_fill_2 FILLER_2_1634 ();
 sg13g2_fill_1 FILLER_2_1645 ();
 sg13g2_fill_2 FILLER_2_1665 ();
 sg13g2_fill_2 FILLER_2_1688 ();
 sg13g2_fill_1 FILLER_2_1690 ();
 sg13g2_fill_2 FILLER_2_1717 ();
 sg13g2_fill_1 FILLER_2_1719 ();
 sg13g2_fill_2 FILLER_2_1741 ();
 sg13g2_fill_2 FILLER_2_1818 ();
 sg13g2_fill_1 FILLER_2_1820 ();
 sg13g2_fill_1 FILLER_2_1848 ();
 sg13g2_fill_1 FILLER_2_1921 ();
 sg13g2_fill_1 FILLER_2_1931 ();
 sg13g2_fill_2 FILLER_2_1977 ();
 sg13g2_decap_8 FILLER_2_2029 ();
 sg13g2_fill_1 FILLER_2_2057 ();
 sg13g2_fill_1 FILLER_2_2094 ();
 sg13g2_fill_2 FILLER_2_2120 ();
 sg13g2_fill_2 FILLER_2_2148 ();
 sg13g2_fill_2 FILLER_2_2176 ();
 sg13g2_fill_1 FILLER_2_2178 ();
 sg13g2_fill_2 FILLER_2_2244 ();
 sg13g2_fill_2 FILLER_2_2288 ();
 sg13g2_fill_1 FILLER_2_2302 ();
 sg13g2_fill_1 FILLER_2_2313 ();
 sg13g2_fill_2 FILLER_2_2318 ();
 sg13g2_fill_1 FILLER_2_2320 ();
 sg13g2_fill_2 FILLER_2_2331 ();
 sg13g2_fill_1 FILLER_2_2333 ();
 sg13g2_decap_4 FILLER_2_2364 ();
 sg13g2_fill_1 FILLER_2_2368 ();
 sg13g2_fill_2 FILLER_2_2379 ();
 sg13g2_fill_2 FILLER_2_2474 ();
 sg13g2_fill_1 FILLER_2_2476 ();
 sg13g2_fill_1 FILLER_2_2518 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_4 FILLER_2_2553 ();
 sg13g2_fill_1 FILLER_2_2557 ();
 sg13g2_fill_2 FILLER_2_2562 ();
 sg13g2_fill_1 FILLER_2_2564 ();
 sg13g2_fill_1 FILLER_2_2570 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_decap_8 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2601 ();
 sg13g2_fill_2 FILLER_2_2608 ();
 sg13g2_fill_1 FILLER_2_2610 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_decap_8 FILLER_2_2622 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_decap_8 FILLER_2_2636 ();
 sg13g2_decap_8 FILLER_2_2643 ();
 sg13g2_decap_8 FILLER_2_2650 ();
 sg13g2_decap_8 FILLER_2_2657 ();
 sg13g2_decap_8 FILLER_2_2664 ();
 sg13g2_fill_2 FILLER_2_2671 ();
 sg13g2_fill_1 FILLER_2_2673 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_93 ();
 sg13g2_fill_2 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_fill_2 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_293 ();
 sg13g2_fill_1 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_380 ();
 sg13g2_fill_1 FILLER_3_416 ();
 sg13g2_fill_1 FILLER_3_434 ();
 sg13g2_fill_1 FILLER_3_461 ();
 sg13g2_fill_1 FILLER_3_492 ();
 sg13g2_fill_2 FILLER_3_541 ();
 sg13g2_fill_1 FILLER_3_543 ();
 sg13g2_fill_2 FILLER_3_568 ();
 sg13g2_fill_1 FILLER_3_649 ();
 sg13g2_fill_1 FILLER_3_676 ();
 sg13g2_fill_1 FILLER_3_729 ();
 sg13g2_fill_1 FILLER_3_756 ();
 sg13g2_fill_1 FILLER_3_772 ();
 sg13g2_fill_1 FILLER_3_881 ();
 sg13g2_fill_2 FILLER_3_942 ();
 sg13g2_fill_1 FILLER_3_944 ();
 sg13g2_fill_1 FILLER_3_954 ();
 sg13g2_fill_2 FILLER_3_980 ();
 sg13g2_fill_2 FILLER_3_1039 ();
 sg13g2_fill_2 FILLER_3_1055 ();
 sg13g2_fill_1 FILLER_3_1057 ();
 sg13g2_fill_2 FILLER_3_1116 ();
 sg13g2_fill_1 FILLER_3_1118 ();
 sg13g2_fill_2 FILLER_3_1193 ();
 sg13g2_fill_1 FILLER_3_1221 ();
 sg13g2_fill_1 FILLER_3_1231 ();
 sg13g2_fill_1 FILLER_3_1241 ();
 sg13g2_fill_1 FILLER_3_1281 ();
 sg13g2_fill_2 FILLER_3_1313 ();
 sg13g2_fill_2 FILLER_3_1411 ();
 sg13g2_fill_1 FILLER_3_1422 ();
 sg13g2_fill_1 FILLER_3_1561 ();
 sg13g2_fill_2 FILLER_3_1574 ();
 sg13g2_fill_1 FILLER_3_1581 ();
 sg13g2_fill_2 FILLER_3_1617 ();
 sg13g2_decap_4 FILLER_3_1645 ();
 sg13g2_fill_2 FILLER_3_1663 ();
 sg13g2_fill_2 FILLER_3_1705 ();
 sg13g2_fill_1 FILLER_3_1707 ();
 sg13g2_fill_1 FILLER_3_1762 ();
 sg13g2_fill_2 FILLER_3_1772 ();
 sg13g2_fill_1 FILLER_3_1774 ();
 sg13g2_fill_1 FILLER_3_1905 ();
 sg13g2_fill_1 FILLER_3_1942 ();
 sg13g2_fill_2 FILLER_3_1989 ();
 sg13g2_fill_2 FILLER_3_2019 ();
 sg13g2_fill_2 FILLER_3_2047 ();
 sg13g2_fill_1 FILLER_3_2049 ();
 sg13g2_fill_2 FILLER_3_2111 ();
 sg13g2_fill_1 FILLER_3_2113 ();
 sg13g2_fill_2 FILLER_3_2124 ();
 sg13g2_fill_2 FILLER_3_2143 ();
 sg13g2_fill_1 FILLER_3_2145 ();
 sg13g2_fill_2 FILLER_3_2165 ();
 sg13g2_fill_1 FILLER_3_2167 ();
 sg13g2_fill_2 FILLER_3_2215 ();
 sg13g2_fill_1 FILLER_3_2217 ();
 sg13g2_fill_2 FILLER_3_2248 ();
 sg13g2_fill_1 FILLER_3_2250 ();
 sg13g2_fill_1 FILLER_3_2277 ();
 sg13g2_fill_2 FILLER_3_2301 ();
 sg13g2_fill_1 FILLER_3_2407 ();
 sg13g2_fill_2 FILLER_3_2458 ();
 sg13g2_fill_1 FILLER_3_2460 ();
 sg13g2_fill_2 FILLER_3_2581 ();
 sg13g2_fill_1 FILLER_3_2583 ();
 sg13g2_decap_8 FILLER_3_2588 ();
 sg13g2_decap_4 FILLER_3_2595 ();
 sg13g2_fill_1 FILLER_3_2599 ();
 sg13g2_decap_8 FILLER_3_2626 ();
 sg13g2_fill_2 FILLER_3_2633 ();
 sg13g2_fill_1 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2662 ();
 sg13g2_decap_4 FILLER_3_2669 ();
 sg13g2_fill_1 FILLER_3_2673 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_4 FILLER_4_84 ();
 sg13g2_fill_2 FILLER_4_154 ();
 sg13g2_fill_1 FILLER_4_156 ();
 sg13g2_fill_2 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_272 ();
 sg13g2_fill_2 FILLER_4_365 ();
 sg13g2_fill_1 FILLER_4_367 ();
 sg13g2_fill_1 FILLER_4_467 ();
 sg13g2_fill_2 FILLER_4_516 ();
 sg13g2_fill_2 FILLER_4_531 ();
 sg13g2_fill_1 FILLER_4_533 ();
 sg13g2_fill_2 FILLER_4_548 ();
 sg13g2_fill_2 FILLER_4_585 ();
 sg13g2_fill_1 FILLER_4_587 ();
 sg13g2_fill_2 FILLER_4_614 ();
 sg13g2_fill_1 FILLER_4_616 ();
 sg13g2_fill_1 FILLER_4_651 ();
 sg13g2_fill_1 FILLER_4_661 ();
 sg13g2_fill_1 FILLER_4_702 ();
 sg13g2_fill_1 FILLER_4_729 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_fill_2 FILLER_4_798 ();
 sg13g2_fill_2 FILLER_4_809 ();
 sg13g2_fill_1 FILLER_4_811 ();
 sg13g2_fill_2 FILLER_4_825 ();
 sg13g2_fill_1 FILLER_4_827 ();
 sg13g2_fill_2 FILLER_4_859 ();
 sg13g2_fill_2 FILLER_4_866 ();
 sg13g2_fill_1 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_895 ();
 sg13g2_fill_1 FILLER_4_897 ();
 sg13g2_fill_1 FILLER_4_912 ();
 sg13g2_fill_1 FILLER_4_966 ();
 sg13g2_fill_1 FILLER_4_1004 ();
 sg13g2_fill_2 FILLER_4_1015 ();
 sg13g2_fill_2 FILLER_4_1069 ();
 sg13g2_fill_1 FILLER_4_1071 ();
 sg13g2_fill_2 FILLER_4_1098 ();
 sg13g2_fill_1 FILLER_4_1100 ();
 sg13g2_fill_1 FILLER_4_1114 ();
 sg13g2_fill_1 FILLER_4_1198 ();
 sg13g2_fill_1 FILLER_4_1297 ();
 sg13g2_fill_2 FILLER_4_1348 ();
 sg13g2_fill_1 FILLER_4_1355 ();
 sg13g2_fill_2 FILLER_4_1402 ();
 sg13g2_fill_2 FILLER_4_1427 ();
 sg13g2_fill_1 FILLER_4_1465 ();
 sg13g2_fill_2 FILLER_4_1486 ();
 sg13g2_fill_2 FILLER_4_1516 ();
 sg13g2_fill_2 FILLER_4_1539 ();
 sg13g2_fill_2 FILLER_4_1578 ();
 sg13g2_fill_1 FILLER_4_1580 ();
 sg13g2_fill_1 FILLER_4_1617 ();
 sg13g2_fill_1 FILLER_4_1709 ();
 sg13g2_fill_2 FILLER_4_1762 ();
 sg13g2_fill_2 FILLER_4_1933 ();
 sg13g2_fill_1 FILLER_4_1935 ();
 sg13g2_fill_2 FILLER_4_1976 ();
 sg13g2_fill_1 FILLER_4_1978 ();
 sg13g2_fill_1 FILLER_4_2044 ();
 sg13g2_decap_8 FILLER_4_2072 ();
 sg13g2_decap_4 FILLER_4_2079 ();
 sg13g2_fill_2 FILLER_4_2093 ();
 sg13g2_fill_2 FILLER_4_2108 ();
 sg13g2_fill_1 FILLER_4_2178 ();
 sg13g2_fill_2 FILLER_4_2183 ();
 sg13g2_fill_2 FILLER_4_2256 ();
 sg13g2_decap_8 FILLER_4_2309 ();
 sg13g2_fill_2 FILLER_4_2316 ();
 sg13g2_decap_8 FILLER_4_2327 ();
 sg13g2_fill_1 FILLER_4_2334 ();
 sg13g2_fill_1 FILLER_4_2345 ();
 sg13g2_fill_2 FILLER_4_2365 ();
 sg13g2_fill_2 FILLER_4_2376 ();
 sg13g2_fill_1 FILLER_4_2378 ();
 sg13g2_fill_2 FILLER_4_2424 ();
 sg13g2_fill_1 FILLER_4_2426 ();
 sg13g2_fill_1 FILLER_4_2484 ();
 sg13g2_fill_1 FILLER_4_2543 ();
 sg13g2_fill_2 FILLER_4_2653 ();
 sg13g2_decap_4 FILLER_4_2668 ();
 sg13g2_fill_2 FILLER_4_2672 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_4 FILLER_5_70 ();
 sg13g2_fill_2 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_fill_1 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_1 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_379 ();
 sg13g2_fill_1 FILLER_5_381 ();
 sg13g2_fill_2 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_5_550 ();
 sg13g2_fill_1 FILLER_5_627 ();
 sg13g2_fill_2 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_701 ();
 sg13g2_fill_1 FILLER_5_729 ();
 sg13g2_fill_1 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_785 ();
 sg13g2_fill_1 FILLER_5_787 ();
 sg13g2_fill_2 FILLER_5_848 ();
 sg13g2_fill_1 FILLER_5_928 ();
 sg13g2_fill_2 FILLER_5_939 ();
 sg13g2_fill_1 FILLER_5_941 ();
 sg13g2_fill_2 FILLER_5_970 ();
 sg13g2_fill_2 FILLER_5_1004 ();
 sg13g2_fill_1 FILLER_5_1006 ();
 sg13g2_fill_1 FILLER_5_1090 ();
 sg13g2_fill_2 FILLER_5_1108 ();
 sg13g2_fill_1 FILLER_5_1110 ();
 sg13g2_fill_2 FILLER_5_1142 ();
 sg13g2_fill_1 FILLER_5_1144 ();
 sg13g2_fill_1 FILLER_5_1155 ();
 sg13g2_fill_2 FILLER_5_1162 ();
 sg13g2_fill_1 FILLER_5_1164 ();
 sg13g2_fill_1 FILLER_5_1188 ();
 sg13g2_fill_1 FILLER_5_1255 ();
 sg13g2_fill_2 FILLER_5_1284 ();
 sg13g2_fill_1 FILLER_5_1295 ();
 sg13g2_fill_1 FILLER_5_1305 ();
 sg13g2_fill_2 FILLER_5_1311 ();
 sg13g2_fill_2 FILLER_5_1330 ();
 sg13g2_fill_1 FILLER_5_1332 ();
 sg13g2_fill_1 FILLER_5_1392 ();
 sg13g2_fill_2 FILLER_5_1437 ();
 sg13g2_fill_1 FILLER_5_1439 ();
 sg13g2_fill_2 FILLER_5_1465 ();
 sg13g2_fill_1 FILLER_5_1535 ();
 sg13g2_fill_2 FILLER_5_1595 ();
 sg13g2_fill_1 FILLER_5_1597 ();
 sg13g2_fill_2 FILLER_5_1603 ();
 sg13g2_fill_1 FILLER_5_1605 ();
 sg13g2_fill_2 FILLER_5_1622 ();
 sg13g2_fill_1 FILLER_5_1624 ();
 sg13g2_fill_1 FILLER_5_1644 ();
 sg13g2_fill_1 FILLER_5_1681 ();
 sg13g2_decap_4 FILLER_5_1696 ();
 sg13g2_fill_2 FILLER_5_1735 ();
 sg13g2_fill_1 FILLER_5_1737 ();
 sg13g2_fill_2 FILLER_5_1837 ();
 sg13g2_fill_1 FILLER_5_1839 ();
 sg13g2_fill_2 FILLER_5_1859 ();
 sg13g2_fill_1 FILLER_5_1861 ();
 sg13g2_fill_2 FILLER_5_1924 ();
 sg13g2_fill_1 FILLER_5_1926 ();
 sg13g2_fill_1 FILLER_5_1931 ();
 sg13g2_fill_1 FILLER_5_1946 ();
 sg13g2_fill_1 FILLER_5_1962 ();
 sg13g2_fill_2 FILLER_5_2067 ();
 sg13g2_fill_1 FILLER_5_2069 ();
 sg13g2_fill_1 FILLER_5_2129 ();
 sg13g2_fill_1 FILLER_5_2187 ();
 sg13g2_fill_1 FILLER_5_2201 ();
 sg13g2_fill_2 FILLER_5_2248 ();
 sg13g2_decap_4 FILLER_5_2289 ();
 sg13g2_fill_1 FILLER_5_2337 ();
 sg13g2_fill_2 FILLER_5_2372 ();
 sg13g2_fill_1 FILLER_5_2374 ();
 sg13g2_fill_2 FILLER_5_2419 ();
 sg13g2_fill_2 FILLER_5_2427 ();
 sg13g2_fill_1 FILLER_5_2429 ();
 sg13g2_decap_4 FILLER_5_2440 ();
 sg13g2_fill_1 FILLER_5_2458 ();
 sg13g2_decap_8 FILLER_5_2478 ();
 sg13g2_fill_1 FILLER_5_2504 ();
 sg13g2_fill_2 FILLER_5_2518 ();
 sg13g2_fill_1 FILLER_5_2520 ();
 sg13g2_fill_2 FILLER_5_2555 ();
 sg13g2_fill_2 FILLER_5_2631 ();
 sg13g2_fill_1 FILLER_5_2633 ();
 sg13g2_decap_4 FILLER_5_2670 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_fill_2 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_103 ();
 sg13g2_fill_1 FILLER_6_105 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_284 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_318 ();
 sg13g2_fill_2 FILLER_6_329 ();
 sg13g2_fill_1 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_fill_2 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_6_399 ();
 sg13g2_fill_1 FILLER_6_426 ();
 sg13g2_fill_1 FILLER_6_442 ();
 sg13g2_fill_2 FILLER_6_467 ();
 sg13g2_fill_2 FILLER_6_522 ();
 sg13g2_fill_1 FILLER_6_524 ();
 sg13g2_fill_2 FILLER_6_598 ();
 sg13g2_fill_1 FILLER_6_600 ();
 sg13g2_fill_1 FILLER_6_697 ();
 sg13g2_fill_2 FILLER_6_703 ();
 sg13g2_fill_1 FILLER_6_705 ();
 sg13g2_fill_2 FILLER_6_737 ();
 sg13g2_fill_1 FILLER_6_774 ();
 sg13g2_fill_1 FILLER_6_801 ();
 sg13g2_fill_1 FILLER_6_858 ();
 sg13g2_fill_1 FILLER_6_873 ();
 sg13g2_fill_2 FILLER_6_930 ();
 sg13g2_fill_1 FILLER_6_932 ();
 sg13g2_fill_2 FILLER_6_959 ();
 sg13g2_fill_2 FILLER_6_1019 ();
 sg13g2_fill_1 FILLER_6_1021 ();
 sg13g2_fill_1 FILLER_6_1141 ();
 sg13g2_fill_2 FILLER_6_1168 ();
 sg13g2_fill_1 FILLER_6_1170 ();
 sg13g2_fill_2 FILLER_6_1197 ();
 sg13g2_fill_1 FILLER_6_1199 ();
 sg13g2_decap_8 FILLER_6_1359 ();
 sg13g2_fill_2 FILLER_6_1366 ();
 sg13g2_fill_2 FILLER_6_1464 ();
 sg13g2_fill_1 FILLER_6_1466 ();
 sg13g2_fill_2 FILLER_6_1498 ();
 sg13g2_fill_1 FILLER_6_1542 ();
 sg13g2_fill_1 FILLER_6_1601 ();
 sg13g2_fill_2 FILLER_6_1615 ();
 sg13g2_fill_1 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1647 ();
 sg13g2_fill_2 FILLER_6_1654 ();
 sg13g2_fill_1 FILLER_6_1660 ();
 sg13g2_decap_4 FILLER_6_1670 ();
 sg13g2_fill_1 FILLER_6_1674 ();
 sg13g2_fill_2 FILLER_6_1711 ();
 sg13g2_fill_2 FILLER_6_1783 ();
 sg13g2_fill_1 FILLER_6_1785 ();
 sg13g2_fill_2 FILLER_6_1895 ();
 sg13g2_fill_1 FILLER_6_1897 ();
 sg13g2_fill_2 FILLER_6_1985 ();
 sg13g2_fill_2 FILLER_6_2212 ();
 sg13g2_fill_2 FILLER_6_2240 ();
 sg13g2_fill_2 FILLER_6_2281 ();
 sg13g2_fill_1 FILLER_6_2309 ();
 sg13g2_fill_2 FILLER_6_2345 ();
 sg13g2_fill_1 FILLER_6_2443 ();
 sg13g2_fill_2 FILLER_6_2532 ();
 sg13g2_fill_1 FILLER_6_2534 ();
 sg13g2_fill_2 FILLER_6_2575 ();
 sg13g2_fill_1 FILLER_6_2577 ();
 sg13g2_fill_1 FILLER_6_2604 ();
 sg13g2_fill_2 FILLER_6_2632 ();
 sg13g2_fill_1 FILLER_6_2634 ();
 sg13g2_fill_2 FILLER_6_2645 ();
 sg13g2_decap_4 FILLER_6_2669 ();
 sg13g2_fill_1 FILLER_6_2673 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_62 ();
 sg13g2_fill_2 FILLER_7_69 ();
 sg13g2_fill_2 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_125 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_fill_1 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_291 ();
 sg13g2_fill_2 FILLER_7_389 ();
 sg13g2_fill_2 FILLER_7_411 ();
 sg13g2_fill_1 FILLER_7_413 ();
 sg13g2_fill_2 FILLER_7_621 ();
 sg13g2_fill_1 FILLER_7_623 ();
 sg13g2_fill_1 FILLER_7_642 ();
 sg13g2_fill_2 FILLER_7_662 ();
 sg13g2_fill_1 FILLER_7_664 ();
 sg13g2_fill_1 FILLER_7_670 ();
 sg13g2_fill_2 FILLER_7_680 ();
 sg13g2_fill_1 FILLER_7_682 ();
 sg13g2_fill_2 FILLER_7_727 ();
 sg13g2_fill_1 FILLER_7_729 ();
 sg13g2_fill_2 FILLER_7_760 ();
 sg13g2_fill_2 FILLER_7_836 ();
 sg13g2_fill_1 FILLER_7_930 ();
 sg13g2_fill_2 FILLER_7_957 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_fill_2 FILLER_7_986 ();
 sg13g2_fill_1 FILLER_7_988 ();
 sg13g2_fill_1 FILLER_7_1034 ();
 sg13g2_fill_1 FILLER_7_1066 ();
 sg13g2_fill_2 FILLER_7_1097 ();
 sg13g2_fill_1 FILLER_7_1099 ();
 sg13g2_fill_2 FILLER_7_1188 ();
 sg13g2_fill_1 FILLER_7_1195 ();
 sg13g2_fill_2 FILLER_7_1237 ();
 sg13g2_fill_1 FILLER_7_1239 ();
 sg13g2_fill_1 FILLER_7_1250 ();
 sg13g2_fill_2 FILLER_7_1335 ();
 sg13g2_fill_1 FILLER_7_1337 ();
 sg13g2_fill_2 FILLER_7_1371 ();
 sg13g2_fill_2 FILLER_7_1382 ();
 sg13g2_fill_1 FILLER_7_1425 ();
 sg13g2_fill_2 FILLER_7_1457 ();
 sg13g2_fill_2 FILLER_7_1484 ();
 sg13g2_fill_1 FILLER_7_1577 ();
 sg13g2_fill_2 FILLER_7_1624 ();
 sg13g2_fill_1 FILLER_7_1626 ();
 sg13g2_decap_4 FILLER_7_1641 ();
 sg13g2_fill_1 FILLER_7_1645 ();
 sg13g2_fill_1 FILLER_7_1682 ();
 sg13g2_fill_1 FILLER_7_1727 ();
 sg13g2_fill_2 FILLER_7_1759 ();
 sg13g2_fill_1 FILLER_7_1761 ();
 sg13g2_fill_1 FILLER_7_1797 ();
 sg13g2_fill_2 FILLER_7_1838 ();
 sg13g2_fill_1 FILLER_7_1855 ();
 sg13g2_decap_4 FILLER_7_1886 ();
 sg13g2_fill_2 FILLER_7_1890 ();
 sg13g2_fill_1 FILLER_7_1900 ();
 sg13g2_fill_2 FILLER_7_1971 ();
 sg13g2_fill_1 FILLER_7_1973 ();
 sg13g2_fill_2 FILLER_7_2000 ();
 sg13g2_fill_2 FILLER_7_2021 ();
 sg13g2_fill_1 FILLER_7_2023 ();
 sg13g2_fill_2 FILLER_7_2076 ();
 sg13g2_fill_1 FILLER_7_2078 ();
 sg13g2_fill_2 FILLER_7_2093 ();
 sg13g2_fill_1 FILLER_7_2095 ();
 sg13g2_fill_2 FILLER_7_2123 ();
 sg13g2_fill_1 FILLER_7_2144 ();
 sg13g2_decap_8 FILLER_7_2185 ();
 sg13g2_decap_4 FILLER_7_2246 ();
 sg13g2_decap_4 FILLER_7_2303 ();
 sg13g2_fill_2 FILLER_7_2329 ();
 sg13g2_fill_1 FILLER_7_2331 ();
 sg13g2_fill_2 FILLER_7_2372 ();
 sg13g2_fill_1 FILLER_7_2388 ();
 sg13g2_decap_4 FILLER_7_2411 ();
 sg13g2_fill_1 FILLER_7_2425 ();
 sg13g2_decap_4 FILLER_7_2439 ();
 sg13g2_fill_2 FILLER_7_2457 ();
 sg13g2_fill_1 FILLER_7_2459 ();
 sg13g2_fill_2 FILLER_7_2485 ();
 sg13g2_fill_1 FILLER_7_2487 ();
 sg13g2_fill_2 FILLER_7_2498 ();
 sg13g2_fill_2 FILLER_7_2551 ();
 sg13g2_fill_2 FILLER_7_2567 ();
 sg13g2_fill_1 FILLER_7_2569 ();
 sg13g2_fill_1 FILLER_7_2589 ();
 sg13g2_fill_1 FILLER_7_2630 ();
 sg13g2_decap_8 FILLER_7_2641 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_fill_2 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_138 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_2 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_2 FILLER_8_450 ();
 sg13g2_fill_1 FILLER_8_452 ();
 sg13g2_fill_2 FILLER_8_483 ();
 sg13g2_fill_1 FILLER_8_485 ();
 sg13g2_fill_2 FILLER_8_534 ();
 sg13g2_fill_1 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_588 ();
 sg13g2_fill_2 FILLER_8_631 ();
 sg13g2_fill_1 FILLER_8_633 ();
 sg13g2_fill_2 FILLER_8_700 ();
 sg13g2_fill_1 FILLER_8_716 ();
 sg13g2_fill_2 FILLER_8_739 ();
 sg13g2_fill_1 FILLER_8_741 ();
 sg13g2_fill_2 FILLER_8_774 ();
 sg13g2_fill_1 FILLER_8_776 ();
 sg13g2_fill_2 FILLER_8_847 ();
 sg13g2_fill_2 FILLER_8_884 ();
 sg13g2_fill_1 FILLER_8_886 ();
 sg13g2_fill_2 FILLER_8_937 ();
 sg13g2_fill_1 FILLER_8_939 ();
 sg13g2_fill_1 FILLER_8_960 ();
 sg13g2_fill_2 FILLER_8_1001 ();
 sg13g2_fill_1 FILLER_8_1003 ();
 sg13g2_fill_1 FILLER_8_1023 ();
 sg13g2_fill_1 FILLER_8_1038 ();
 sg13g2_fill_1 FILLER_8_1091 ();
 sg13g2_fill_1 FILLER_8_1148 ();
 sg13g2_fill_1 FILLER_8_1154 ();
 sg13g2_fill_2 FILLER_8_1357 ();
 sg13g2_fill_1 FILLER_8_1359 ();
 sg13g2_fill_2 FILLER_8_1401 ();
 sg13g2_fill_1 FILLER_8_1403 ();
 sg13g2_fill_2 FILLER_8_1448 ();
 sg13g2_fill_2 FILLER_8_1483 ();
 sg13g2_fill_1 FILLER_8_1485 ();
 sg13g2_fill_2 FILLER_8_1564 ();
 sg13g2_fill_1 FILLER_8_1566 ();
 sg13g2_fill_1 FILLER_8_1592 ();
 sg13g2_fill_1 FILLER_8_1619 ();
 sg13g2_fill_2 FILLER_8_1628 ();
 sg13g2_fill_2 FILLER_8_1647 ();
 sg13g2_fill_1 FILLER_8_1649 ();
 sg13g2_fill_1 FILLER_8_1738 ();
 sg13g2_fill_1 FILLER_8_1819 ();
 sg13g2_decap_8 FILLER_8_1872 ();
 sg13g2_fill_1 FILLER_8_1921 ();
 sg13g2_fill_2 FILLER_8_1956 ();
 sg13g2_fill_1 FILLER_8_1958 ();
 sg13g2_fill_2 FILLER_8_2030 ();
 sg13g2_fill_1 FILLER_8_2058 ();
 sg13g2_fill_2 FILLER_8_2095 ();
 sg13g2_fill_1 FILLER_8_2097 ();
 sg13g2_fill_1 FILLER_8_2124 ();
 sg13g2_fill_1 FILLER_8_2168 ();
 sg13g2_fill_1 FILLER_8_2240 ();
 sg13g2_fill_2 FILLER_8_2271 ();
 sg13g2_fill_1 FILLER_8_2273 ();
 sg13g2_fill_2 FILLER_8_2380 ();
 sg13g2_fill_2 FILLER_8_2490 ();
 sg13g2_fill_1 FILLER_8_2492 ();
 sg13g2_fill_2 FILLER_8_2547 ();
 sg13g2_fill_1 FILLER_8_2597 ();
 sg13g2_fill_2 FILLER_8_2608 ();
 sg13g2_fill_1 FILLER_8_2610 ();
 sg13g2_fill_2 FILLER_8_2671 ();
 sg13g2_fill_1 FILLER_8_2673 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_2 FILLER_9_263 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_2 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_513 ();
 sg13g2_fill_1 FILLER_9_515 ();
 sg13g2_fill_1 FILLER_9_521 ();
 sg13g2_fill_1 FILLER_9_532 ();
 sg13g2_fill_2 FILLER_9_543 ();
 sg13g2_fill_1 FILLER_9_545 ();
 sg13g2_fill_2 FILLER_9_577 ();
 sg13g2_fill_1 FILLER_9_579 ();
 sg13g2_fill_1 FILLER_9_629 ();
 sg13g2_fill_2 FILLER_9_640 ();
 sg13g2_fill_1 FILLER_9_667 ();
 sg13g2_fill_1 FILLER_9_688 ();
 sg13g2_fill_1 FILLER_9_738 ();
 sg13g2_fill_2 FILLER_9_773 ();
 sg13g2_fill_2 FILLER_9_816 ();
 sg13g2_fill_1 FILLER_9_818 ();
 sg13g2_fill_1 FILLER_9_823 ();
 sg13g2_fill_2 FILLER_9_829 ();
 sg13g2_fill_1 FILLER_9_831 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_fill_2 FILLER_9_871 ();
 sg13g2_fill_1 FILLER_9_912 ();
 sg13g2_fill_2 FILLER_9_965 ();
 sg13g2_fill_1 FILLER_9_967 ();
 sg13g2_fill_2 FILLER_9_994 ();
 sg13g2_fill_1 FILLER_9_1022 ();
 sg13g2_fill_2 FILLER_9_1049 ();
 sg13g2_fill_2 FILLER_9_1108 ();
 sg13g2_fill_1 FILLER_9_1110 ();
 sg13g2_fill_2 FILLER_9_1143 ();
 sg13g2_fill_2 FILLER_9_1266 ();
 sg13g2_fill_1 FILLER_9_1268 ();
 sg13g2_fill_1 FILLER_9_1274 ();
 sg13g2_fill_2 FILLER_9_1318 ();
 sg13g2_fill_1 FILLER_9_1335 ();
 sg13g2_decap_4 FILLER_9_1346 ();
 sg13g2_fill_2 FILLER_9_1369 ();
 sg13g2_fill_1 FILLER_9_1371 ();
 sg13g2_fill_2 FILLER_9_1441 ();
 sg13g2_decap_8 FILLER_9_1464 ();
 sg13g2_fill_2 FILLER_9_1471 ();
 sg13g2_fill_1 FILLER_9_1473 ();
 sg13g2_decap_4 FILLER_9_1489 ();
 sg13g2_fill_2 FILLER_9_1493 ();
 sg13g2_fill_2 FILLER_9_1518 ();
 sg13g2_fill_1 FILLER_9_1520 ();
 sg13g2_fill_1 FILLER_9_1534 ();
 sg13g2_fill_2 FILLER_9_1547 ();
 sg13g2_fill_2 FILLER_9_1582 ();
 sg13g2_fill_1 FILLER_9_1598 ();
 sg13g2_fill_1 FILLER_9_1608 ();
 sg13g2_fill_2 FILLER_9_1679 ();
 sg13g2_fill_2 FILLER_9_1808 ();
 sg13g2_fill_2 FILLER_9_1843 ();
 sg13g2_fill_1 FILLER_9_1845 ();
 sg13g2_decap_8 FILLER_9_1863 ();
 sg13g2_fill_1 FILLER_9_1870 ();
 sg13g2_fill_2 FILLER_9_1875 ();
 sg13g2_fill_1 FILLER_9_1877 ();
 sg13g2_fill_2 FILLER_9_1910 ();
 sg13g2_fill_1 FILLER_9_1912 ();
 sg13g2_fill_2 FILLER_9_1932 ();
 sg13g2_fill_1 FILLER_9_2025 ();
 sg13g2_fill_2 FILLER_9_2054 ();
 sg13g2_fill_1 FILLER_9_2056 ();
 sg13g2_fill_2 FILLER_9_2067 ();
 sg13g2_fill_2 FILLER_9_2149 ();
 sg13g2_fill_1 FILLER_9_2151 ();
 sg13g2_fill_1 FILLER_9_2188 ();
 sg13g2_fill_1 FILLER_9_2234 ();
 sg13g2_fill_1 FILLER_9_2268 ();
 sg13g2_fill_2 FILLER_9_2317 ();
 sg13g2_fill_2 FILLER_9_2356 ();
 sg13g2_fill_1 FILLER_9_2358 ();
 sg13g2_fill_2 FILLER_9_2415 ();
 sg13g2_fill_1 FILLER_9_2417 ();
 sg13g2_fill_1 FILLER_9_2427 ();
 sg13g2_fill_2 FILLER_9_2490 ();
 sg13g2_fill_1 FILLER_9_2492 ();
 sg13g2_fill_2 FILLER_9_2519 ();
 sg13g2_fill_1 FILLER_9_2521 ();
 sg13g2_fill_2 FILLER_9_2552 ();
 sg13g2_fill_2 FILLER_9_2639 ();
 sg13g2_fill_1 FILLER_9_2641 ();
 sg13g2_decap_4 FILLER_9_2668 ();
 sg13g2_fill_2 FILLER_9_2672 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_82 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_291 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_fill_2 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_fill_2 FILLER_10_388 ();
 sg13g2_fill_1 FILLER_10_390 ();
 sg13g2_fill_1 FILLER_10_422 ();
 sg13g2_fill_2 FILLER_10_439 ();
 sg13g2_fill_2 FILLER_10_467 ();
 sg13g2_fill_2 FILLER_10_490 ();
 sg13g2_fill_1 FILLER_10_492 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_549 ();
 sg13g2_fill_2 FILLER_10_559 ();
 sg13g2_fill_1 FILLER_10_561 ();
 sg13g2_fill_1 FILLER_10_589 ();
 sg13g2_fill_2 FILLER_10_598 ();
 sg13g2_fill_2 FILLER_10_622 ();
 sg13g2_fill_2 FILLER_10_637 ();
 sg13g2_fill_1 FILLER_10_639 ();
 sg13g2_fill_1 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_656 ();
 sg13g2_fill_1 FILLER_10_658 ();
 sg13g2_fill_2 FILLER_10_685 ();
 sg13g2_fill_1 FILLER_10_687 ();
 sg13g2_fill_2 FILLER_10_723 ();
 sg13g2_fill_1 FILLER_10_725 ();
 sg13g2_fill_2 FILLER_10_735 ();
 sg13g2_fill_1 FILLER_10_737 ();
 sg13g2_fill_1 FILLER_10_777 ();
 sg13g2_fill_2 FILLER_10_845 ();
 sg13g2_fill_1 FILLER_10_847 ();
 sg13g2_fill_1 FILLER_10_874 ();
 sg13g2_fill_1 FILLER_10_889 ();
 sg13g2_fill_1 FILLER_10_975 ();
 sg13g2_fill_1 FILLER_10_1017 ();
 sg13g2_fill_1 FILLER_10_1050 ();
 sg13g2_fill_1 FILLER_10_1078 ();
 sg13g2_fill_1 FILLER_10_1089 ();
 sg13g2_fill_1 FILLER_10_1184 ();
 sg13g2_fill_2 FILLER_10_1233 ();
 sg13g2_fill_1 FILLER_10_1235 ();
 sg13g2_fill_2 FILLER_10_1254 ();
 sg13g2_fill_1 FILLER_10_1291 ();
 sg13g2_fill_1 FILLER_10_1333 ();
 sg13g2_fill_2 FILLER_10_1352 ();
 sg13g2_fill_1 FILLER_10_1354 ();
 sg13g2_fill_1 FILLER_10_1387 ();
 sg13g2_fill_1 FILLER_10_1416 ();
 sg13g2_fill_1 FILLER_10_1425 ();
 sg13g2_fill_2 FILLER_10_1457 ();
 sg13g2_fill_2 FILLER_10_1475 ();
 sg13g2_fill_2 FILLER_10_1503 ();
 sg13g2_fill_1 FILLER_10_1505 ();
 sg13g2_fill_1 FILLER_10_1536 ();
 sg13g2_fill_1 FILLER_10_1550 ();
 sg13g2_decap_4 FILLER_10_1563 ();
 sg13g2_fill_1 FILLER_10_1567 ();
 sg13g2_fill_2 FILLER_10_1617 ();
 sg13g2_fill_2 FILLER_10_1675 ();
 sg13g2_fill_1 FILLER_10_1687 ();
 sg13g2_fill_2 FILLER_10_1701 ();
 sg13g2_fill_1 FILLER_10_1703 ();
 sg13g2_fill_2 FILLER_10_1718 ();
 sg13g2_fill_1 FILLER_10_1720 ();
 sg13g2_fill_1 FILLER_10_1771 ();
 sg13g2_fill_2 FILLER_10_1797 ();
 sg13g2_fill_1 FILLER_10_1799 ();
 sg13g2_decap_4 FILLER_10_1858 ();
 sg13g2_fill_2 FILLER_10_1862 ();
 sg13g2_fill_1 FILLER_10_1966 ();
 sg13g2_fill_1 FILLER_10_1987 ();
 sg13g2_fill_2 FILLER_10_2018 ();
 sg13g2_fill_1 FILLER_10_2088 ();
 sg13g2_fill_2 FILLER_10_2143 ();
 sg13g2_fill_1 FILLER_10_2145 ();
 sg13g2_fill_2 FILLER_10_2180 ();
 sg13g2_fill_1 FILLER_10_2182 ();
 sg13g2_decap_4 FILLER_10_2219 ();
 sg13g2_fill_1 FILLER_10_2223 ();
 sg13g2_decap_8 FILLER_10_2312 ();
 sg13g2_fill_2 FILLER_10_2319 ();
 sg13g2_fill_1 FILLER_10_2366 ();
 sg13g2_fill_2 FILLER_10_2438 ();
 sg13g2_fill_1 FILLER_10_2440 ();
 sg13g2_decap_4 FILLER_10_2457 ();
 sg13g2_fill_2 FILLER_10_2461 ();
 sg13g2_fill_1 FILLER_10_2467 ();
 sg13g2_fill_2 FILLER_10_2588 ();
 sg13g2_fill_2 FILLER_10_2671 ();
 sg13g2_fill_1 FILLER_10_2673 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_18 ();
 sg13g2_fill_1 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_435 ();
 sg13g2_fill_1 FILLER_11_474 ();
 sg13g2_fill_1 FILLER_11_490 ();
 sg13g2_fill_1 FILLER_11_496 ();
 sg13g2_fill_1 FILLER_11_507 ();
 sg13g2_fill_2 FILLER_11_539 ();
 sg13g2_fill_1 FILLER_11_541 ();
 sg13g2_fill_2 FILLER_11_550 ();
 sg13g2_fill_1 FILLER_11_552 ();
 sg13g2_fill_2 FILLER_11_568 ();
 sg13g2_fill_1 FILLER_11_570 ();
 sg13g2_fill_1 FILLER_11_589 ();
 sg13g2_fill_2 FILLER_11_616 ();
 sg13g2_fill_2 FILLER_11_629 ();
 sg13g2_fill_1 FILLER_11_631 ();
 sg13g2_fill_1 FILLER_11_668 ();
 sg13g2_fill_2 FILLER_11_689 ();
 sg13g2_fill_1 FILLER_11_696 ();
 sg13g2_fill_2 FILLER_11_703 ();
 sg13g2_fill_1 FILLER_11_705 ();
 sg13g2_fill_1 FILLER_11_737 ();
 sg13g2_fill_1 FILLER_11_764 ();
 sg13g2_fill_1 FILLER_11_818 ();
 sg13g2_fill_2 FILLER_11_833 ();
 sg13g2_fill_2 FILLER_11_850 ();
 sg13g2_fill_2 FILLER_11_958 ();
 sg13g2_fill_2 FILLER_11_995 ();
 sg13g2_fill_1 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1029 ();
 sg13g2_fill_2 FILLER_11_1122 ();
 sg13g2_fill_1 FILLER_11_1124 ();
 sg13g2_fill_1 FILLER_11_1161 ();
 sg13g2_fill_1 FILLER_11_1229 ();
 sg13g2_fill_2 FILLER_11_1235 ();
 sg13g2_fill_1 FILLER_11_1237 ();
 sg13g2_fill_2 FILLER_11_1255 ();
 sg13g2_fill_1 FILLER_11_1257 ();
 sg13g2_fill_2 FILLER_11_1284 ();
 sg13g2_fill_1 FILLER_11_1286 ();
 sg13g2_fill_2 FILLER_11_1297 ();
 sg13g2_fill_1 FILLER_11_1299 ();
 sg13g2_fill_2 FILLER_11_1305 ();
 sg13g2_fill_2 FILLER_11_1320 ();
 sg13g2_decap_8 FILLER_11_1330 ();
 sg13g2_decap_4 FILLER_11_1337 ();
 sg13g2_fill_1 FILLER_11_1368 ();
 sg13g2_decap_8 FILLER_11_1381 ();
 sg13g2_decap_8 FILLER_11_1388 ();
 sg13g2_fill_1 FILLER_11_1395 ();
 sg13g2_fill_2 FILLER_11_1406 ();
 sg13g2_fill_1 FILLER_11_1408 ();
 sg13g2_fill_2 FILLER_11_1418 ();
 sg13g2_fill_1 FILLER_11_1420 ();
 sg13g2_fill_1 FILLER_11_1430 ();
 sg13g2_fill_2 FILLER_11_1443 ();
 sg13g2_fill_2 FILLER_11_1451 ();
 sg13g2_fill_2 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1507 ();
 sg13g2_fill_2 FILLER_11_1530 ();
 sg13g2_fill_1 FILLER_11_1532 ();
 sg13g2_fill_1 FILLER_11_1537 ();
 sg13g2_decap_8 FILLER_11_1542 ();
 sg13g2_decap_8 FILLER_11_1579 ();
 sg13g2_decap_8 FILLER_11_1586 ();
 sg13g2_decap_4 FILLER_11_1593 ();
 sg13g2_fill_1 FILLER_11_1597 ();
 sg13g2_decap_4 FILLER_11_1606 ();
 sg13g2_fill_2 FILLER_11_1629 ();
 sg13g2_fill_1 FILLER_11_1644 ();
 sg13g2_decap_4 FILLER_11_1671 ();
 sg13g2_fill_1 FILLER_11_1675 ();
 sg13g2_fill_1 FILLER_11_1721 ();
 sg13g2_fill_2 FILLER_11_1842 ();
 sg13g2_fill_1 FILLER_11_1853 ();
 sg13g2_fill_1 FILLER_11_1880 ();
 sg13g2_fill_1 FILLER_11_1939 ();
 sg13g2_fill_1 FILLER_11_1949 ();
 sg13g2_fill_2 FILLER_11_1968 ();
 sg13g2_fill_1 FILLER_11_1970 ();
 sg13g2_fill_2 FILLER_11_2001 ();
 sg13g2_fill_1 FILLER_11_2003 ();
 sg13g2_fill_2 FILLER_11_2039 ();
 sg13g2_fill_1 FILLER_11_2041 ();
 sg13g2_fill_2 FILLER_11_2050 ();
 sg13g2_fill_1 FILLER_11_2052 ();
 sg13g2_fill_2 FILLER_11_2066 ();
 sg13g2_fill_1 FILLER_11_2068 ();
 sg13g2_fill_1 FILLER_11_2092 ();
 sg13g2_fill_1 FILLER_11_2130 ();
 sg13g2_fill_1 FILLER_11_2189 ();
 sg13g2_decap_4 FILLER_11_2232 ();
 sg13g2_fill_1 FILLER_11_2236 ();
 sg13g2_fill_2 FILLER_11_2256 ();
 sg13g2_fill_1 FILLER_11_2311 ();
 sg13g2_fill_2 FILLER_11_2352 ();
 sg13g2_fill_2 FILLER_11_2415 ();
 sg13g2_fill_1 FILLER_11_2417 ();
 sg13g2_fill_2 FILLER_11_2424 ();
 sg13g2_fill_1 FILLER_11_2426 ();
 sg13g2_fill_1 FILLER_11_2478 ();
 sg13g2_fill_2 FILLER_11_2519 ();
 sg13g2_fill_1 FILLER_11_2521 ();
 sg13g2_fill_2 FILLER_11_2557 ();
 sg13g2_fill_1 FILLER_11_2595 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_260 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_fill_1 FILLER_12_328 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_fill_2 FILLER_12_372 ();
 sg13g2_fill_1 FILLER_12_434 ();
 sg13g2_fill_1 FILLER_12_448 ();
 sg13g2_fill_2 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_12_479 ();
 sg13g2_fill_1 FILLER_12_486 ();
 sg13g2_fill_2 FILLER_12_619 ();
 sg13g2_fill_2 FILLER_12_640 ();
 sg13g2_fill_1 FILLER_12_662 ();
 sg13g2_fill_2 FILLER_12_699 ();
 sg13g2_fill_1 FILLER_12_742 ();
 sg13g2_fill_1 FILLER_12_774 ();
 sg13g2_fill_1 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_852 ();
 sg13g2_fill_2 FILLER_12_867 ();
 sg13g2_fill_1 FILLER_12_869 ();
 sg13g2_fill_1 FILLER_12_889 ();
 sg13g2_fill_1 FILLER_12_899 ();
 sg13g2_fill_2 FILLER_12_936 ();
 sg13g2_fill_1 FILLER_12_938 ();
 sg13g2_fill_1 FILLER_12_969 ();
 sg13g2_fill_1 FILLER_12_995 ();
 sg13g2_fill_2 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1041 ();
 sg13g2_fill_2 FILLER_12_1080 ();
 sg13g2_fill_1 FILLER_12_1082 ();
 sg13g2_fill_2 FILLER_12_1087 ();
 sg13g2_fill_2 FILLER_12_1107 ();
 sg13g2_fill_2 FILLER_12_1132 ();
 sg13g2_fill_1 FILLER_12_1134 ();
 sg13g2_fill_1 FILLER_12_1170 ();
 sg13g2_fill_2 FILLER_12_1188 ();
 sg13g2_fill_1 FILLER_12_1239 ();
 sg13g2_fill_2 FILLER_12_1278 ();
 sg13g2_fill_2 FILLER_12_1330 ();
 sg13g2_fill_1 FILLER_12_1332 ();
 sg13g2_decap_8 FILLER_12_1390 ();
 sg13g2_decap_8 FILLER_12_1397 ();
 sg13g2_fill_2 FILLER_12_1426 ();
 sg13g2_fill_2 FILLER_12_1451 ();
 sg13g2_fill_1 FILLER_12_1453 ();
 sg13g2_fill_2 FILLER_12_1469 ();
 sg13g2_fill_1 FILLER_12_1475 ();
 sg13g2_decap_4 FILLER_12_1484 ();
 sg13g2_decap_8 FILLER_12_1516 ();
 sg13g2_decap_4 FILLER_12_1523 ();
 sg13g2_fill_1 FILLER_12_1527 ();
 sg13g2_fill_1 FILLER_12_1554 ();
 sg13g2_fill_2 FILLER_12_1568 ();
 sg13g2_fill_1 FILLER_12_1570 ();
 sg13g2_fill_2 FILLER_12_1576 ();
 sg13g2_fill_1 FILLER_12_1578 ();
 sg13g2_fill_1 FILLER_12_1583 ();
 sg13g2_decap_4 FILLER_12_1594 ();
 sg13g2_fill_1 FILLER_12_1598 ();
 sg13g2_decap_4 FILLER_12_1609 ();
 sg13g2_fill_1 FILLER_12_1621 ();
 sg13g2_fill_2 FILLER_12_1627 ();
 sg13g2_decap_8 FILLER_12_1637 ();
 sg13g2_decap_4 FILLER_12_1644 ();
 sg13g2_fill_1 FILLER_12_1648 ();
 sg13g2_fill_2 FILLER_12_1679 ();
 sg13g2_fill_1 FILLER_12_1691 ();
 sg13g2_fill_1 FILLER_12_1755 ();
 sg13g2_fill_2 FILLER_12_1765 ();
 sg13g2_fill_2 FILLER_12_1840 ();
 sg13g2_fill_1 FILLER_12_1842 ();
 sg13g2_fill_1 FILLER_12_1921 ();
 sg13g2_fill_2 FILLER_12_1962 ();
 sg13g2_fill_1 FILLER_12_1964 ();
 sg13g2_fill_2 FILLER_12_1991 ();
 sg13g2_fill_2 FILLER_12_2019 ();
 sg13g2_fill_1 FILLER_12_2061 ();
 sg13g2_fill_1 FILLER_12_2113 ();
 sg13g2_fill_1 FILLER_12_2142 ();
 sg13g2_fill_2 FILLER_12_2176 ();
 sg13g2_fill_1 FILLER_12_2178 ();
 sg13g2_decap_4 FILLER_12_2221 ();
 sg13g2_fill_2 FILLER_12_2225 ();
 sg13g2_fill_2 FILLER_12_2283 ();
 sg13g2_decap_4 FILLER_12_2333 ();
 sg13g2_fill_1 FILLER_12_2337 ();
 sg13g2_fill_1 FILLER_12_2387 ();
 sg13g2_fill_1 FILLER_12_2424 ();
 sg13g2_fill_1 FILLER_12_2440 ();
 sg13g2_fill_1 FILLER_12_2451 ();
 sg13g2_fill_1 FILLER_12_2548 ();
 sg13g2_fill_2 FILLER_12_2563 ();
 sg13g2_fill_1 FILLER_12_2596 ();
 sg13g2_fill_2 FILLER_12_2629 ();
 sg13g2_fill_2 FILLER_12_2649 ();
 sg13g2_fill_1 FILLER_12_2673 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_396 ();
 sg13g2_fill_1 FILLER_13_434 ();
 sg13g2_fill_2 FILLER_13_471 ();
 sg13g2_fill_2 FILLER_13_486 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_fill_2 FILLER_13_504 ();
 sg13g2_fill_2 FILLER_13_586 ();
 sg13g2_fill_1 FILLER_13_588 ();
 sg13g2_fill_2 FILLER_13_673 ();
 sg13g2_fill_1 FILLER_13_675 ();
 sg13g2_fill_2 FILLER_13_696 ();
 sg13g2_fill_1 FILLER_13_698 ();
 sg13g2_fill_1 FILLER_13_717 ();
 sg13g2_fill_2 FILLER_13_760 ();
 sg13g2_fill_2 FILLER_13_784 ();
 sg13g2_fill_1 FILLER_13_797 ();
 sg13g2_fill_2 FILLER_13_807 ();
 sg13g2_fill_2 FILLER_13_822 ();
 sg13g2_fill_1 FILLER_13_853 ();
 sg13g2_fill_2 FILLER_13_921 ();
 sg13g2_fill_2 FILLER_13_960 ();
 sg13g2_fill_2 FILLER_13_1059 ();
 sg13g2_fill_1 FILLER_13_1087 ();
 sg13g2_fill_1 FILLER_13_1105 ();
 sg13g2_fill_2 FILLER_13_1112 ();
 sg13g2_fill_2 FILLER_13_1140 ();
 sg13g2_fill_2 FILLER_13_1172 ();
 sg13g2_fill_1 FILLER_13_1174 ();
 sg13g2_fill_2 FILLER_13_1215 ();
 sg13g2_fill_2 FILLER_13_1263 ();
 sg13g2_fill_1 FILLER_13_1300 ();
 sg13g2_fill_1 FILLER_13_1309 ();
 sg13g2_decap_8 FILLER_13_1314 ();
 sg13g2_decap_4 FILLER_13_1321 ();
 sg13g2_fill_1 FILLER_13_1325 ();
 sg13g2_decap_4 FILLER_13_1336 ();
 sg13g2_fill_2 FILLER_13_1340 ();
 sg13g2_fill_1 FILLER_13_1409 ();
 sg13g2_decap_4 FILLER_13_1414 ();
 sg13g2_fill_1 FILLER_13_1426 ();
 sg13g2_decap_8 FILLER_13_1437 ();
 sg13g2_decap_4 FILLER_13_1444 ();
 sg13g2_fill_2 FILLER_13_1465 ();
 sg13g2_decap_4 FILLER_13_1493 ();
 sg13g2_fill_2 FILLER_13_1518 ();
 sg13g2_fill_2 FILLER_13_1528 ();
 sg13g2_fill_2 FILLER_13_1540 ();
 sg13g2_fill_2 FILLER_13_1550 ();
 sg13g2_fill_1 FILLER_13_1577 ();
 sg13g2_fill_2 FILLER_13_1666 ();
 sg13g2_fill_1 FILLER_13_1668 ();
 sg13g2_fill_1 FILLER_13_1683 ();
 sg13g2_fill_2 FILLER_13_1728 ();
 sg13g2_fill_2 FILLER_13_1790 ();
 sg13g2_fill_1 FILLER_13_1792 ();
 sg13g2_fill_1 FILLER_13_1833 ();
 sg13g2_fill_1 FILLER_13_1934 ();
 sg13g2_fill_2 FILLER_13_1963 ();
 sg13g2_fill_1 FILLER_13_1965 ();
 sg13g2_fill_2 FILLER_13_1998 ();
 sg13g2_fill_1 FILLER_13_2000 ();
 sg13g2_fill_1 FILLER_13_2045 ();
 sg13g2_fill_1 FILLER_13_2084 ();
 sg13g2_decap_4 FILLER_13_2098 ();
 sg13g2_fill_1 FILLER_13_2102 ();
 sg13g2_fill_2 FILLER_13_2157 ();
 sg13g2_fill_2 FILLER_13_2185 ();
 sg13g2_fill_1 FILLER_13_2187 ();
 sg13g2_fill_1 FILLER_13_2198 ();
 sg13g2_decap_4 FILLER_13_2218 ();
 sg13g2_fill_2 FILLER_13_2232 ();
 sg13g2_fill_1 FILLER_13_2234 ();
 sg13g2_fill_1 FILLER_13_2254 ();
 sg13g2_fill_1 FILLER_13_2278 ();
 sg13g2_fill_2 FILLER_13_2288 ();
 sg13g2_fill_2 FILLER_13_2304 ();
 sg13g2_decap_8 FILLER_13_2332 ();
 sg13g2_fill_2 FILLER_13_2339 ();
 sg13g2_fill_1 FILLER_13_2412 ();
 sg13g2_fill_2 FILLER_13_2448 ();
 sg13g2_fill_1 FILLER_13_2450 ();
 sg13g2_fill_2 FILLER_13_2486 ();
 sg13g2_fill_1 FILLER_13_2488 ();
 sg13g2_fill_2 FILLER_13_2515 ();
 sg13g2_fill_1 FILLER_13_2517 ();
 sg13g2_fill_1 FILLER_13_2673 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_91 ();
 sg13g2_fill_1 FILLER_14_93 ();
 sg13g2_fill_1 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_466 ();
 sg13g2_fill_1 FILLER_14_583 ();
 sg13g2_fill_2 FILLER_14_593 ();
 sg13g2_fill_1 FILLER_14_595 ();
 sg13g2_fill_2 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_617 ();
 sg13g2_fill_2 FILLER_14_638 ();
 sg13g2_fill_2 FILLER_14_650 ();
 sg13g2_fill_1 FILLER_14_652 ();
 sg13g2_fill_2 FILLER_14_687 ();
 sg13g2_fill_1 FILLER_14_720 ();
 sg13g2_fill_2 FILLER_14_776 ();
 sg13g2_fill_1 FILLER_14_786 ();
 sg13g2_fill_2 FILLER_14_813 ();
 sg13g2_fill_1 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_862 ();
 sg13g2_fill_1 FILLER_14_883 ();
 sg13g2_fill_2 FILLER_14_897 ();
 sg13g2_fill_1 FILLER_14_899 ();
 sg13g2_fill_1 FILLER_14_913 ();
 sg13g2_fill_2 FILLER_14_963 ();
 sg13g2_fill_2 FILLER_14_1025 ();
 sg13g2_fill_2 FILLER_14_1054 ();
 sg13g2_fill_1 FILLER_14_1056 ();
 sg13g2_fill_2 FILLER_14_1070 ();
 sg13g2_fill_1 FILLER_14_1172 ();
 sg13g2_fill_2 FILLER_14_1181 ();
 sg13g2_fill_1 FILLER_14_1183 ();
 sg13g2_fill_2 FILLER_14_1236 ();
 sg13g2_fill_1 FILLER_14_1238 ();
 sg13g2_fill_2 FILLER_14_1273 ();
 sg13g2_fill_1 FILLER_14_1275 ();
 sg13g2_fill_2 FILLER_14_1280 ();
 sg13g2_fill_1 FILLER_14_1282 ();
 sg13g2_decap_8 FILLER_14_1287 ();
 sg13g2_fill_2 FILLER_14_1304 ();
 sg13g2_fill_2 FILLER_14_1310 ();
 sg13g2_fill_1 FILLER_14_1338 ();
 sg13g2_decap_8 FILLER_14_1395 ();
 sg13g2_fill_2 FILLER_14_1402 ();
 sg13g2_fill_1 FILLER_14_1428 ();
 sg13g2_fill_1 FILLER_14_1435 ();
 sg13g2_fill_2 FILLER_14_1455 ();
 sg13g2_decap_8 FILLER_14_1465 ();
 sg13g2_decap_8 FILLER_14_1472 ();
 sg13g2_fill_2 FILLER_14_1479 ();
 sg13g2_fill_1 FILLER_14_1481 ();
 sg13g2_fill_2 FILLER_14_1499 ();
 sg13g2_fill_2 FILLER_14_1523 ();
 sg13g2_fill_1 FILLER_14_1525 ();
 sg13g2_fill_2 FILLER_14_1539 ();
 sg13g2_fill_2 FILLER_14_1549 ();
 sg13g2_fill_1 FILLER_14_1559 ();
 sg13g2_fill_1 FILLER_14_1569 ();
 sg13g2_decap_4 FILLER_14_1579 ();
 sg13g2_fill_1 FILLER_14_1587 ();
 sg13g2_fill_1 FILLER_14_1645 ();
 sg13g2_fill_2 FILLER_14_1656 ();
 sg13g2_fill_2 FILLER_14_1697 ();
 sg13g2_fill_2 FILLER_14_1787 ();
 sg13g2_fill_2 FILLER_14_1829 ();
 sg13g2_fill_1 FILLER_14_1831 ();
 sg13g2_fill_2 FILLER_14_1917 ();
 sg13g2_fill_1 FILLER_14_1919 ();
 sg13g2_fill_2 FILLER_14_1972 ();
 sg13g2_fill_1 FILLER_14_2000 ();
 sg13g2_fill_1 FILLER_14_2033 ();
 sg13g2_fill_1 FILLER_14_2054 ();
 sg13g2_fill_2 FILLER_14_2069 ();
 sg13g2_fill_1 FILLER_14_2071 ();
 sg13g2_fill_2 FILLER_14_2082 ();
 sg13g2_fill_1 FILLER_14_2084 ();
 sg13g2_decap_4 FILLER_14_2112 ();
 sg13g2_fill_2 FILLER_14_2116 ();
 sg13g2_fill_1 FILLER_14_2173 ();
 sg13g2_fill_2 FILLER_14_2307 ();
 sg13g2_fill_2 FILLER_14_2326 ();
 sg13g2_fill_1 FILLER_14_2351 ();
 sg13g2_fill_1 FILLER_14_2415 ();
 sg13g2_fill_1 FILLER_14_2559 ();
 sg13g2_fill_2 FILLER_14_2564 ();
 sg13g2_fill_1 FILLER_14_2576 ();
 sg13g2_fill_1 FILLER_14_2641 ();
 sg13g2_fill_2 FILLER_14_2672 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_2 FILLER_15_29 ();
 sg13g2_fill_1 FILLER_15_41 ();
 sg13g2_fill_2 FILLER_15_104 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_302 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_330 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_fill_1 FILLER_15_391 ();
 sg13g2_fill_2 FILLER_15_441 ();
 sg13g2_fill_1 FILLER_15_473 ();
 sg13g2_fill_1 FILLER_15_487 ();
 sg13g2_fill_1 FILLER_15_502 ();
 sg13g2_fill_1 FILLER_15_517 ();
 sg13g2_fill_2 FILLER_15_629 ();
 sg13g2_fill_2 FILLER_15_713 ();
 sg13g2_fill_2 FILLER_15_720 ();
 sg13g2_fill_1 FILLER_15_722 ();
 sg13g2_fill_2 FILLER_15_796 ();
 sg13g2_fill_2 FILLER_15_811 ();
 sg13g2_fill_1 FILLER_15_813 ();
 sg13g2_fill_2 FILLER_15_828 ();
 sg13g2_fill_2 FILLER_15_839 ();
 sg13g2_fill_1 FILLER_15_841 ();
 sg13g2_fill_2 FILLER_15_884 ();
 sg13g2_fill_1 FILLER_15_886 ();
 sg13g2_fill_1 FILLER_15_950 ();
 sg13g2_fill_1 FILLER_15_1000 ();
 sg13g2_fill_2 FILLER_15_1016 ();
 sg13g2_fill_1 FILLER_15_1018 ();
 sg13g2_fill_1 FILLER_15_1038 ();
 sg13g2_fill_2 FILLER_15_1048 ();
 sg13g2_fill_2 FILLER_15_1098 ();
 sg13g2_fill_1 FILLER_15_1100 ();
 sg13g2_fill_2 FILLER_15_1144 ();
 sg13g2_fill_1 FILLER_15_1146 ();
 sg13g2_fill_1 FILLER_15_1161 ();
 sg13g2_fill_2 FILLER_15_1217 ();
 sg13g2_fill_1 FILLER_15_1219 ();
 sg13g2_fill_1 FILLER_15_1326 ();
 sg13g2_fill_2 FILLER_15_1336 ();
 sg13g2_decap_8 FILLER_15_1361 ();
 sg13g2_fill_2 FILLER_15_1368 ();
 sg13g2_fill_2 FILLER_15_1409 ();
 sg13g2_decap_4 FILLER_15_1419 ();
 sg13g2_fill_1 FILLER_15_1427 ();
 sg13g2_fill_1 FILLER_15_1433 ();
 sg13g2_fill_1 FILLER_15_1449 ();
 sg13g2_fill_2 FILLER_15_1454 ();
 sg13g2_fill_1 FILLER_15_1456 ();
 sg13g2_decap_4 FILLER_15_1480 ();
 sg13g2_fill_2 FILLER_15_1500 ();
 sg13g2_decap_4 FILLER_15_1533 ();
 sg13g2_fill_1 FILLER_15_1537 ();
 sg13g2_decap_8 FILLER_15_1553 ();
 sg13g2_decap_8 FILLER_15_1560 ();
 sg13g2_fill_2 FILLER_15_1614 ();
 sg13g2_fill_1 FILLER_15_1642 ();
 sg13g2_fill_2 FILLER_15_1679 ();
 sg13g2_fill_1 FILLER_15_1681 ();
 sg13g2_fill_2 FILLER_15_1701 ();
 sg13g2_fill_1 FILLER_15_1713 ();
 sg13g2_fill_2 FILLER_15_1748 ();
 sg13g2_fill_2 FILLER_15_1763 ();
 sg13g2_fill_1 FILLER_15_1765 ();
 sg13g2_fill_1 FILLER_15_1822 ();
 sg13g2_fill_2 FILLER_15_1850 ();
 sg13g2_fill_2 FILLER_15_1879 ();
 sg13g2_fill_1 FILLER_15_1881 ();
 sg13g2_fill_2 FILLER_15_1907 ();
 sg13g2_fill_1 FILLER_15_1909 ();
 sg13g2_fill_2 FILLER_15_1946 ();
 sg13g2_fill_2 FILLER_15_1988 ();
 sg13g2_fill_1 FILLER_15_1990 ();
 sg13g2_fill_2 FILLER_15_2025 ();
 sg13g2_fill_1 FILLER_15_2027 ();
 sg13g2_fill_1 FILLER_15_2156 ();
 sg13g2_fill_1 FILLER_15_2163 ();
 sg13g2_fill_1 FILLER_15_2193 ();
 sg13g2_fill_1 FILLER_15_2269 ();
 sg13g2_fill_2 FILLER_15_2291 ();
 sg13g2_decap_4 FILLER_15_2363 ();
 sg13g2_decap_4 FILLER_15_2424 ();
 sg13g2_fill_2 FILLER_15_2428 ();
 sg13g2_fill_1 FILLER_15_2436 ();
 sg13g2_fill_2 FILLER_15_2470 ();
 sg13g2_fill_1 FILLER_15_2476 ();
 sg13g2_fill_1 FILLER_15_2521 ();
 sg13g2_fill_2 FILLER_15_2586 ();
 sg13g2_fill_1 FILLER_15_2588 ();
 sg13g2_fill_2 FILLER_15_2617 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_27 ();
 sg13g2_fill_1 FILLER_16_29 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_2 FILLER_16_454 ();
 sg13g2_fill_2 FILLER_16_474 ();
 sg13g2_fill_1 FILLER_16_490 ();
 sg13g2_fill_2 FILLER_16_538 ();
 sg13g2_fill_2 FILLER_16_566 ();
 sg13g2_fill_1 FILLER_16_568 ();
 sg13g2_fill_2 FILLER_16_590 ();
 sg13g2_fill_1 FILLER_16_592 ();
 sg13g2_fill_1 FILLER_16_616 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_2 FILLER_16_710 ();
 sg13g2_fill_1 FILLER_16_752 ();
 sg13g2_fill_1 FILLER_16_848 ();
 sg13g2_fill_2 FILLER_16_904 ();
 sg13g2_fill_1 FILLER_16_906 ();
 sg13g2_fill_2 FILLER_16_956 ();
 sg13g2_fill_2 FILLER_16_963 ();
 sg13g2_fill_1 FILLER_16_965 ();
 sg13g2_fill_2 FILLER_16_975 ();
 sg13g2_fill_1 FILLER_16_977 ();
 sg13g2_fill_1 FILLER_16_1013 ();
 sg13g2_fill_1 FILLER_16_1118 ();
 sg13g2_fill_2 FILLER_16_1173 ();
 sg13g2_fill_2 FILLER_16_1198 ();
 sg13g2_fill_2 FILLER_16_1245 ();
 sg13g2_fill_2 FILLER_16_1297 ();
 sg13g2_fill_1 FILLER_16_1325 ();
 sg13g2_fill_2 FILLER_16_1330 ();
 sg13g2_fill_1 FILLER_16_1332 ();
 sg13g2_fill_2 FILLER_16_1338 ();
 sg13g2_fill_1 FILLER_16_1340 ();
 sg13g2_fill_1 FILLER_16_1350 ();
 sg13g2_fill_2 FILLER_16_1356 ();
 sg13g2_fill_1 FILLER_16_1358 ();
 sg13g2_fill_2 FILLER_16_1371 ();
 sg13g2_fill_1 FILLER_16_1373 ();
 sg13g2_fill_2 FILLER_16_1392 ();
 sg13g2_fill_2 FILLER_16_1467 ();
 sg13g2_fill_1 FILLER_16_1469 ();
 sg13g2_fill_2 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1494 ();
 sg13g2_decap_4 FILLER_16_1501 ();
 sg13g2_fill_2 FILLER_16_1523 ();
 sg13g2_fill_1 FILLER_16_1549 ();
 sg13g2_fill_2 FILLER_16_1590 ();
 sg13g2_fill_2 FILLER_16_1601 ();
 sg13g2_decap_4 FILLER_16_1618 ();
 sg13g2_fill_1 FILLER_16_1622 ();
 sg13g2_decap_8 FILLER_16_1635 ();
 sg13g2_fill_2 FILLER_16_1642 ();
 sg13g2_fill_2 FILLER_16_1777 ();
 sg13g2_fill_1 FILLER_16_1779 ();
 sg13g2_fill_2 FILLER_16_1797 ();
 sg13g2_fill_1 FILLER_16_1809 ();
 sg13g2_decap_4 FILLER_16_1842 ();
 sg13g2_fill_1 FILLER_16_1846 ();
 sg13g2_fill_1 FILLER_16_1890 ();
 sg13g2_fill_1 FILLER_16_1987 ();
 sg13g2_fill_1 FILLER_16_2042 ();
 sg13g2_fill_2 FILLER_16_2075 ();
 sg13g2_fill_2 FILLER_16_2091 ();
 sg13g2_fill_1 FILLER_16_2093 ();
 sg13g2_fill_2 FILLER_16_2136 ();
 sg13g2_fill_1 FILLER_16_2253 ();
 sg13g2_fill_2 FILLER_16_2322 ();
 sg13g2_fill_2 FILLER_16_2379 ();
 sg13g2_fill_1 FILLER_16_2381 ();
 sg13g2_decap_4 FILLER_16_2412 ();
 sg13g2_fill_2 FILLER_16_2416 ();
 sg13g2_fill_2 FILLER_16_2424 ();
 sg13g2_fill_1 FILLER_16_2426 ();
 sg13g2_fill_2 FILLER_16_2489 ();
 sg13g2_fill_1 FILLER_16_2496 ();
 sg13g2_fill_2 FILLER_16_2510 ();
 sg13g2_fill_2 FILLER_16_2580 ();
 sg13g2_fill_1 FILLER_16_2582 ();
 sg13g2_fill_1 FILLER_16_2623 ();
 sg13g2_fill_1 FILLER_16_2637 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_44 ();
 sg13g2_fill_2 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_284 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_fill_2 FILLER_17_402 ();
 sg13g2_fill_1 FILLER_17_410 ();
 sg13g2_fill_2 FILLER_17_450 ();
 sg13g2_fill_2 FILLER_17_624 ();
 sg13g2_fill_1 FILLER_17_626 ();
 sg13g2_fill_1 FILLER_17_639 ();
 sg13g2_fill_1 FILLER_17_659 ();
 sg13g2_fill_2 FILLER_17_720 ();
 sg13g2_fill_1 FILLER_17_728 ();
 sg13g2_fill_1 FILLER_17_738 ();
 sg13g2_fill_2 FILLER_17_789 ();
 sg13g2_fill_1 FILLER_17_831 ();
 sg13g2_fill_2 FILLER_17_837 ();
 sg13g2_fill_2 FILLER_17_848 ();
 sg13g2_fill_1 FILLER_17_850 ();
 sg13g2_fill_1 FILLER_17_911 ();
 sg13g2_fill_2 FILLER_17_952 ();
 sg13g2_fill_1 FILLER_17_954 ();
 sg13g2_fill_1 FILLER_17_965 ();
 sg13g2_fill_1 FILLER_17_996 ();
 sg13g2_fill_2 FILLER_17_1019 ();
 sg13g2_fill_2 FILLER_17_1064 ();
 sg13g2_fill_1 FILLER_17_1066 ();
 sg13g2_fill_2 FILLER_17_1076 ();
 sg13g2_fill_1 FILLER_17_1078 ();
 sg13g2_fill_1 FILLER_17_1104 ();
 sg13g2_fill_1 FILLER_17_1121 ();
 sg13g2_fill_2 FILLER_17_1154 ();
 sg13g2_fill_2 FILLER_17_1165 ();
 sg13g2_fill_1 FILLER_17_1181 ();
 sg13g2_fill_2 FILLER_17_1208 ();
 sg13g2_fill_1 FILLER_17_1210 ();
 sg13g2_fill_1 FILLER_17_1220 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_fill_2 FILLER_17_1279 ();
 sg13g2_fill_1 FILLER_17_1281 ();
 sg13g2_fill_1 FILLER_17_1303 ();
 sg13g2_fill_2 FILLER_17_1312 ();
 sg13g2_fill_1 FILLER_17_1314 ();
 sg13g2_fill_2 FILLER_17_1370 ();
 sg13g2_fill_2 FILLER_17_1392 ();
 sg13g2_fill_1 FILLER_17_1394 ();
 sg13g2_decap_4 FILLER_17_1421 ();
 sg13g2_fill_1 FILLER_17_1438 ();
 sg13g2_fill_1 FILLER_17_1447 ();
 sg13g2_fill_2 FILLER_17_1457 ();
 sg13g2_fill_2 FILLER_17_1464 ();
 sg13g2_fill_1 FILLER_17_1466 ();
 sg13g2_fill_2 FILLER_17_1476 ();
 sg13g2_fill_1 FILLER_17_1478 ();
 sg13g2_decap_4 FILLER_17_1485 ();
 sg13g2_fill_1 FILLER_17_1489 ();
 sg13g2_decap_4 FILLER_17_1498 ();
 sg13g2_fill_2 FILLER_17_1502 ();
 sg13g2_fill_2 FILLER_17_1536 ();
 sg13g2_fill_1 FILLER_17_1538 ();
 sg13g2_fill_2 FILLER_17_1556 ();
 sg13g2_decap_4 FILLER_17_1571 ();
 sg13g2_fill_2 FILLER_17_1580 ();
 sg13g2_fill_1 FILLER_17_1582 ();
 sg13g2_fill_2 FILLER_17_1596 ();
 sg13g2_fill_2 FILLER_17_1616 ();
 sg13g2_fill_1 FILLER_17_1618 ();
 sg13g2_fill_2 FILLER_17_1655 ();
 sg13g2_fill_1 FILLER_17_1680 ();
 sg13g2_fill_2 FILLER_17_1702 ();
 sg13g2_fill_2 FILLER_17_1748 ();
 sg13g2_fill_1 FILLER_17_1750 ();
 sg13g2_fill_2 FILLER_17_1849 ();
 sg13g2_fill_1 FILLER_17_1851 ();
 sg13g2_decap_4 FILLER_17_1856 ();
 sg13g2_fill_1 FILLER_17_1860 ();
 sg13g2_decap_4 FILLER_17_1869 ();
 sg13g2_fill_2 FILLER_17_1879 ();
 sg13g2_fill_1 FILLER_17_1881 ();
 sg13g2_fill_2 FILLER_17_1961 ();
 sg13g2_fill_1 FILLER_17_1963 ();
 sg13g2_fill_2 FILLER_17_2017 ();
 sg13g2_fill_2 FILLER_17_2071 ();
 sg13g2_fill_1 FILLER_17_2073 ();
 sg13g2_fill_2 FILLER_17_2118 ();
 sg13g2_decap_4 FILLER_17_2124 ();
 sg13g2_fill_1 FILLER_17_2128 ();
 sg13g2_fill_2 FILLER_17_2168 ();
 sg13g2_fill_1 FILLER_17_2170 ();
 sg13g2_decap_4 FILLER_17_2234 ();
 sg13g2_fill_1 FILLER_17_2362 ();
 sg13g2_fill_1 FILLER_17_2407 ();
 sg13g2_decap_4 FILLER_17_2444 ();
 sg13g2_fill_2 FILLER_17_2512 ();
 sg13g2_fill_2 FILLER_17_2546 ();
 sg13g2_fill_1 FILLER_17_2548 ();
 sg13g2_fill_2 FILLER_17_2581 ();
 sg13g2_fill_2 FILLER_17_2595 ();
 sg13g2_fill_2 FILLER_17_2628 ();
 sg13g2_fill_2 FILLER_17_2651 ();
 sg13g2_fill_1 FILLER_17_2653 ();
 sg13g2_fill_2 FILLER_17_2671 ();
 sg13g2_fill_1 FILLER_17_2673 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_30 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_389 ();
 sg13g2_fill_1 FILLER_18_517 ();
 sg13g2_fill_2 FILLER_18_529 ();
 sg13g2_fill_1 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_537 ();
 sg13g2_fill_2 FILLER_18_547 ();
 sg13g2_fill_1 FILLER_18_549 ();
 sg13g2_fill_2 FILLER_18_573 ();
 sg13g2_fill_1 FILLER_18_575 ();
 sg13g2_fill_2 FILLER_18_598 ();
 sg13g2_fill_1 FILLER_18_600 ();
 sg13g2_fill_1 FILLER_18_625 ();
 sg13g2_fill_1 FILLER_18_694 ();
 sg13g2_fill_1 FILLER_18_698 ();
 sg13g2_fill_1 FILLER_18_729 ();
 sg13g2_fill_2 FILLER_18_828 ();
 sg13g2_fill_2 FILLER_18_835 ();
 sg13g2_fill_2 FILLER_18_847 ();
 sg13g2_fill_1 FILLER_18_849 ();
 sg13g2_fill_2 FILLER_18_860 ();
 sg13g2_fill_2 FILLER_18_909 ();
 sg13g2_fill_1 FILLER_18_911 ();
 sg13g2_fill_2 FILLER_18_938 ();
 sg13g2_fill_1 FILLER_18_945 ();
 sg13g2_fill_2 FILLER_18_1049 ();
 sg13g2_fill_1 FILLER_18_1051 ();
 sg13g2_fill_2 FILLER_18_1066 ();
 sg13g2_fill_2 FILLER_18_1094 ();
 sg13g2_fill_1 FILLER_18_1096 ();
 sg13g2_fill_1 FILLER_18_1123 ();
 sg13g2_fill_2 FILLER_18_1172 ();
 sg13g2_fill_1 FILLER_18_1174 ();
 sg13g2_fill_1 FILLER_18_1196 ();
 sg13g2_fill_2 FILLER_18_1209 ();
 sg13g2_fill_1 FILLER_18_1211 ();
 sg13g2_fill_2 FILLER_18_1238 ();
 sg13g2_fill_1 FILLER_18_1284 ();
 sg13g2_fill_1 FILLER_18_1309 ();
 sg13g2_fill_2 FILLER_18_1344 ();
 sg13g2_fill_2 FILLER_18_1361 ();
 sg13g2_fill_1 FILLER_18_1363 ();
 sg13g2_decap_8 FILLER_18_1407 ();
 sg13g2_fill_2 FILLER_18_1414 ();
 sg13g2_fill_1 FILLER_18_1416 ();
 sg13g2_decap_8 FILLER_18_1430 ();
 sg13g2_fill_2 FILLER_18_1437 ();
 sg13g2_fill_1 FILLER_18_1439 ();
 sg13g2_fill_2 FILLER_18_1445 ();
 sg13g2_decap_4 FILLER_18_1455 ();
 sg13g2_decap_4 FILLER_18_1489 ();
 sg13g2_decap_4 FILLER_18_1524 ();
 sg13g2_fill_2 FILLER_18_1538 ();
 sg13g2_decap_4 FILLER_18_1553 ();
 sg13g2_fill_1 FILLER_18_1557 ();
 sg13g2_decap_4 FILLER_18_1574 ();
 sg13g2_fill_1 FILLER_18_1578 ();
 sg13g2_fill_2 FILLER_18_1592 ();
 sg13g2_fill_1 FILLER_18_1594 ();
 sg13g2_decap_8 FILLER_18_1615 ();
 sg13g2_decap_4 FILLER_18_1626 ();
 sg13g2_decap_4 FILLER_18_1638 ();
 sg13g2_fill_2 FILLER_18_1642 ();
 sg13g2_fill_2 FILLER_18_1751 ();
 sg13g2_fill_2 FILLER_18_1787 ();
 sg13g2_fill_1 FILLER_18_1789 ();
 sg13g2_fill_2 FILLER_18_1820 ();
 sg13g2_fill_2 FILLER_18_1837 ();
 sg13g2_fill_1 FILLER_18_1839 ();
 sg13g2_decap_8 FILLER_18_1900 ();
 sg13g2_fill_1 FILLER_18_1907 ();
 sg13g2_decap_4 FILLER_18_1934 ();
 sg13g2_fill_2 FILLER_18_1969 ();
 sg13g2_fill_1 FILLER_18_1971 ();
 sg13g2_fill_1 FILLER_18_2008 ();
 sg13g2_fill_2 FILLER_18_2035 ();
 sg13g2_fill_1 FILLER_18_2037 ();
 sg13g2_fill_2 FILLER_18_2051 ();
 sg13g2_fill_1 FILLER_18_2053 ();
 sg13g2_fill_2 FILLER_18_2107 ();
 sg13g2_fill_1 FILLER_18_2109 ();
 sg13g2_fill_1 FILLER_18_2180 ();
 sg13g2_fill_1 FILLER_18_2295 ();
 sg13g2_fill_1 FILLER_18_2345 ();
 sg13g2_fill_1 FILLER_18_2370 ();
 sg13g2_fill_2 FILLER_18_2461 ();
 sg13g2_fill_1 FILLER_18_2463 ();
 sg13g2_fill_2 FILLER_18_2491 ();
 sg13g2_fill_2 FILLER_18_2558 ();
 sg13g2_fill_1 FILLER_18_2569 ();
 sg13g2_fill_2 FILLER_18_2609 ();
 sg13g2_fill_1 FILLER_18_2647 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_376 ();
 sg13g2_fill_2 FILLER_19_418 ();
 sg13g2_fill_2 FILLER_19_486 ();
 sg13g2_fill_2 FILLER_19_587 ();
 sg13g2_fill_1 FILLER_19_627 ();
 sg13g2_fill_1 FILLER_19_650 ();
 sg13g2_fill_1 FILLER_19_703 ();
 sg13g2_fill_2 FILLER_19_718 ();
 sg13g2_fill_2 FILLER_19_725 ();
 sg13g2_fill_1 FILLER_19_727 ();
 sg13g2_fill_2 FILLER_19_741 ();
 sg13g2_fill_2 FILLER_19_752 ();
 sg13g2_fill_2 FILLER_19_819 ();
 sg13g2_fill_2 FILLER_19_839 ();
 sg13g2_fill_2 FILLER_19_850 ();
 sg13g2_fill_1 FILLER_19_865 ();
 sg13g2_fill_2 FILLER_19_880 ();
 sg13g2_fill_1 FILLER_19_882 ();
 sg13g2_fill_1 FILLER_19_927 ();
 sg13g2_fill_2 FILLER_19_947 ();
 sg13g2_fill_1 FILLER_19_954 ();
 sg13g2_fill_1 FILLER_19_968 ();
 sg13g2_fill_2 FILLER_19_979 ();
 sg13g2_fill_1 FILLER_19_1018 ();
 sg13g2_fill_2 FILLER_19_1031 ();
 sg13g2_fill_2 FILLER_19_1077 ();
 sg13g2_fill_2 FILLER_19_1096 ();
 sg13g2_fill_2 FILLER_19_1107 ();
 sg13g2_fill_2 FILLER_19_1126 ();
 sg13g2_fill_2 FILLER_19_1137 ();
 sg13g2_fill_2 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1149 ();
 sg13g2_fill_1 FILLER_19_1171 ();
 sg13g2_fill_1 FILLER_19_1180 ();
 sg13g2_fill_1 FILLER_19_1220 ();
 sg13g2_decap_4 FILLER_19_1261 ();
 sg13g2_decap_8 FILLER_19_1283 ();
 sg13g2_fill_2 FILLER_19_1290 ();
 sg13g2_fill_1 FILLER_19_1292 ();
 sg13g2_decap_4 FILLER_19_1311 ();
 sg13g2_fill_1 FILLER_19_1315 ();
 sg13g2_decap_8 FILLER_19_1358 ();
 sg13g2_fill_1 FILLER_19_1365 ();
 sg13g2_decap_8 FILLER_19_1370 ();
 sg13g2_decap_8 FILLER_19_1377 ();
 sg13g2_decap_8 FILLER_19_1389 ();
 sg13g2_fill_2 FILLER_19_1396 ();
 sg13g2_fill_2 FILLER_19_1436 ();
 sg13g2_fill_1 FILLER_19_1438 ();
 sg13g2_decap_4 FILLER_19_1486 ();
 sg13g2_fill_2 FILLER_19_1498 ();
 sg13g2_decap_4 FILLER_19_1510 ();
 sg13g2_fill_1 FILLER_19_1514 ();
 sg13g2_fill_1 FILLER_19_1520 ();
 sg13g2_fill_2 FILLER_19_1569 ();
 sg13g2_fill_1 FILLER_19_1571 ();
 sg13g2_fill_1 FILLER_19_1580 ();
 sg13g2_decap_4 FILLER_19_1585 ();
 sg13g2_fill_1 FILLER_19_1589 ();
 sg13g2_decap_4 FILLER_19_1594 ();
 sg13g2_fill_2 FILLER_19_1598 ();
 sg13g2_decap_4 FILLER_19_1634 ();
 sg13g2_fill_2 FILLER_19_1638 ();
 sg13g2_decap_4 FILLER_19_1653 ();
 sg13g2_fill_1 FILLER_19_1657 ();
 sg13g2_decap_8 FILLER_19_1677 ();
 sg13g2_fill_1 FILLER_19_1684 ();
 sg13g2_fill_2 FILLER_19_1772 ();
 sg13g2_fill_1 FILLER_19_1804 ();
 sg13g2_fill_2 FILLER_19_1873 ();
 sg13g2_fill_1 FILLER_19_1875 ();
 sg13g2_decap_4 FILLER_19_1901 ();
 sg13g2_fill_2 FILLER_19_1918 ();
 sg13g2_fill_1 FILLER_19_1920 ();
 sg13g2_fill_1 FILLER_19_1928 ();
 sg13g2_decap_4 FILLER_19_1938 ();
 sg13g2_fill_2 FILLER_19_1955 ();
 sg13g2_fill_2 FILLER_19_1995 ();
 sg13g2_fill_1 FILLER_19_1997 ();
 sg13g2_fill_1 FILLER_19_2029 ();
 sg13g2_fill_2 FILLER_19_2074 ();
 sg13g2_fill_1 FILLER_19_2076 ();
 sg13g2_decap_4 FILLER_19_2113 ();
 sg13g2_fill_1 FILLER_19_2117 ();
 sg13g2_fill_2 FILLER_19_2154 ();
 sg13g2_fill_1 FILLER_19_2156 ();
 sg13g2_fill_1 FILLER_19_2162 ();
 sg13g2_fill_2 FILLER_19_2203 ();
 sg13g2_fill_2 FILLER_19_2215 ();
 sg13g2_fill_1 FILLER_19_2217 ();
 sg13g2_fill_2 FILLER_19_2258 ();
 sg13g2_fill_1 FILLER_19_2260 ();
 sg13g2_fill_1 FILLER_19_2279 ();
 sg13g2_fill_2 FILLER_19_2291 ();
 sg13g2_fill_1 FILLER_19_2293 ();
 sg13g2_fill_1 FILLER_19_2324 ();
 sg13g2_fill_1 FILLER_19_2338 ();
 sg13g2_fill_2 FILLER_19_2368 ();
 sg13g2_fill_1 FILLER_19_2370 ();
 sg13g2_fill_2 FILLER_19_2414 ();
 sg13g2_fill_1 FILLER_19_2433 ();
 sg13g2_fill_2 FILLER_19_2444 ();
 sg13g2_fill_1 FILLER_19_2446 ();
 sg13g2_fill_2 FILLER_19_2477 ();
 sg13g2_fill_1 FILLER_19_2531 ();
 sg13g2_fill_1 FILLER_19_2548 ();
 sg13g2_fill_2 FILLER_19_2590 ();
 sg13g2_fill_1 FILLER_19_2592 ();
 sg13g2_fill_2 FILLER_19_2603 ();
 sg13g2_fill_1 FILLER_19_2637 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_452 ();
 sg13g2_fill_1 FILLER_20_489 ();
 sg13g2_fill_2 FILLER_20_527 ();
 sg13g2_fill_2 FILLER_20_538 ();
 sg13g2_fill_1 FILLER_20_540 ();
 sg13g2_fill_2 FILLER_20_630 ();
 sg13g2_fill_1 FILLER_20_632 ();
 sg13g2_fill_2 FILLER_20_724 ();
 sg13g2_fill_1 FILLER_20_726 ();
 sg13g2_fill_1 FILLER_20_739 ();
 sg13g2_fill_1 FILLER_20_794 ();
 sg13g2_fill_2 FILLER_20_805 ();
 sg13g2_fill_2 FILLER_20_811 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_2 FILLER_20_1039 ();
 sg13g2_fill_1 FILLER_20_1041 ();
 sg13g2_fill_2 FILLER_20_1052 ();
 sg13g2_fill_1 FILLER_20_1054 ();
 sg13g2_fill_2 FILLER_20_1117 ();
 sg13g2_fill_1 FILLER_20_1119 ();
 sg13g2_fill_2 FILLER_20_1156 ();
 sg13g2_fill_1 FILLER_20_1158 ();
 sg13g2_fill_1 FILLER_20_1198 ();
 sg13g2_fill_2 FILLER_20_1221 ();
 sg13g2_fill_1 FILLER_20_1256 ();
 sg13g2_decap_4 FILLER_20_1314 ();
 sg13g2_fill_1 FILLER_20_1326 ();
 sg13g2_decap_4 FILLER_20_1341 ();
 sg13g2_fill_1 FILLER_20_1345 ();
 sg13g2_decap_4 FILLER_20_1434 ();
 sg13g2_fill_1 FILLER_20_1438 ();
 sg13g2_fill_2 FILLER_20_1462 ();
 sg13g2_fill_1 FILLER_20_1490 ();
 sg13g2_fill_2 FILLER_20_1495 ();
 sg13g2_fill_1 FILLER_20_1497 ();
 sg13g2_decap_4 FILLER_20_1503 ();
 sg13g2_fill_1 FILLER_20_1507 ();
 sg13g2_decap_8 FILLER_20_1512 ();
 sg13g2_fill_1 FILLER_20_1519 ();
 sg13g2_decap_4 FILLER_20_1554 ();
 sg13g2_fill_1 FILLER_20_1570 ();
 sg13g2_fill_2 FILLER_20_1612 ();
 sg13g2_fill_1 FILLER_20_1614 ();
 sg13g2_fill_1 FILLER_20_1620 ();
 sg13g2_fill_2 FILLER_20_1642 ();
 sg13g2_fill_1 FILLER_20_1644 ();
 sg13g2_fill_2 FILLER_20_1649 ();
 sg13g2_decap_4 FILLER_20_1677 ();
 sg13g2_fill_2 FILLER_20_1681 ();
 sg13g2_fill_2 FILLER_20_1693 ();
 sg13g2_fill_2 FILLER_20_1718 ();
 sg13g2_fill_1 FILLER_20_1726 ();
 sg13g2_fill_1 FILLER_20_1785 ();
 sg13g2_fill_2 FILLER_20_1796 ();
 sg13g2_fill_1 FILLER_20_1798 ();
 sg13g2_decap_4 FILLER_20_1826 ();
 sg13g2_fill_2 FILLER_20_1830 ();
 sg13g2_fill_2 FILLER_20_1904 ();
 sg13g2_decap_4 FILLER_20_1932 ();
 sg13g2_fill_1 FILLER_20_1936 ();
 sg13g2_fill_2 FILLER_20_1982 ();
 sg13g2_fill_2 FILLER_20_2016 ();
 sg13g2_fill_2 FILLER_20_2023 ();
 sg13g2_fill_1 FILLER_20_2025 ();
 sg13g2_fill_2 FILLER_20_2035 ();
 sg13g2_fill_2 FILLER_20_2082 ();
 sg13g2_fill_1 FILLER_20_2084 ();
 sg13g2_decap_4 FILLER_20_2106 ();
 sg13g2_fill_1 FILLER_20_2132 ();
 sg13g2_fill_1 FILLER_20_2238 ();
 sg13g2_fill_2 FILLER_20_2348 ();
 sg13g2_fill_1 FILLER_20_2350 ();
 sg13g2_fill_1 FILLER_20_2388 ();
 sg13g2_fill_2 FILLER_20_2477 ();
 sg13g2_fill_1 FILLER_20_2479 ();
 sg13g2_fill_2 FILLER_20_2490 ();
 sg13g2_fill_1 FILLER_20_2492 ();
 sg13g2_fill_2 FILLER_20_2533 ();
 sg13g2_fill_1 FILLER_20_2535 ();
 sg13g2_fill_2 FILLER_20_2580 ();
 sg13g2_fill_2 FILLER_20_2636 ();
 sg13g2_fill_2 FILLER_20_2654 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_86 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_432 ();
 sg13g2_fill_2 FILLER_21_456 ();
 sg13g2_fill_2 FILLER_21_474 ();
 sg13g2_fill_1 FILLER_21_476 ();
 sg13g2_fill_1 FILLER_21_561 ();
 sg13g2_fill_1 FILLER_21_619 ();
 sg13g2_fill_2 FILLER_21_655 ();
 sg13g2_fill_1 FILLER_21_657 ();
 sg13g2_fill_2 FILLER_21_715 ();
 sg13g2_fill_1 FILLER_21_717 ();
 sg13g2_fill_2 FILLER_21_740 ();
 sg13g2_fill_2 FILLER_21_751 ();
 sg13g2_fill_2 FILLER_21_832 ();
 sg13g2_fill_1 FILLER_21_834 ();
 sg13g2_fill_1 FILLER_21_847 ();
 sg13g2_fill_2 FILLER_21_861 ();
 sg13g2_fill_2 FILLER_21_871 ();
 sg13g2_fill_1 FILLER_21_882 ();
 sg13g2_fill_2 FILLER_21_894 ();
 sg13g2_fill_2 FILLER_21_911 ();
 sg13g2_fill_1 FILLER_21_913 ();
 sg13g2_fill_2 FILLER_21_932 ();
 sg13g2_fill_1 FILLER_21_934 ();
 sg13g2_fill_2 FILLER_21_940 ();
 sg13g2_fill_1 FILLER_21_942 ();
 sg13g2_fill_1 FILLER_21_965 ();
 sg13g2_fill_2 FILLER_21_1053 ();
 sg13g2_fill_2 FILLER_21_1085 ();
 sg13g2_fill_1 FILLER_21_1087 ();
 sg13g2_fill_1 FILLER_21_1101 ();
 sg13g2_fill_2 FILLER_21_1119 ();
 sg13g2_fill_1 FILLER_21_1121 ();
 sg13g2_fill_1 FILLER_21_1132 ();
 sg13g2_fill_2 FILLER_21_1159 ();
 sg13g2_fill_1 FILLER_21_1176 ();
 sg13g2_fill_2 FILLER_21_1241 ();
 sg13g2_fill_1 FILLER_21_1243 ();
 sg13g2_fill_2 FILLER_21_1275 ();
 sg13g2_decap_4 FILLER_21_1291 ();
 sg13g2_fill_2 FILLER_21_1295 ();
 sg13g2_fill_2 FILLER_21_1329 ();
 sg13g2_fill_1 FILLER_21_1331 ();
 sg13g2_fill_1 FILLER_21_1337 ();
 sg13g2_decap_8 FILLER_21_1343 ();
 sg13g2_fill_2 FILLER_21_1350 ();
 sg13g2_fill_2 FILLER_21_1359 ();
 sg13g2_fill_2 FILLER_21_1366 ();
 sg13g2_decap_8 FILLER_21_1389 ();
 sg13g2_fill_2 FILLER_21_1396 ();
 sg13g2_fill_2 FILLER_21_1415 ();
 sg13g2_fill_2 FILLER_21_1533 ();
 sg13g2_fill_1 FILLER_21_1564 ();
 sg13g2_fill_2 FILLER_21_1622 ();
 sg13g2_fill_1 FILLER_21_1624 ();
 sg13g2_fill_2 FILLER_21_1660 ();
 sg13g2_fill_2 FILLER_21_1666 ();
 sg13g2_fill_2 FILLER_21_1724 ();
 sg13g2_fill_1 FILLER_21_1726 ();
 sg13g2_fill_2 FILLER_21_1745 ();
 sg13g2_fill_1 FILLER_21_1787 ();
 sg13g2_fill_1 FILLER_21_1843 ();
 sg13g2_fill_2 FILLER_21_1874 ();
 sg13g2_fill_1 FILLER_21_1876 ();
 sg13g2_fill_2 FILLER_21_1887 ();
 sg13g2_fill_1 FILLER_21_1889 ();
 sg13g2_fill_2 FILLER_21_1921 ();
 sg13g2_fill_1 FILLER_21_1923 ();
 sg13g2_fill_2 FILLER_21_1975 ();
 sg13g2_fill_1 FILLER_21_1977 ();
 sg13g2_fill_2 FILLER_21_2014 ();
 sg13g2_fill_1 FILLER_21_2016 ();
 sg13g2_fill_1 FILLER_21_2077 ();
 sg13g2_fill_2 FILLER_21_2132 ();
 sg13g2_fill_1 FILLER_21_2134 ();
 sg13g2_fill_2 FILLER_21_2143 ();
 sg13g2_fill_1 FILLER_21_2145 ();
 sg13g2_fill_2 FILLER_21_2162 ();
 sg13g2_fill_1 FILLER_21_2215 ();
 sg13g2_fill_2 FILLER_21_2277 ();
 sg13g2_fill_2 FILLER_21_2325 ();
 sg13g2_fill_1 FILLER_21_2327 ();
 sg13g2_fill_1 FILLER_21_2362 ();
 sg13g2_fill_2 FILLER_21_2409 ();
 sg13g2_fill_2 FILLER_21_2541 ();
 sg13g2_fill_1 FILLER_21_2543 ();
 sg13g2_fill_2 FILLER_21_2560 ();
 sg13g2_fill_1 FILLER_21_2587 ();
 sg13g2_fill_2 FILLER_21_2627 ();
 sg13g2_fill_2 FILLER_21_2645 ();
 sg13g2_fill_1 FILLER_21_2647 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_277 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_fill_2 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_411 ();
 sg13g2_fill_2 FILLER_22_487 ();
 sg13g2_fill_2 FILLER_22_542 ();
 sg13g2_fill_1 FILLER_22_544 ();
 sg13g2_fill_2 FILLER_22_777 ();
 sg13g2_fill_1 FILLER_22_779 ();
 sg13g2_fill_2 FILLER_22_839 ();
 sg13g2_fill_2 FILLER_22_895 ();
 sg13g2_fill_1 FILLER_22_897 ();
 sg13g2_fill_2 FILLER_22_924 ();
 sg13g2_fill_1 FILLER_22_926 ();
 sg13g2_fill_2 FILLER_22_990 ();
 sg13g2_fill_1 FILLER_22_992 ();
 sg13g2_fill_2 FILLER_22_1017 ();
 sg13g2_fill_1 FILLER_22_1039 ();
 sg13g2_fill_1 FILLER_22_1057 ();
 sg13g2_fill_2 FILLER_22_1102 ();
 sg13g2_fill_1 FILLER_22_1104 ();
 sg13g2_fill_2 FILLER_22_1131 ();
 sg13g2_fill_1 FILLER_22_1133 ();
 sg13g2_fill_1 FILLER_22_1160 ();
 sg13g2_fill_2 FILLER_22_1166 ();
 sg13g2_fill_1 FILLER_22_1208 ();
 sg13g2_fill_1 FILLER_22_1218 ();
 sg13g2_fill_1 FILLER_22_1255 ();
 sg13g2_decap_8 FILLER_22_1298 ();
 sg13g2_fill_1 FILLER_22_1305 ();
 sg13g2_fill_2 FILLER_22_1327 ();
 sg13g2_fill_1 FILLER_22_1376 ();
 sg13g2_fill_2 FILLER_22_1416 ();
 sg13g2_fill_1 FILLER_22_1418 ();
 sg13g2_fill_2 FILLER_22_1428 ();
 sg13g2_fill_2 FILLER_22_1486 ();
 sg13g2_fill_1 FILLER_22_1558 ();
 sg13g2_fill_2 FILLER_22_1577 ();
 sg13g2_fill_1 FILLER_22_1579 ();
 sg13g2_fill_2 FILLER_22_1593 ();
 sg13g2_fill_1 FILLER_22_1606 ();
 sg13g2_fill_2 FILLER_22_1642 ();
 sg13g2_fill_1 FILLER_22_1644 ();
 sg13g2_fill_1 FILLER_22_1691 ();
 sg13g2_fill_1 FILLER_22_1738 ();
 sg13g2_fill_2 FILLER_22_1770 ();
 sg13g2_fill_2 FILLER_22_1861 ();
 sg13g2_fill_1 FILLER_22_1863 ();
 sg13g2_fill_2 FILLER_22_1874 ();
 sg13g2_fill_1 FILLER_22_1876 ();
 sg13g2_fill_1 FILLER_22_1887 ();
 sg13g2_fill_2 FILLER_22_1914 ();
 sg13g2_fill_2 FILLER_22_1920 ();
 sg13g2_fill_1 FILLER_22_1922 ();
 sg13g2_fill_2 FILLER_22_1942 ();
 sg13g2_fill_2 FILLER_22_1958 ();
 sg13g2_fill_1 FILLER_22_2005 ();
 sg13g2_fill_1 FILLER_22_2143 ();
 sg13g2_fill_2 FILLER_22_2152 ();
 sg13g2_fill_1 FILLER_22_2180 ();
 sg13g2_fill_2 FILLER_22_2210 ();
 sg13g2_fill_2 FILLER_22_2248 ();
 sg13g2_fill_1 FILLER_22_2250 ();
 sg13g2_decap_4 FILLER_22_2265 ();
 sg13g2_fill_1 FILLER_22_2349 ();
 sg13g2_fill_1 FILLER_22_2399 ();
 sg13g2_fill_2 FILLER_22_2433 ();
 sg13g2_fill_2 FILLER_22_2492 ();
 sg13g2_fill_1 FILLER_22_2494 ();
 sg13g2_fill_2 FILLER_22_2546 ();
 sg13g2_fill_1 FILLER_22_2548 ();
 sg13g2_fill_1 FILLER_22_2590 ();
 sg13g2_fill_1 FILLER_22_2626 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_405 ();
 sg13g2_fill_1 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_534 ();
 sg13g2_fill_1 FILLER_23_562 ();
 sg13g2_fill_1 FILLER_23_573 ();
 sg13g2_fill_2 FILLER_23_583 ();
 sg13g2_fill_2 FILLER_23_595 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_fill_1 FILLER_23_612 ();
 sg13g2_fill_2 FILLER_23_673 ();
 sg13g2_fill_2 FILLER_23_683 ();
 sg13g2_fill_1 FILLER_23_711 ();
 sg13g2_fill_2 FILLER_23_737 ();
 sg13g2_fill_2 FILLER_23_744 ();
 sg13g2_fill_1 FILLER_23_746 ();
 sg13g2_fill_1 FILLER_23_810 ();
 sg13g2_fill_2 FILLER_23_865 ();
 sg13g2_fill_2 FILLER_23_879 ();
 sg13g2_fill_1 FILLER_23_881 ();
 sg13g2_fill_2 FILLER_23_913 ();
 sg13g2_fill_1 FILLER_23_915 ();
 sg13g2_fill_2 FILLER_23_948 ();
 sg13g2_fill_1 FILLER_23_950 ();
 sg13g2_fill_1 FILLER_23_964 ();
 sg13g2_fill_1 FILLER_23_1002 ();
 sg13g2_fill_2 FILLER_23_1081 ();
 sg13g2_fill_1 FILLER_23_1083 ();
 sg13g2_fill_2 FILLER_23_1129 ();
 sg13g2_fill_1 FILLER_23_1136 ();
 sg13g2_fill_2 FILLER_23_1141 ();
 sg13g2_fill_1 FILLER_23_1143 ();
 sg13g2_fill_2 FILLER_23_1174 ();
 sg13g2_fill_1 FILLER_23_1176 ();
 sg13g2_fill_1 FILLER_23_1196 ();
 sg13g2_fill_2 FILLER_23_1208 ();
 sg13g2_fill_1 FILLER_23_1210 ();
 sg13g2_fill_2 FILLER_23_1306 ();
 sg13g2_fill_1 FILLER_23_1308 ();
 sg13g2_fill_2 FILLER_23_1372 ();
 sg13g2_fill_1 FILLER_23_1374 ();
 sg13g2_decap_8 FILLER_23_1391 ();
 sg13g2_fill_1 FILLER_23_1398 ();
 sg13g2_fill_2 FILLER_23_1407 ();
 sg13g2_fill_1 FILLER_23_1409 ();
 sg13g2_fill_2 FILLER_23_1462 ();
 sg13g2_fill_2 FILLER_23_1512 ();
 sg13g2_fill_1 FILLER_23_1514 ();
 sg13g2_fill_2 FILLER_23_1532 ();
 sg13g2_fill_1 FILLER_23_1542 ();
 sg13g2_fill_1 FILLER_23_1552 ();
 sg13g2_fill_1 FILLER_23_1567 ();
 sg13g2_decap_8 FILLER_23_1576 ();
 sg13g2_decap_4 FILLER_23_1605 ();
 sg13g2_fill_1 FILLER_23_1634 ();
 sg13g2_decap_4 FILLER_23_1654 ();
 sg13g2_fill_1 FILLER_23_1658 ();
 sg13g2_fill_2 FILLER_23_1686 ();
 sg13g2_fill_2 FILLER_23_1791 ();
 sg13g2_fill_2 FILLER_23_1840 ();
 sg13g2_decap_8 FILLER_23_1915 ();
 sg13g2_fill_2 FILLER_23_1977 ();
 sg13g2_fill_1 FILLER_23_1979 ();
 sg13g2_fill_1 FILLER_23_2023 ();
 sg13g2_fill_1 FILLER_23_2067 ();
 sg13g2_fill_2 FILLER_23_2112 ();
 sg13g2_fill_2 FILLER_23_2119 ();
 sg13g2_fill_2 FILLER_23_2231 ();
 sg13g2_fill_1 FILLER_23_2233 ();
 sg13g2_decap_8 FILLER_23_2360 ();
 sg13g2_fill_1 FILLER_23_2393 ();
 sg13g2_fill_2 FILLER_23_2445 ();
 sg13g2_fill_2 FILLER_23_2536 ();
 sg13g2_fill_2 FILLER_23_2559 ();
 sg13g2_fill_1 FILLER_23_2643 ();
 sg13g2_fill_2 FILLER_23_2671 ();
 sg13g2_fill_1 FILLER_23_2673 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_433 ();
 sg13g2_fill_2 FILLER_24_462 ();
 sg13g2_fill_2 FILLER_24_530 ();
 sg13g2_fill_1 FILLER_24_532 ();
 sg13g2_fill_1 FILLER_24_543 ();
 sg13g2_fill_2 FILLER_24_595 ();
 sg13g2_fill_2 FILLER_24_612 ();
 sg13g2_fill_1 FILLER_24_614 ();
 sg13g2_fill_2 FILLER_24_655 ();
 sg13g2_fill_1 FILLER_24_657 ();
 sg13g2_fill_2 FILLER_24_694 ();
 sg13g2_fill_2 FILLER_24_783 ();
 sg13g2_fill_1 FILLER_24_785 ();
 sg13g2_fill_1 FILLER_24_790 ();
 sg13g2_fill_2 FILLER_24_802 ();
 sg13g2_fill_1 FILLER_24_825 ();
 sg13g2_fill_1 FILLER_24_856 ();
 sg13g2_fill_1 FILLER_24_885 ();
 sg13g2_fill_2 FILLER_24_892 ();
 sg13g2_fill_2 FILLER_24_907 ();
 sg13g2_fill_2 FILLER_24_917 ();
 sg13g2_fill_1 FILLER_24_919 ();
 sg13g2_fill_2 FILLER_24_938 ();
 sg13g2_fill_1 FILLER_24_940 ();
 sg13g2_fill_2 FILLER_24_946 ();
 sg13g2_fill_1 FILLER_24_948 ();
 sg13g2_fill_2 FILLER_24_960 ();
 sg13g2_fill_1 FILLER_24_1001 ();
 sg13g2_fill_1 FILLER_24_1037 ();
 sg13g2_fill_1 FILLER_24_1069 ();
 sg13g2_fill_1 FILLER_24_1096 ();
 sg13g2_fill_2 FILLER_24_1163 ();
 sg13g2_fill_1 FILLER_24_1165 ();
 sg13g2_fill_2 FILLER_24_1192 ();
 sg13g2_fill_1 FILLER_24_1251 ();
 sg13g2_fill_1 FILLER_24_1257 ();
 sg13g2_fill_1 FILLER_24_1275 ();
 sg13g2_fill_2 FILLER_24_1351 ();
 sg13g2_decap_4 FILLER_24_1371 ();
 sg13g2_fill_1 FILLER_24_1375 ();
 sg13g2_decap_8 FILLER_24_1393 ();
 sg13g2_fill_1 FILLER_24_1400 ();
 sg13g2_decap_8 FILLER_24_1405 ();
 sg13g2_decap_4 FILLER_24_1412 ();
 sg13g2_fill_1 FILLER_24_1416 ();
 sg13g2_fill_2 FILLER_24_1433 ();
 sg13g2_fill_1 FILLER_24_1435 ();
 sg13g2_fill_2 FILLER_24_1512 ();
 sg13g2_fill_2 FILLER_24_1533 ();
 sg13g2_fill_2 FILLER_24_1551 ();
 sg13g2_fill_1 FILLER_24_1561 ();
 sg13g2_decap_4 FILLER_24_1587 ();
 sg13g2_fill_1 FILLER_24_1591 ();
 sg13g2_fill_2 FILLER_24_1609 ();
 sg13g2_fill_1 FILLER_24_1611 ();
 sg13g2_fill_2 FILLER_24_1664 ();
 sg13g2_fill_1 FILLER_24_1666 ();
 sg13g2_fill_2 FILLER_24_1693 ();
 sg13g2_fill_2 FILLER_24_1724 ();
 sg13g2_fill_1 FILLER_24_1801 ();
 sg13g2_fill_1 FILLER_24_1810 ();
 sg13g2_fill_2 FILLER_24_1821 ();
 sg13g2_fill_2 FILLER_24_1836 ();
 sg13g2_fill_1 FILLER_24_1860 ();
 sg13g2_fill_2 FILLER_24_1884 ();
 sg13g2_fill_1 FILLER_24_1910 ();
 sg13g2_fill_2 FILLER_24_1945 ();
 sg13g2_fill_2 FILLER_24_2040 ();
 sg13g2_fill_1 FILLER_24_2042 ();
 sg13g2_fill_1 FILLER_24_2079 ();
 sg13g2_fill_1 FILLER_24_2090 ();
 sg13g2_fill_1 FILLER_24_2114 ();
 sg13g2_fill_2 FILLER_24_2157 ();
 sg13g2_fill_2 FILLER_24_2191 ();
 sg13g2_fill_1 FILLER_24_2193 ();
 sg13g2_fill_2 FILLER_24_2284 ();
 sg13g2_fill_2 FILLER_24_2322 ();
 sg13g2_fill_1 FILLER_24_2384 ();
 sg13g2_fill_2 FILLER_24_2447 ();
 sg13g2_fill_1 FILLER_24_2449 ();
 sg13g2_fill_2 FILLER_24_2485 ();
 sg13g2_fill_1 FILLER_24_2545 ();
 sg13g2_fill_1 FILLER_24_2673 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_decap_4 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_44 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_fill_2 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_25_421 ();
 sg13g2_fill_1 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_453 ();
 sg13g2_fill_2 FILLER_25_514 ();
 sg13g2_fill_1 FILLER_25_516 ();
 sg13g2_fill_2 FILLER_25_566 ();
 sg13g2_fill_1 FILLER_25_568 ();
 sg13g2_fill_2 FILLER_25_676 ();
 sg13g2_fill_2 FILLER_25_741 ();
 sg13g2_fill_1 FILLER_25_743 ();
 sg13g2_fill_2 FILLER_25_753 ();
 sg13g2_fill_1 FILLER_25_755 ();
 sg13g2_fill_2 FILLER_25_760 ();
 sg13g2_fill_1 FILLER_25_762 ();
 sg13g2_fill_2 FILLER_25_776 ();
 sg13g2_fill_2 FILLER_25_782 ();
 sg13g2_fill_1 FILLER_25_784 ();
 sg13g2_fill_1 FILLER_25_847 ();
 sg13g2_fill_2 FILLER_25_874 ();
 sg13g2_fill_1 FILLER_25_876 ();
 sg13g2_fill_2 FILLER_25_889 ();
 sg13g2_fill_2 FILLER_25_972 ();
 sg13g2_fill_1 FILLER_25_1003 ();
 sg13g2_fill_2 FILLER_25_1021 ();
 sg13g2_fill_1 FILLER_25_1023 ();
 sg13g2_fill_2 FILLER_25_1033 ();
 sg13g2_fill_2 FILLER_25_1104 ();
 sg13g2_fill_2 FILLER_25_1137 ();
 sg13g2_fill_2 FILLER_25_1175 ();
 sg13g2_fill_1 FILLER_25_1177 ();
 sg13g2_fill_2 FILLER_25_1183 ();
 sg13g2_fill_2 FILLER_25_1206 ();
 sg13g2_fill_1 FILLER_25_1222 ();
 sg13g2_fill_2 FILLER_25_1240 ();
 sg13g2_fill_1 FILLER_25_1326 ();
 sg13g2_decap_4 FILLER_25_1369 ();
 sg13g2_fill_1 FILLER_25_1416 ();
 sg13g2_fill_2 FILLER_25_1428 ();
 sg13g2_fill_1 FILLER_25_1430 ();
 sg13g2_fill_2 FILLER_25_1460 ();
 sg13g2_fill_1 FILLER_25_1470 ();
 sg13g2_fill_2 FILLER_25_1502 ();
 sg13g2_decap_8 FILLER_25_1524 ();
 sg13g2_fill_1 FILLER_25_1556 ();
 sg13g2_fill_1 FILLER_25_1611 ();
 sg13g2_fill_2 FILLER_25_1637 ();
 sg13g2_fill_1 FILLER_25_1639 ();
 sg13g2_fill_1 FILLER_25_1654 ();
 sg13g2_fill_2 FILLER_25_1673 ();
 sg13g2_fill_1 FILLER_25_1708 ();
 sg13g2_fill_1 FILLER_25_1775 ();
 sg13g2_fill_1 FILLER_25_1812 ();
 sg13g2_fill_1 FILLER_25_1843 ();
 sg13g2_fill_1 FILLER_25_1880 ();
 sg13g2_fill_1 FILLER_25_1921 ();
 sg13g2_fill_2 FILLER_25_2011 ();
 sg13g2_fill_2 FILLER_25_2031 ();
 sg13g2_fill_1 FILLER_25_2033 ();
 sg13g2_decap_8 FILLER_25_2063 ();
 sg13g2_fill_2 FILLER_25_2125 ();
 sg13g2_fill_1 FILLER_25_2127 ();
 sg13g2_fill_2 FILLER_25_2187 ();
 sg13g2_fill_1 FILLER_25_2219 ();
 sg13g2_fill_2 FILLER_25_2230 ();
 sg13g2_decap_4 FILLER_25_2284 ();
 sg13g2_fill_2 FILLER_25_2320 ();
 sg13g2_fill_1 FILLER_25_2327 ();
 sg13g2_fill_1 FILLER_25_2335 ();
 sg13g2_decap_4 FILLER_25_2345 ();
 sg13g2_fill_1 FILLER_25_2349 ();
 sg13g2_decap_4 FILLER_25_2389 ();
 sg13g2_fill_1 FILLER_25_2393 ();
 sg13g2_fill_1 FILLER_25_2408 ();
 sg13g2_fill_2 FILLER_25_2419 ();
 sg13g2_fill_2 FILLER_25_2467 ();
 sg13g2_fill_2 FILLER_25_2505 ();
 sg13g2_fill_1 FILLER_25_2507 ();
 sg13g2_fill_2 FILLER_25_2530 ();
 sg13g2_fill_2 FILLER_25_2577 ();
 sg13g2_fill_1 FILLER_25_2579 ();
 sg13g2_fill_1 FILLER_25_2590 ();
 sg13g2_fill_2 FILLER_25_2606 ();
 sg13g2_fill_1 FILLER_25_2627 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_418 ();
 sg13g2_fill_2 FILLER_26_478 ();
 sg13g2_fill_1 FILLER_26_512 ();
 sg13g2_fill_1 FILLER_26_539 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_fill_2 FILLER_26_590 ();
 sg13g2_fill_1 FILLER_26_592 ();
 sg13g2_fill_2 FILLER_26_598 ();
 sg13g2_fill_1 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_609 ();
 sg13g2_fill_2 FILLER_26_628 ();
 sg13g2_fill_2 FILLER_26_651 ();
 sg13g2_fill_1 FILLER_26_653 ();
 sg13g2_fill_2 FILLER_26_814 ();
 sg13g2_fill_1 FILLER_26_816 ();
 sg13g2_fill_2 FILLER_26_830 ();
 sg13g2_fill_1 FILLER_26_832 ();
 sg13g2_fill_2 FILLER_26_842 ();
 sg13g2_fill_1 FILLER_26_863 ();
 sg13g2_fill_2 FILLER_26_904 ();
 sg13g2_decap_4 FILLER_26_1001 ();
 sg13g2_fill_1 FILLER_26_1005 ();
 sg13g2_fill_2 FILLER_26_1015 ();
 sg13g2_fill_1 FILLER_26_1017 ();
 sg13g2_fill_2 FILLER_26_1024 ();
 sg13g2_fill_1 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1053 ();
 sg13g2_fill_2 FILLER_26_1064 ();
 sg13g2_fill_1 FILLER_26_1093 ();
 sg13g2_fill_2 FILLER_26_1098 ();
 sg13g2_fill_2 FILLER_26_1108 ();
 sg13g2_fill_2 FILLER_26_1146 ();
 sg13g2_fill_2 FILLER_26_1162 ();
 sg13g2_fill_1 FILLER_26_1164 ();
 sg13g2_fill_2 FILLER_26_1245 ();
 sg13g2_fill_1 FILLER_26_1293 ();
 sg13g2_fill_1 FILLER_26_1326 ();
 sg13g2_fill_2 FILLER_26_1340 ();
 sg13g2_fill_1 FILLER_26_1342 ();
 sg13g2_fill_1 FILLER_26_1358 ();
 sg13g2_fill_2 FILLER_26_1414 ();
 sg13g2_fill_2 FILLER_26_1455 ();
 sg13g2_decap_8 FILLER_26_1465 ();
 sg13g2_fill_2 FILLER_26_1472 ();
 sg13g2_fill_1 FILLER_26_1474 ();
 sg13g2_fill_2 FILLER_26_1480 ();
 sg13g2_fill_2 FILLER_26_1516 ();
 sg13g2_fill_1 FILLER_26_1518 ();
 sg13g2_fill_1 FILLER_26_1542 ();
 sg13g2_decap_4 FILLER_26_1563 ();
 sg13g2_fill_2 FILLER_26_1582 ();
 sg13g2_fill_2 FILLER_26_1603 ();
 sg13g2_fill_1 FILLER_26_1605 ();
 sg13g2_fill_2 FILLER_26_1637 ();
 sg13g2_fill_1 FILLER_26_1746 ();
 sg13g2_fill_1 FILLER_26_1776 ();
 sg13g2_fill_2 FILLER_26_1798 ();
 sg13g2_fill_1 FILLER_26_1804 ();
 sg13g2_decap_4 FILLER_26_1815 ();
 sg13g2_fill_1 FILLER_26_1824 ();
 sg13g2_fill_1 FILLER_26_1929 ();
 sg13g2_fill_1 FILLER_26_1971 ();
 sg13g2_fill_2 FILLER_26_1982 ();
 sg13g2_fill_1 FILLER_26_1984 ();
 sg13g2_fill_1 FILLER_26_2021 ();
 sg13g2_fill_2 FILLER_26_2156 ();
 sg13g2_fill_1 FILLER_26_2227 ();
 sg13g2_fill_1 FILLER_26_2251 ();
 sg13g2_decap_4 FILLER_26_2292 ();
 sg13g2_fill_1 FILLER_26_2322 ();
 sg13g2_fill_1 FILLER_26_2368 ();
 sg13g2_fill_2 FILLER_26_2395 ();
 sg13g2_fill_1 FILLER_26_2397 ();
 sg13g2_fill_2 FILLER_26_2424 ();
 sg13g2_fill_1 FILLER_26_2426 ();
 sg13g2_fill_2 FILLER_26_2446 ();
 sg13g2_fill_2 FILLER_26_2467 ();
 sg13g2_fill_1 FILLER_26_2469 ();
 sg13g2_fill_2 FILLER_26_2484 ();
 sg13g2_fill_1 FILLER_26_2568 ();
 sg13g2_fill_2 FILLER_26_2612 ();
 sg13g2_decap_4 FILLER_26_2644 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_fill_1 FILLER_27_397 ();
 sg13g2_fill_2 FILLER_27_440 ();
 sg13g2_fill_1 FILLER_27_442 ();
 sg13g2_fill_1 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_597 ();
 sg13g2_fill_1 FILLER_27_599 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_640 ();
 sg13g2_fill_2 FILLER_27_683 ();
 sg13g2_fill_2 FILLER_27_690 ();
 sg13g2_fill_1 FILLER_27_692 ();
 sg13g2_fill_1 FILLER_27_701 ();
 sg13g2_fill_2 FILLER_27_715 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_fill_1 FILLER_27_727 ();
 sg13g2_fill_1 FILLER_27_733 ();
 sg13g2_fill_2 FILLER_27_742 ();
 sg13g2_fill_1 FILLER_27_744 ();
 sg13g2_fill_2 FILLER_27_754 ();
 sg13g2_decap_4 FILLER_27_771 ();
 sg13g2_fill_2 FILLER_27_810 ();
 sg13g2_fill_2 FILLER_27_874 ();
 sg13g2_fill_1 FILLER_27_876 ();
 sg13g2_fill_2 FILLER_27_883 ();
 sg13g2_fill_2 FILLER_27_920 ();
 sg13g2_fill_1 FILLER_27_922 ();
 sg13g2_fill_2 FILLER_27_979 ();
 sg13g2_fill_1 FILLER_27_981 ();
 sg13g2_fill_2 FILLER_27_990 ();
 sg13g2_fill_1 FILLER_27_992 ();
 sg13g2_fill_2 FILLER_27_998 ();
 sg13g2_fill_2 FILLER_27_1039 ();
 sg13g2_fill_1 FILLER_27_1059 ();
 sg13g2_fill_2 FILLER_27_1070 ();
 sg13g2_fill_1 FILLER_27_1072 ();
 sg13g2_fill_2 FILLER_27_1129 ();
 sg13g2_fill_1 FILLER_27_1176 ();
 sg13g2_fill_1 FILLER_27_1190 ();
 sg13g2_fill_2 FILLER_27_1263 ();
 sg13g2_fill_2 FILLER_27_1279 ();
 sg13g2_fill_1 FILLER_27_1326 ();
 sg13g2_decap_4 FILLER_27_1418 ();
 sg13g2_fill_1 FILLER_27_1422 ();
 sg13g2_fill_2 FILLER_27_1444 ();
 sg13g2_fill_1 FILLER_27_1446 ();
 sg13g2_fill_2 FILLER_27_1451 ();
 sg13g2_fill_2 FILLER_27_1461 ();
 sg13g2_fill_2 FILLER_27_1471 ();
 sg13g2_fill_1 FILLER_27_1473 ();
 sg13g2_fill_1 FILLER_27_1500 ();
 sg13g2_fill_2 FILLER_27_1514 ();
 sg13g2_fill_1 FILLER_27_1516 ();
 sg13g2_fill_2 FILLER_27_1525 ();
 sg13g2_fill_1 FILLER_27_1527 ();
 sg13g2_fill_1 FILLER_27_1536 ();
 sg13g2_fill_2 FILLER_27_1548 ();
 sg13g2_fill_1 FILLER_27_1563 ();
 sg13g2_fill_2 FILLER_27_1594 ();
 sg13g2_fill_1 FILLER_27_1596 ();
 sg13g2_fill_1 FILLER_27_1621 ();
 sg13g2_fill_2 FILLER_27_1630 ();
 sg13g2_fill_1 FILLER_27_1632 ();
 sg13g2_decap_8 FILLER_27_1641 ();
 sg13g2_fill_2 FILLER_27_1648 ();
 sg13g2_fill_1 FILLER_27_1654 ();
 sg13g2_decap_4 FILLER_27_1690 ();
 sg13g2_fill_2 FILLER_27_1694 ();
 sg13g2_fill_1 FILLER_27_1710 ();
 sg13g2_fill_2 FILLER_27_1755 ();
 sg13g2_fill_1 FILLER_27_1757 ();
 sg13g2_fill_1 FILLER_27_1788 ();
 sg13g2_fill_1 FILLER_27_1847 ();
 sg13g2_fill_2 FILLER_27_1894 ();
 sg13g2_fill_2 FILLER_27_1958 ();
 sg13g2_fill_1 FILLER_27_2056 ();
 sg13g2_fill_1 FILLER_27_2132 ();
 sg13g2_fill_1 FILLER_27_2146 ();
 sg13g2_fill_2 FILLER_27_2178 ();
 sg13g2_fill_2 FILLER_27_2262 ();
 sg13g2_fill_2 FILLER_27_2364 ();
 sg13g2_decap_8 FILLER_27_2374 ();
 sg13g2_fill_2 FILLER_27_2381 ();
 sg13g2_decap_4 FILLER_27_2388 ();
 sg13g2_fill_1 FILLER_27_2392 ();
 sg13g2_fill_1 FILLER_27_2406 ();
 sg13g2_fill_1 FILLER_27_2459 ();
 sg13g2_fill_1 FILLER_27_2468 ();
 sg13g2_fill_2 FILLER_27_2490 ();
 sg13g2_fill_1 FILLER_27_2492 ();
 sg13g2_decap_4 FILLER_27_2525 ();
 sg13g2_fill_1 FILLER_27_2542 ();
 sg13g2_fill_1 FILLER_27_2590 ();
 sg13g2_decap_4 FILLER_27_2651 ();
 sg13g2_fill_2 FILLER_27_2655 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_17 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_57 ();
 sg13g2_decap_4 FILLER_28_73 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_fill_2 FILLER_28_481 ();
 sg13g2_fill_1 FILLER_28_493 ();
 sg13g2_fill_2 FILLER_28_505 ();
 sg13g2_fill_2 FILLER_28_521 ();
 sg13g2_fill_1 FILLER_28_523 ();
 sg13g2_fill_2 FILLER_28_539 ();
 sg13g2_fill_2 FILLER_28_572 ();
 sg13g2_fill_1 FILLER_28_574 ();
 sg13g2_fill_2 FILLER_28_592 ();
 sg13g2_fill_2 FILLER_28_599 ();
 sg13g2_decap_4 FILLER_28_761 ();
 sg13g2_fill_1 FILLER_28_765 ();
 sg13g2_fill_2 FILLER_28_784 ();
 sg13g2_fill_1 FILLER_28_786 ();
 sg13g2_fill_2 FILLER_28_847 ();
 sg13g2_fill_2 FILLER_28_864 ();
 sg13g2_fill_1 FILLER_28_866 ();
 sg13g2_fill_2 FILLER_28_877 ();
 sg13g2_fill_2 FILLER_28_885 ();
 sg13g2_fill_1 FILLER_28_887 ();
 sg13g2_fill_1 FILLER_28_912 ();
 sg13g2_fill_2 FILLER_28_948 ();
 sg13g2_fill_1 FILLER_28_971 ();
 sg13g2_fill_2 FILLER_28_1003 ();
 sg13g2_fill_1 FILLER_28_1005 ();
 sg13g2_fill_2 FILLER_28_1016 ();
 sg13g2_fill_1 FILLER_28_1018 ();
 sg13g2_fill_1 FILLER_28_1029 ();
 sg13g2_fill_1 FILLER_28_1067 ();
 sg13g2_fill_2 FILLER_28_1094 ();
 sg13g2_fill_2 FILLER_28_1126 ();
 sg13g2_fill_2 FILLER_28_1142 ();
 sg13g2_fill_2 FILLER_28_1210 ();
 sg13g2_fill_2 FILLER_28_1242 ();
 sg13g2_fill_2 FILLER_28_1310 ();
 sg13g2_fill_1 FILLER_28_1312 ();
 sg13g2_fill_1 FILLER_28_1318 ();
 sg13g2_fill_2 FILLER_28_1329 ();
 sg13g2_decap_8 FILLER_28_1352 ();
 sg13g2_decap_8 FILLER_28_1359 ();
 sg13g2_fill_1 FILLER_28_1366 ();
 sg13g2_fill_2 FILLER_28_1410 ();
 sg13g2_decap_4 FILLER_28_1424 ();
 sg13g2_fill_1 FILLER_28_1428 ();
 sg13g2_fill_2 FILLER_28_1444 ();
 sg13g2_fill_1 FILLER_28_1446 ();
 sg13g2_fill_1 FILLER_28_1452 ();
 sg13g2_fill_1 FILLER_28_1459 ();
 sg13g2_fill_2 FILLER_28_1482 ();
 sg13g2_fill_1 FILLER_28_1484 ();
 sg13g2_fill_1 FILLER_28_1516 ();
 sg13g2_fill_2 FILLER_28_1523 ();
 sg13g2_decap_4 FILLER_28_1535 ();
 sg13g2_decap_8 FILLER_28_1545 ();
 sg13g2_fill_1 FILLER_28_1552 ();
 sg13g2_decap_8 FILLER_28_1561 ();
 sg13g2_fill_1 FILLER_28_1568 ();
 sg13g2_fill_1 FILLER_28_1574 ();
 sg13g2_fill_2 FILLER_28_1587 ();
 sg13g2_fill_1 FILLER_28_1589 ();
 sg13g2_fill_1 FILLER_28_1596 ();
 sg13g2_fill_1 FILLER_28_1601 ();
 sg13g2_decap_8 FILLER_28_1613 ();
 sg13g2_decap_8 FILLER_28_1648 ();
 sg13g2_fill_2 FILLER_28_1685 ();
 sg13g2_fill_2 FILLER_28_1691 ();
 sg13g2_fill_1 FILLER_28_1708 ();
 sg13g2_fill_1 FILLER_28_1739 ();
 sg13g2_fill_2 FILLER_28_1744 ();
 sg13g2_fill_2 FILLER_28_1767 ();
 sg13g2_fill_1 FILLER_28_1782 ();
 sg13g2_fill_2 FILLER_28_1806 ();
 sg13g2_fill_1 FILLER_28_1808 ();
 sg13g2_fill_1 FILLER_28_1821 ();
 sg13g2_fill_2 FILLER_28_1858 ();
 sg13g2_fill_2 FILLER_28_1866 ();
 sg13g2_fill_1 FILLER_28_1895 ();
 sg13g2_fill_2 FILLER_28_1966 ();
 sg13g2_fill_1 FILLER_28_1968 ();
 sg13g2_fill_2 FILLER_28_1983 ();
 sg13g2_fill_1 FILLER_28_2063 ();
 sg13g2_fill_2 FILLER_28_2115 ();
 sg13g2_decap_4 FILLER_28_2161 ();
 sg13g2_fill_1 FILLER_28_2165 ();
 sg13g2_fill_1 FILLER_28_2219 ();
 sg13g2_fill_2 FILLER_28_2230 ();
 sg13g2_fill_1 FILLER_28_2237 ();
 sg13g2_fill_1 FILLER_28_2295 ();
 sg13g2_fill_2 FILLER_28_2322 ();
 sg13g2_fill_1 FILLER_28_2324 ();
 sg13g2_fill_2 FILLER_28_2383 ();
 sg13g2_fill_1 FILLER_28_2441 ();
 sg13g2_fill_2 FILLER_28_2468 ();
 sg13g2_fill_1 FILLER_28_2470 ();
 sg13g2_fill_2 FILLER_28_2511 ();
 sg13g2_fill_1 FILLER_28_2563 ();
 sg13g2_fill_2 FILLER_28_2573 ();
 sg13g2_fill_1 FILLER_28_2575 ();
 sg13g2_fill_1 FILLER_28_2612 ();
 sg13g2_fill_2 FILLER_28_2645 ();
 sg13g2_fill_1 FILLER_28_2673 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_29 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_287 ();
 sg13g2_fill_1 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_372 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_fill_1 FILLER_29_414 ();
 sg13g2_fill_1 FILLER_29_450 ();
 sg13g2_fill_2 FILLER_29_482 ();
 sg13g2_fill_1 FILLER_29_484 ();
 sg13g2_fill_1 FILLER_29_502 ();
 sg13g2_fill_2 FILLER_29_539 ();
 sg13g2_fill_1 FILLER_29_541 ();
 sg13g2_fill_1 FILLER_29_549 ();
 sg13g2_fill_1 FILLER_29_561 ();
 sg13g2_fill_2 FILLER_29_597 ();
 sg13g2_fill_1 FILLER_29_599 ();
 sg13g2_fill_2 FILLER_29_605 ();
 sg13g2_fill_2 FILLER_29_652 ();
 sg13g2_fill_2 FILLER_29_667 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_fill_2 FILLER_29_838 ();
 sg13g2_fill_1 FILLER_29_840 ();
 sg13g2_fill_2 FILLER_29_930 ();
 sg13g2_fill_2 FILLER_29_937 ();
 sg13g2_fill_2 FILLER_29_1037 ();
 sg13g2_fill_2 FILLER_29_1048 ();
 sg13g2_fill_2 FILLER_29_1092 ();
 sg13g2_fill_1 FILLER_29_1094 ();
 sg13g2_fill_2 FILLER_29_1121 ();
 sg13g2_fill_1 FILLER_29_1131 ();
 sg13g2_fill_1 FILLER_29_1163 ();
 sg13g2_fill_2 FILLER_29_1169 ();
 sg13g2_fill_1 FILLER_29_1171 ();
 sg13g2_fill_2 FILLER_29_1202 ();
 sg13g2_fill_2 FILLER_29_1245 ();
 sg13g2_fill_2 FILLER_29_1268 ();
 sg13g2_fill_2 FILLER_29_1279 ();
 sg13g2_decap_8 FILLER_29_1346 ();
 sg13g2_decap_8 FILLER_29_1353 ();
 sg13g2_decap_4 FILLER_29_1440 ();
 sg13g2_fill_1 FILLER_29_1444 ();
 sg13g2_fill_1 FILLER_29_1472 ();
 sg13g2_fill_2 FILLER_29_1487 ();
 sg13g2_fill_1 FILLER_29_1489 ();
 sg13g2_fill_1 FILLER_29_1507 ();
 sg13g2_decap_4 FILLER_29_1549 ();
 sg13g2_decap_4 FILLER_29_1577 ();
 sg13g2_fill_1 FILLER_29_1581 ();
 sg13g2_decap_4 FILLER_29_1590 ();
 sg13g2_fill_1 FILLER_29_1594 ();
 sg13g2_fill_2 FILLER_29_1599 ();
 sg13g2_fill_1 FILLER_29_1601 ();
 sg13g2_fill_2 FILLER_29_1632 ();
 sg13g2_fill_2 FILLER_29_1670 ();
 sg13g2_fill_1 FILLER_29_1754 ();
 sg13g2_fill_2 FILLER_29_1791 ();
 sg13g2_fill_1 FILLER_29_1818 ();
 sg13g2_fill_1 FILLER_29_1870 ();
 sg13g2_fill_2 FILLER_29_1877 ();
 sg13g2_fill_1 FILLER_29_1879 ();
 sg13g2_fill_1 FILLER_29_1895 ();
 sg13g2_fill_2 FILLER_29_1902 ();
 sg13g2_fill_2 FILLER_29_1926 ();
 sg13g2_fill_1 FILLER_29_1928 ();
 sg13g2_fill_2 FILLER_29_1983 ();
 sg13g2_fill_1 FILLER_29_1985 ();
 sg13g2_fill_1 FILLER_29_2027 ();
 sg13g2_fill_1 FILLER_29_2068 ();
 sg13g2_fill_1 FILLER_29_2095 ();
 sg13g2_fill_2 FILLER_29_2122 ();
 sg13g2_fill_2 FILLER_29_2153 ();
 sg13g2_fill_1 FILLER_29_2155 ();
 sg13g2_fill_1 FILLER_29_2173 ();
 sg13g2_fill_2 FILLER_29_2180 ();
 sg13g2_fill_2 FILLER_29_2207 ();
 sg13g2_fill_1 FILLER_29_2209 ();
 sg13g2_fill_2 FILLER_29_2224 ();
 sg13g2_fill_2 FILLER_29_2265 ();
 sg13g2_fill_1 FILLER_29_2288 ();
 sg13g2_fill_2 FILLER_29_2315 ();
 sg13g2_fill_2 FILLER_29_2329 ();
 sg13g2_fill_2 FILLER_29_2339 ();
 sg13g2_fill_1 FILLER_29_2341 ();
 sg13g2_decap_4 FILLER_29_2364 ();
 sg13g2_fill_1 FILLER_29_2368 ();
 sg13g2_fill_2 FILLER_29_2405 ();
 sg13g2_fill_1 FILLER_29_2407 ();
 sg13g2_fill_2 FILLER_29_2418 ();
 sg13g2_fill_2 FILLER_29_2425 ();
 sg13g2_fill_1 FILLER_29_2437 ();
 sg13g2_fill_1 FILLER_29_2443 ();
 sg13g2_fill_2 FILLER_29_2454 ();
 sg13g2_fill_1 FILLER_29_2456 ();
 sg13g2_fill_2 FILLER_29_2467 ();
 sg13g2_fill_2 FILLER_29_2493 ();
 sg13g2_decap_4 FILLER_29_2590 ();
 sg13g2_fill_1 FILLER_29_2594 ();
 sg13g2_fill_1 FILLER_29_2656 ();
 sg13g2_decap_4 FILLER_29_2670 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_36 ();
 sg13g2_fill_1 FILLER_30_38 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_2 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_30_434 ();
 sg13g2_fill_1 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_479 ();
 sg13g2_fill_1 FILLER_30_481 ();
 sg13g2_fill_1 FILLER_30_556 ();
 sg13g2_fill_2 FILLER_30_583 ();
 sg13g2_fill_1 FILLER_30_599 ();
 sg13g2_fill_1 FILLER_30_669 ();
 sg13g2_fill_2 FILLER_30_693 ();
 sg13g2_fill_2 FILLER_30_727 ();
 sg13g2_fill_1 FILLER_30_729 ();
 sg13g2_fill_1 FILLER_30_747 ();
 sg13g2_fill_1 FILLER_30_771 ();
 sg13g2_fill_2 FILLER_30_792 ();
 sg13g2_fill_1 FILLER_30_807 ();
 sg13g2_fill_2 FILLER_30_838 ();
 sg13g2_fill_1 FILLER_30_840 ();
 sg13g2_fill_2 FILLER_30_859 ();
 sg13g2_fill_1 FILLER_30_870 ();
 sg13g2_fill_2 FILLER_30_899 ();
 sg13g2_fill_2 FILLER_30_910 ();
 sg13g2_fill_1 FILLER_30_921 ();
 sg13g2_fill_1 FILLER_30_939 ();
 sg13g2_fill_1 FILLER_30_966 ();
 sg13g2_fill_2 FILLER_30_977 ();
 sg13g2_fill_2 FILLER_30_997 ();
 sg13g2_fill_1 FILLER_30_1004 ();
 sg13g2_fill_2 FILLER_30_1132 ();
 sg13g2_fill_2 FILLER_30_1149 ();
 sg13g2_fill_2 FILLER_30_1161 ();
 sg13g2_fill_1 FILLER_30_1163 ();
 sg13g2_fill_1 FILLER_30_1204 ();
 sg13g2_decap_8 FILLER_30_1241 ();
 sg13g2_decap_8 FILLER_30_1248 ();
 sg13g2_fill_1 FILLER_30_1255 ();
 sg13g2_fill_2 FILLER_30_1306 ();
 sg13g2_fill_2 FILLER_30_1360 ();
 sg13g2_fill_1 FILLER_30_1362 ();
 sg13g2_decap_4 FILLER_30_1424 ();
 sg13g2_fill_2 FILLER_30_1446 ();
 sg13g2_fill_1 FILLER_30_1448 ();
 sg13g2_fill_2 FILLER_30_1463 ();
 sg13g2_decap_4 FILLER_30_1473 ();
 sg13g2_decap_8 FILLER_30_1504 ();
 sg13g2_decap_8 FILLER_30_1511 ();
 sg13g2_decap_4 FILLER_30_1558 ();
 sg13g2_fill_1 FILLER_30_1666 ();
 sg13g2_fill_2 FILLER_30_1686 ();
 sg13g2_decap_8 FILLER_30_1698 ();
 sg13g2_fill_2 FILLER_30_1735 ();
 sg13g2_decap_4 FILLER_30_1751 ();
 sg13g2_fill_1 FILLER_30_1818 ();
 sg13g2_fill_2 FILLER_30_1855 ();
 sg13g2_fill_2 FILLER_30_1869 ();
 sg13g2_fill_1 FILLER_30_1871 ();
 sg13g2_fill_2 FILLER_30_1918 ();
 sg13g2_fill_2 FILLER_30_1963 ();
 sg13g2_fill_1 FILLER_30_1965 ();
 sg13g2_fill_1 FILLER_30_2007 ();
 sg13g2_fill_2 FILLER_30_2043 ();
 sg13g2_fill_2 FILLER_30_2061 ();
 sg13g2_fill_1 FILLER_30_2099 ();
 sg13g2_fill_1 FILLER_30_2133 ();
 sg13g2_fill_2 FILLER_30_2153 ();
 sg13g2_fill_1 FILLER_30_2155 ();
 sg13g2_fill_2 FILLER_30_2169 ();
 sg13g2_fill_1 FILLER_30_2171 ();
 sg13g2_fill_2 FILLER_30_2178 ();
 sg13g2_fill_1 FILLER_30_2180 ();
 sg13g2_fill_2 FILLER_30_2189 ();
 sg13g2_fill_1 FILLER_30_2191 ();
 sg13g2_fill_2 FILLER_30_2249 ();
 sg13g2_fill_1 FILLER_30_2321 ();
 sg13g2_fill_1 FILLER_30_2389 ();
 sg13g2_fill_1 FILLER_30_2546 ();
 sg13g2_fill_1 FILLER_30_2565 ();
 sg13g2_fill_1 FILLER_30_2585 ();
 sg13g2_fill_2 FILLER_30_2633 ();
 sg13g2_decap_4 FILLER_30_2670 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_decap_4 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_22 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_fill_1 FILLER_31_457 ();
 sg13g2_fill_1 FILLER_31_481 ();
 sg13g2_fill_2 FILLER_31_491 ();
 sg13g2_fill_1 FILLER_31_493 ();
 sg13g2_fill_1 FILLER_31_507 ();
 sg13g2_fill_2 FILLER_31_518 ();
 sg13g2_fill_1 FILLER_31_529 ();
 sg13g2_fill_2 FILLER_31_572 ();
 sg13g2_fill_1 FILLER_31_574 ();
 sg13g2_fill_2 FILLER_31_596 ();
 sg13g2_fill_1 FILLER_31_603 ();
 sg13g2_decap_4 FILLER_31_617 ();
 sg13g2_fill_1 FILLER_31_621 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_fill_2 FILLER_31_649 ();
 sg13g2_fill_1 FILLER_31_651 ();
 sg13g2_fill_2 FILLER_31_657 ();
 sg13g2_fill_1 FILLER_31_659 ();
 sg13g2_fill_1 FILLER_31_669 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_fill_1 FILLER_31_698 ();
 sg13g2_fill_2 FILLER_31_725 ();
 sg13g2_fill_2 FILLER_31_847 ();
 sg13g2_fill_2 FILLER_31_875 ();
 sg13g2_fill_2 FILLER_31_935 ();
 sg13g2_fill_1 FILLER_31_963 ();
 sg13g2_fill_1 FILLER_31_1020 ();
 sg13g2_fill_2 FILLER_31_1039 ();
 sg13g2_fill_2 FILLER_31_1050 ();
 sg13g2_fill_1 FILLER_31_1052 ();
 sg13g2_fill_2 FILLER_31_1067 ();
 sg13g2_fill_1 FILLER_31_1069 ();
 sg13g2_fill_1 FILLER_31_1084 ();
 sg13g2_fill_2 FILLER_31_1125 ();
 sg13g2_fill_2 FILLER_31_1153 ();
 sg13g2_fill_1 FILLER_31_1155 ();
 sg13g2_fill_2 FILLER_31_1182 ();
 sg13g2_fill_1 FILLER_31_1184 ();
 sg13g2_decap_8 FILLER_31_1208 ();
 sg13g2_decap_8 FILLER_31_1232 ();
 sg13g2_fill_2 FILLER_31_1245 ();
 sg13g2_fill_2 FILLER_31_1269 ();
 sg13g2_fill_1 FILLER_31_1271 ();
 sg13g2_fill_2 FILLER_31_1336 ();
 sg13g2_fill_1 FILLER_31_1352 ();
 sg13g2_fill_1 FILLER_31_1362 ();
 sg13g2_fill_1 FILLER_31_1372 ();
 sg13g2_fill_2 FILLER_31_1406 ();
 sg13g2_decap_4 FILLER_31_1470 ();
 sg13g2_fill_1 FILLER_31_1474 ();
 sg13g2_fill_2 FILLER_31_1485 ();
 sg13g2_fill_1 FILLER_31_1487 ();
 sg13g2_fill_1 FILLER_31_1497 ();
 sg13g2_decap_4 FILLER_31_1519 ();
 sg13g2_fill_1 FILLER_31_1523 ();
 sg13g2_decap_4 FILLER_31_1537 ();
 sg13g2_fill_2 FILLER_31_1541 ();
 sg13g2_decap_4 FILLER_31_1547 ();
 sg13g2_fill_1 FILLER_31_1551 ();
 sg13g2_fill_2 FILLER_31_1562 ();
 sg13g2_fill_2 FILLER_31_1587 ();
 sg13g2_fill_1 FILLER_31_1639 ();
 sg13g2_decap_4 FILLER_31_1666 ();
 sg13g2_fill_2 FILLER_31_1771 ();
 sg13g2_fill_1 FILLER_31_1773 ();
 sg13g2_fill_2 FILLER_31_1784 ();
 sg13g2_fill_1 FILLER_31_1786 ();
 sg13g2_fill_2 FILLER_31_1792 ();
 sg13g2_fill_1 FILLER_31_1794 ();
 sg13g2_decap_8 FILLER_31_1800 ();
 sg13g2_fill_2 FILLER_31_1821 ();
 sg13g2_decap_8 FILLER_31_1856 ();
 sg13g2_fill_1 FILLER_31_1863 ();
 sg13g2_fill_2 FILLER_31_1872 ();
 sg13g2_fill_1 FILLER_31_1874 ();
 sg13g2_fill_2 FILLER_31_1890 ();
 sg13g2_fill_2 FILLER_31_1913 ();
 sg13g2_fill_1 FILLER_31_1915 ();
 sg13g2_decap_4 FILLER_31_1942 ();
 sg13g2_fill_1 FILLER_31_1946 ();
 sg13g2_fill_2 FILLER_31_1976 ();
 sg13g2_fill_1 FILLER_31_1978 ();
 sg13g2_fill_1 FILLER_31_1994 ();
 sg13g2_fill_1 FILLER_31_2071 ();
 sg13g2_fill_1 FILLER_31_2088 ();
 sg13g2_fill_1 FILLER_31_2138 ();
 sg13g2_fill_1 FILLER_31_2147 ();
 sg13g2_fill_2 FILLER_31_2192 ();
 sg13g2_fill_2 FILLER_31_2216 ();
 sg13g2_fill_1 FILLER_31_2218 ();
 sg13g2_fill_2 FILLER_31_2237 ();
 sg13g2_fill_1 FILLER_31_2239 ();
 sg13g2_fill_2 FILLER_31_2275 ();
 sg13g2_fill_2 FILLER_31_2292 ();
 sg13g2_fill_1 FILLER_31_2294 ();
 sg13g2_fill_2 FILLER_31_2333 ();
 sg13g2_fill_1 FILLER_31_2335 ();
 sg13g2_decap_4 FILLER_31_2348 ();
 sg13g2_fill_2 FILLER_31_2450 ();
 sg13g2_fill_1 FILLER_31_2469 ();
 sg13g2_fill_2 FILLER_31_2491 ();
 sg13g2_fill_1 FILLER_31_2493 ();
 sg13g2_fill_2 FILLER_31_2508 ();
 sg13g2_fill_2 FILLER_31_2542 ();
 sg13g2_decap_8 FILLER_31_2556 ();
 sg13g2_fill_1 FILLER_31_2563 ();
 sg13g2_decap_4 FILLER_31_2653 ();
 sg13g2_decap_4 FILLER_31_2670 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_24 ();
 sg13g2_decap_4 FILLER_32_31 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_169 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_369 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_443 ();
 sg13g2_fill_1 FILLER_32_476 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_1 FILLER_32_675 ();
 sg13g2_decap_8 FILLER_32_685 ();
 sg13g2_decap_4 FILLER_32_692 ();
 sg13g2_fill_1 FILLER_32_696 ();
 sg13g2_fill_2 FILLER_32_724 ();
 sg13g2_fill_1 FILLER_32_726 ();
 sg13g2_fill_2 FILLER_32_740 ();
 sg13g2_fill_1 FILLER_32_742 ();
 sg13g2_fill_2 FILLER_32_752 ();
 sg13g2_fill_1 FILLER_32_770 ();
 sg13g2_fill_2 FILLER_32_889 ();
 sg13g2_fill_2 FILLER_32_907 ();
 sg13g2_fill_1 FILLER_32_909 ();
 sg13g2_fill_2 FILLER_32_915 ();
 sg13g2_fill_2 FILLER_32_986 ();
 sg13g2_fill_2 FILLER_32_1007 ();
 sg13g2_fill_2 FILLER_32_1028 ();
 sg13g2_fill_1 FILLER_32_1030 ();
 sg13g2_fill_2 FILLER_32_1082 ();
 sg13g2_fill_1 FILLER_32_1120 ();
 sg13g2_decap_4 FILLER_32_1178 ();
 sg13g2_fill_1 FILLER_32_1182 ();
 sg13g2_fill_2 FILLER_32_1235 ();
 sg13g2_decap_4 FILLER_32_1251 ();
 sg13g2_fill_1 FILLER_32_1259 ();
 sg13g2_fill_1 FILLER_32_1298 ();
 sg13g2_decap_4 FILLER_32_1304 ();
 sg13g2_fill_1 FILLER_32_1308 ();
 sg13g2_decap_4 FILLER_32_1391 ();
 sg13g2_decap_8 FILLER_32_1403 ();
 sg13g2_decap_4 FILLER_32_1410 ();
 sg13g2_decap_4 FILLER_32_1423 ();
 sg13g2_fill_2 FILLER_32_1427 ();
 sg13g2_fill_2 FILLER_32_1450 ();
 sg13g2_fill_1 FILLER_32_1452 ();
 sg13g2_fill_2 FILLER_32_1466 ();
 sg13g2_decap_8 FILLER_32_1478 ();
 sg13g2_fill_1 FILLER_32_1549 ();
 sg13g2_decap_4 FILLER_32_1566 ();
 sg13g2_fill_2 FILLER_32_1616 ();
 sg13g2_decap_8 FILLER_32_1622 ();
 sg13g2_fill_2 FILLER_32_1629 ();
 sg13g2_fill_2 FILLER_32_1635 ();
 sg13g2_fill_1 FILLER_32_1637 ();
 sg13g2_decap_8 FILLER_32_1644 ();
 sg13g2_decap_8 FILLER_32_1671 ();
 sg13g2_fill_2 FILLER_32_1678 ();
 sg13g2_decap_8 FILLER_32_1693 ();
 sg13g2_fill_1 FILLER_32_1700 ();
 sg13g2_fill_2 FILLER_32_1705 ();
 sg13g2_fill_1 FILLER_32_1716 ();
 sg13g2_fill_1 FILLER_32_1753 ();
 sg13g2_fill_2 FILLER_32_1831 ();
 sg13g2_decap_4 FILLER_32_1864 ();
 sg13g2_fill_2 FILLER_32_1868 ();
 sg13g2_fill_2 FILLER_32_1896 ();
 sg13g2_fill_2 FILLER_32_1924 ();
 sg13g2_fill_1 FILLER_32_1926 ();
 sg13g2_decap_8 FILLER_32_1935 ();
 sg13g2_decap_8 FILLER_32_1942 ();
 sg13g2_decap_8 FILLER_32_1949 ();
 sg13g2_fill_1 FILLER_32_1956 ();
 sg13g2_fill_2 FILLER_32_1996 ();
 sg13g2_fill_2 FILLER_32_2034 ();
 sg13g2_fill_1 FILLER_32_2049 ();
 sg13g2_decap_4 FILLER_32_2055 ();
 sg13g2_fill_1 FILLER_32_2106 ();
 sg13g2_fill_1 FILLER_32_2162 ();
 sg13g2_fill_2 FILLER_32_2229 ();
 sg13g2_fill_1 FILLER_32_2320 ();
 sg13g2_fill_2 FILLER_32_2367 ();
 sg13g2_fill_1 FILLER_32_2388 ();
 sg13g2_fill_1 FILLER_32_2432 ();
 sg13g2_decap_4 FILLER_32_2454 ();
 sg13g2_fill_2 FILLER_32_2458 ();
 sg13g2_fill_1 FILLER_32_2464 ();
 sg13g2_fill_1 FILLER_32_2551 ();
 sg13g2_fill_2 FILLER_32_2582 ();
 sg13g2_fill_1 FILLER_32_2584 ();
 sg13g2_fill_2 FILLER_32_2634 ();
 sg13g2_fill_1 FILLER_32_2636 ();
 sg13g2_fill_1 FILLER_32_2647 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_24 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_54 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_decap_4 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_435 ();
 sg13g2_fill_2 FILLER_33_454 ();
 sg13g2_fill_2 FILLER_33_465 ();
 sg13g2_fill_1 FILLER_33_467 ();
 sg13g2_fill_2 FILLER_33_478 ();
 sg13g2_decap_8 FILLER_33_500 ();
 sg13g2_decap_8 FILLER_33_524 ();
 sg13g2_decap_4 FILLER_33_535 ();
 sg13g2_fill_1 FILLER_33_539 ();
 sg13g2_fill_2 FILLER_33_563 ();
 sg13g2_fill_1 FILLER_33_565 ();
 sg13g2_decap_8 FILLER_33_596 ();
 sg13g2_fill_2 FILLER_33_616 ();
 sg13g2_decap_4 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_658 ();
 sg13g2_fill_2 FILLER_33_664 ();
 sg13g2_fill_2 FILLER_33_674 ();
 sg13g2_decap_4 FILLER_33_682 ();
 sg13g2_fill_2 FILLER_33_730 ();
 sg13g2_fill_2 FILLER_33_767 ();
 sg13g2_fill_2 FILLER_33_778 ();
 sg13g2_fill_1 FILLER_33_780 ();
 sg13g2_fill_2 FILLER_33_786 ();
 sg13g2_fill_1 FILLER_33_788 ();
 sg13g2_fill_2 FILLER_33_794 ();
 sg13g2_fill_1 FILLER_33_796 ();
 sg13g2_fill_2 FILLER_33_801 ();
 sg13g2_fill_2 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_813 ();
 sg13g2_fill_2 FILLER_33_823 ();
 sg13g2_fill_2 FILLER_33_834 ();
 sg13g2_fill_1 FILLER_33_836 ();
 sg13g2_fill_1 FILLER_33_846 ();
 sg13g2_fill_2 FILLER_33_934 ();
 sg13g2_fill_1 FILLER_33_936 ();
 sg13g2_fill_2 FILLER_33_1007 ();
 sg13g2_fill_1 FILLER_33_1009 ();
 sg13g2_fill_2 FILLER_33_1072 ();
 sg13g2_fill_2 FILLER_33_1127 ();
 sg13g2_fill_2 FILLER_33_1195 ();
 sg13g2_fill_1 FILLER_33_1197 ();
 sg13g2_fill_2 FILLER_33_1234 ();
 sg13g2_fill_1 FILLER_33_1236 ();
 sg13g2_fill_1 FILLER_33_1270 ();
 sg13g2_decap_4 FILLER_33_1277 ();
 sg13g2_fill_2 FILLER_33_1281 ();
 sg13g2_decap_4 FILLER_33_1312 ();
 sg13g2_fill_1 FILLER_33_1316 ();
 sg13g2_decap_8 FILLER_33_1322 ();
 sg13g2_fill_1 FILLER_33_1329 ();
 sg13g2_decap_4 FILLER_33_1334 ();
 sg13g2_fill_1 FILLER_33_1338 ();
 sg13g2_decap_8 FILLER_33_1344 ();
 sg13g2_decap_4 FILLER_33_1351 ();
 sg13g2_fill_2 FILLER_33_1355 ();
 sg13g2_fill_1 FILLER_33_1362 ();
 sg13g2_fill_1 FILLER_33_1379 ();
 sg13g2_fill_1 FILLER_33_1406 ();
 sg13g2_decap_4 FILLER_33_1433 ();
 sg13g2_decap_4 FILLER_33_1458 ();
 sg13g2_fill_1 FILLER_33_1462 ();
 sg13g2_fill_2 FILLER_33_1534 ();
 sg13g2_fill_1 FILLER_33_1536 ();
 sg13g2_decap_4 FILLER_33_1551 ();
 sg13g2_fill_2 FILLER_33_1569 ();
 sg13g2_fill_1 FILLER_33_1571 ();
 sg13g2_fill_2 FILLER_33_1586 ();
 sg13g2_fill_1 FILLER_33_1653 ();
 sg13g2_fill_1 FILLER_33_1680 ();
 sg13g2_decap_4 FILLER_33_1696 ();
 sg13g2_fill_2 FILLER_33_1725 ();
 sg13g2_fill_1 FILLER_33_1727 ();
 sg13g2_fill_2 FILLER_33_1748 ();
 sg13g2_fill_2 FILLER_33_1776 ();
 sg13g2_fill_1 FILLER_33_1778 ();
 sg13g2_fill_1 FILLER_33_1800 ();
 sg13g2_fill_2 FILLER_33_1853 ();
 sg13g2_decap_8 FILLER_33_1872 ();
 sg13g2_fill_1 FILLER_33_1902 ();
 sg13g2_fill_1 FILLER_33_1926 ();
 sg13g2_fill_2 FILLER_33_1935 ();
 sg13g2_decap_8 FILLER_33_1953 ();
 sg13g2_fill_2 FILLER_33_1960 ();
 sg13g2_fill_2 FILLER_33_1966 ();
 sg13g2_fill_1 FILLER_33_1991 ();
 sg13g2_decap_4 FILLER_33_2015 ();
 sg13g2_fill_1 FILLER_33_2023 ();
 sg13g2_fill_2 FILLER_33_2048 ();
 sg13g2_fill_1 FILLER_33_2050 ();
 sg13g2_fill_2 FILLER_33_2083 ();
 sg13g2_fill_1 FILLER_33_2085 ();
 sg13g2_fill_2 FILLER_33_2135 ();
 sg13g2_fill_1 FILLER_33_2154 ();
 sg13g2_fill_2 FILLER_33_2238 ();
 sg13g2_fill_2 FILLER_33_2270 ();
 sg13g2_fill_1 FILLER_33_2272 ();
 sg13g2_fill_1 FILLER_33_2278 ();
 sg13g2_decap_4 FILLER_33_2315 ();
 sg13g2_fill_2 FILLER_33_2319 ();
 sg13g2_fill_1 FILLER_33_2345 ();
 sg13g2_fill_1 FILLER_33_2365 ();
 sg13g2_fill_1 FILLER_33_2380 ();
 sg13g2_fill_2 FILLER_33_2400 ();
 sg13g2_fill_1 FILLER_33_2402 ();
 sg13g2_fill_1 FILLER_33_2408 ();
 sg13g2_fill_2 FILLER_33_2423 ();
 sg13g2_fill_2 FILLER_33_2484 ();
 sg13g2_fill_1 FILLER_33_2536 ();
 sg13g2_fill_1 FILLER_33_2558 ();
 sg13g2_fill_2 FILLER_33_2564 ();
 sg13g2_fill_2 FILLER_33_2570 ();
 sg13g2_fill_1 FILLER_33_2572 ();
 sg13g2_fill_1 FILLER_33_2647 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_11 ();
 sg13g2_fill_2 FILLER_34_23 ();
 sg13g2_fill_1 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_fill_2 FILLER_34_398 ();
 sg13g2_fill_1 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_fill_2 FILLER_34_470 ();
 sg13g2_fill_1 FILLER_34_472 ();
 sg13g2_decap_8 FILLER_34_499 ();
 sg13g2_fill_1 FILLER_34_545 ();
 sg13g2_fill_1 FILLER_34_625 ();
 sg13g2_decap_4 FILLER_34_660 ();
 sg13g2_fill_2 FILLER_34_741 ();
 sg13g2_fill_2 FILLER_34_783 ();
 sg13g2_fill_1 FILLER_34_785 ();
 sg13g2_fill_1 FILLER_34_887 ();
 sg13g2_fill_2 FILLER_34_923 ();
 sg13g2_fill_1 FILLER_34_962 ();
 sg13g2_fill_1 FILLER_34_968 ();
 sg13g2_fill_2 FILLER_34_1025 ();
 sg13g2_fill_2 FILLER_34_1041 ();
 sg13g2_fill_1 FILLER_34_1103 ();
 sg13g2_fill_2 FILLER_34_1117 ();
 sg13g2_fill_1 FILLER_34_1145 ();
 sg13g2_fill_2 FILLER_34_1151 ();
 sg13g2_fill_2 FILLER_34_1157 ();
 sg13g2_fill_1 FILLER_34_1159 ();
 sg13g2_fill_1 FILLER_34_1164 ();
 sg13g2_decap_4 FILLER_34_1193 ();
 sg13g2_fill_1 FILLER_34_1197 ();
 sg13g2_decap_8 FILLER_34_1210 ();
 sg13g2_fill_1 FILLER_34_1217 ();
 sg13g2_decap_4 FILLER_34_1236 ();
 sg13g2_fill_2 FILLER_34_1307 ();
 sg13g2_fill_2 FILLER_34_1330 ();
 sg13g2_fill_1 FILLER_34_1332 ();
 sg13g2_fill_2 FILLER_34_1338 ();
 sg13g2_fill_1 FILLER_34_1350 ();
 sg13g2_fill_1 FILLER_34_1369 ();
 sg13g2_fill_1 FILLER_34_1389 ();
 sg13g2_fill_1 FILLER_34_1394 ();
 sg13g2_fill_1 FILLER_34_1404 ();
 sg13g2_decap_4 FILLER_34_1434 ();
 sg13g2_fill_1 FILLER_34_1460 ();
 sg13g2_fill_1 FILLER_34_1472 ();
 sg13g2_fill_2 FILLER_34_1492 ();
 sg13g2_fill_2 FILLER_34_1511 ();
 sg13g2_decap_4 FILLER_34_1557 ();
 sg13g2_fill_2 FILLER_34_1561 ();
 sg13g2_decap_4 FILLER_34_1569 ();
 sg13g2_fill_1 FILLER_34_1573 ();
 sg13g2_decap_4 FILLER_34_1583 ();
 sg13g2_decap_4 FILLER_34_1603 ();
 sg13g2_decap_8 FILLER_34_1611 ();
 sg13g2_fill_2 FILLER_34_1618 ();
 sg13g2_fill_2 FILLER_34_1634 ();
 sg13g2_decap_8 FILLER_34_1685 ();
 sg13g2_decap_4 FILLER_34_1718 ();
 sg13g2_fill_1 FILLER_34_1722 ();
 sg13g2_decap_4 FILLER_34_1749 ();
 sg13g2_decap_8 FILLER_34_1802 ();
 sg13g2_decap_4 FILLER_34_1809 ();
 sg13g2_fill_2 FILLER_34_1813 ();
 sg13g2_fill_2 FILLER_34_1859 ();
 sg13g2_decap_4 FILLER_34_1998 ();
 sg13g2_decap_8 FILLER_34_2006 ();
 sg13g2_fill_1 FILLER_34_2013 ();
 sg13g2_fill_1 FILLER_34_2041 ();
 sg13g2_fill_1 FILLER_34_2048 ();
 sg13g2_fill_2 FILLER_34_2076 ();
 sg13g2_fill_1 FILLER_34_2078 ();
 sg13g2_fill_1 FILLER_34_2124 ();
 sg13g2_decap_8 FILLER_34_2173 ();
 sg13g2_fill_2 FILLER_34_2180 ();
 sg13g2_fill_2 FILLER_34_2202 ();
 sg13g2_fill_2 FILLER_34_2212 ();
 sg13g2_fill_1 FILLER_34_2214 ();
 sg13g2_fill_2 FILLER_34_2229 ();
 sg13g2_fill_1 FILLER_34_2231 ();
 sg13g2_fill_2 FILLER_34_2268 ();
 sg13g2_fill_1 FILLER_34_2270 ();
 sg13g2_fill_1 FILLER_34_2275 ();
 sg13g2_fill_2 FILLER_34_2281 ();
 sg13g2_fill_1 FILLER_34_2283 ();
 sg13g2_fill_1 FILLER_34_2320 ();
 sg13g2_fill_2 FILLER_34_2370 ();
 sg13g2_fill_2 FILLER_34_2424 ();
 sg13g2_fill_1 FILLER_34_2466 ();
 sg13g2_fill_1 FILLER_34_2495 ();
 sg13g2_fill_1 FILLER_34_2554 ();
 sg13g2_fill_2 FILLER_34_2581 ();
 sg13g2_fill_2 FILLER_34_2622 ();
 sg13g2_fill_1 FILLER_34_2673 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_15 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_decap_8 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_fill_2 FILLER_35_66 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_decap_4 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_321 ();
 sg13g2_decap_4 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_fill_2 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_fill_1 FILLER_35_421 ();
 sg13g2_fill_1 FILLER_35_435 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_466 ();
 sg13g2_fill_1 FILLER_35_468 ();
 sg13g2_fill_2 FILLER_35_490 ();
 sg13g2_fill_2 FILLER_35_557 ();
 sg13g2_decap_8 FILLER_35_594 ();
 sg13g2_fill_1 FILLER_35_601 ();
 sg13g2_fill_1 FILLER_35_606 ();
 sg13g2_fill_2 FILLER_35_623 ();
 sg13g2_fill_1 FILLER_35_625 ();
 sg13g2_fill_2 FILLER_35_647 ();
 sg13g2_fill_1 FILLER_35_649 ();
 sg13g2_decap_4 FILLER_35_662 ();
 sg13g2_fill_2 FILLER_35_666 ();
 sg13g2_decap_4 FILLER_35_674 ();
 sg13g2_fill_2 FILLER_35_678 ();
 sg13g2_fill_1 FILLER_35_723 ();
 sg13g2_fill_2 FILLER_35_758 ();
 sg13g2_fill_1 FILLER_35_760 ();
 sg13g2_fill_1 FILLER_35_863 ();
 sg13g2_fill_1 FILLER_35_873 ();
 sg13g2_fill_2 FILLER_35_904 ();
 sg13g2_fill_1 FILLER_35_906 ();
 sg13g2_fill_2 FILLER_35_968 ();
 sg13g2_fill_2 FILLER_35_1023 ();
 sg13g2_fill_1 FILLER_35_1025 ();
 sg13g2_fill_2 FILLER_35_1057 ();
 sg13g2_fill_1 FILLER_35_1059 ();
 sg13g2_fill_2 FILLER_35_1126 ();
 sg13g2_fill_1 FILLER_35_1136 ();
 sg13g2_fill_2 FILLER_35_1189 ();
 sg13g2_fill_1 FILLER_35_1191 ();
 sg13g2_fill_1 FILLER_35_1228 ();
 sg13g2_decap_4 FILLER_35_1233 ();
 sg13g2_fill_2 FILLER_35_1254 ();
 sg13g2_fill_1 FILLER_35_1256 ();
 sg13g2_fill_2 FILLER_35_1274 ();
 sg13g2_decap_4 FILLER_35_1316 ();
 sg13g2_fill_1 FILLER_35_1320 ();
 sg13g2_fill_1 FILLER_35_1333 ();
 sg13g2_fill_2 FILLER_35_1375 ();
 sg13g2_fill_1 FILLER_35_1377 ();
 sg13g2_fill_2 FILLER_35_1388 ();
 sg13g2_decap_8 FILLER_35_1395 ();
 sg13g2_fill_1 FILLER_35_1402 ();
 sg13g2_fill_2 FILLER_35_1445 ();
 sg13g2_fill_1 FILLER_35_1447 ();
 sg13g2_decap_4 FILLER_35_1454 ();
 sg13g2_fill_2 FILLER_35_1477 ();
 sg13g2_decap_8 FILLER_35_1549 ();
 sg13g2_fill_1 FILLER_35_1556 ();
 sg13g2_decap_4 FILLER_35_1601 ();
 sg13g2_fill_2 FILLER_35_1613 ();
 sg13g2_decap_4 FILLER_35_1619 ();
 sg13g2_fill_2 FILLER_35_1659 ();
 sg13g2_fill_1 FILLER_35_1669 ();
 sg13g2_decap_8 FILLER_35_1709 ();
 sg13g2_fill_2 FILLER_35_1728 ();
 sg13g2_fill_2 FILLER_35_1748 ();
 sg13g2_fill_1 FILLER_35_1760 ();
 sg13g2_decap_4 FILLER_35_1791 ();
 sg13g2_fill_1 FILLER_35_1795 ();
 sg13g2_decap_4 FILLER_35_1830 ();
 sg13g2_fill_2 FILLER_35_1834 ();
 sg13g2_fill_2 FILLER_35_1862 ();
 sg13g2_fill_1 FILLER_35_1980 ();
 sg13g2_decap_4 FILLER_35_2017 ();
 sg13g2_fill_2 FILLER_35_2053 ();
 sg13g2_decap_8 FILLER_35_2102 ();
 sg13g2_fill_2 FILLER_35_2144 ();
 sg13g2_fill_1 FILLER_35_2146 ();
 sg13g2_decap_8 FILLER_35_2160 ();
 sg13g2_fill_1 FILLER_35_2167 ();
 sg13g2_fill_2 FILLER_35_2202 ();
 sg13g2_fill_2 FILLER_35_2251 ();
 sg13g2_fill_1 FILLER_35_2253 ();
 sg13g2_fill_2 FILLER_35_2289 ();
 sg13g2_decap_8 FILLER_35_2317 ();
 sg13g2_fill_2 FILLER_35_2350 ();
 sg13g2_fill_1 FILLER_35_2352 ();
 sg13g2_fill_1 FILLER_35_2414 ();
 sg13g2_fill_1 FILLER_35_2471 ();
 sg13g2_fill_2 FILLER_35_2535 ();
 sg13g2_fill_1 FILLER_35_2618 ();
 sg13g2_decap_8 FILLER_35_2640 ();
 sg13g2_fill_1 FILLER_35_2673 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_2 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_454 ();
 sg13g2_fill_2 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_567 ();
 sg13g2_fill_1 FILLER_36_569 ();
 sg13g2_fill_1 FILLER_36_579 ();
 sg13g2_fill_2 FILLER_36_618 ();
 sg13g2_decap_4 FILLER_36_633 ();
 sg13g2_fill_2 FILLER_36_643 ();
 sg13g2_fill_2 FILLER_36_656 ();
 sg13g2_fill_1 FILLER_36_658 ();
 sg13g2_fill_2 FILLER_36_671 ();
 sg13g2_decap_4 FILLER_36_681 ();
 sg13g2_fill_2 FILLER_36_720 ();
 sg13g2_fill_1 FILLER_36_722 ();
 sg13g2_fill_2 FILLER_36_759 ();
 sg13g2_fill_1 FILLER_36_774 ();
 sg13g2_decap_4 FILLER_36_802 ();
 sg13g2_fill_1 FILLER_36_806 ();
 sg13g2_decap_4 FILLER_36_811 ();
 sg13g2_fill_2 FILLER_36_815 ();
 sg13g2_fill_1 FILLER_36_830 ();
 sg13g2_fill_2 FILLER_36_842 ();
 sg13g2_fill_1 FILLER_36_880 ();
 sg13g2_decap_8 FILLER_36_904 ();
 sg13g2_decap_4 FILLER_36_924 ();
 sg13g2_fill_1 FILLER_36_928 ();
 sg13g2_fill_2 FILLER_36_945 ();
 sg13g2_decap_4 FILLER_36_956 ();
 sg13g2_fill_1 FILLER_36_960 ();
 sg13g2_decap_4 FILLER_36_975 ();
 sg13g2_fill_2 FILLER_36_979 ();
 sg13g2_decap_8 FILLER_36_989 ();
 sg13g2_fill_2 FILLER_36_1009 ();
 sg13g2_fill_1 FILLER_36_1011 ();
 sg13g2_decap_4 FILLER_36_1052 ();
 sg13g2_fill_1 FILLER_36_1056 ();
 sg13g2_fill_2 FILLER_36_1067 ();
 sg13g2_fill_1 FILLER_36_1069 ();
 sg13g2_fill_2 FILLER_36_1123 ();
 sg13g2_fill_1 FILLER_36_1125 ();
 sg13g2_fill_2 FILLER_36_1138 ();
 sg13g2_fill_1 FILLER_36_1140 ();
 sg13g2_fill_2 FILLER_36_1164 ();
 sg13g2_fill_1 FILLER_36_1166 ();
 sg13g2_fill_2 FILLER_36_1180 ();
 sg13g2_fill_1 FILLER_36_1197 ();
 sg13g2_decap_4 FILLER_36_1234 ();
 sg13g2_fill_2 FILLER_36_1288 ();
 sg13g2_fill_1 FILLER_36_1290 ();
 sg13g2_fill_2 FILLER_36_1332 ();
 sg13g2_fill_2 FILLER_36_1339 ();
 sg13g2_fill_1 FILLER_36_1341 ();
 sg13g2_decap_8 FILLER_36_1350 ();
 sg13g2_fill_2 FILLER_36_1357 ();
 sg13g2_fill_2 FILLER_36_1374 ();
 sg13g2_fill_2 FILLER_36_1439 ();
 sg13g2_decap_8 FILLER_36_1489 ();
 sg13g2_decap_4 FILLER_36_1496 ();
 sg13g2_fill_1 FILLER_36_1500 ();
 sg13g2_fill_2 FILLER_36_1517 ();
 sg13g2_fill_1 FILLER_36_1519 ();
 sg13g2_decap_8 FILLER_36_1541 ();
 sg13g2_decap_4 FILLER_36_1560 ();
 sg13g2_fill_1 FILLER_36_1572 ();
 sg13g2_fill_2 FILLER_36_1578 ();
 sg13g2_fill_2 FILLER_36_1630 ();
 sg13g2_fill_1 FILLER_36_1632 ();
 sg13g2_decap_4 FILLER_36_1684 ();
 sg13g2_decap_4 FILLER_36_1780 ();
 sg13g2_decap_4 FILLER_36_1793 ();
 sg13g2_fill_2 FILLER_36_1827 ();
 sg13g2_fill_1 FILLER_36_1829 ();
 sg13g2_fill_2 FILLER_36_1861 ();
 sg13g2_fill_2 FILLER_36_1903 ();
 sg13g2_fill_1 FILLER_36_1905 ();
 sg13g2_fill_2 FILLER_36_2005 ();
 sg13g2_fill_2 FILLER_36_2020 ();
 sg13g2_fill_1 FILLER_36_2022 ();
 sg13g2_fill_1 FILLER_36_2059 ();
 sg13g2_fill_2 FILLER_36_2101 ();
 sg13g2_fill_2 FILLER_36_2128 ();
 sg13g2_fill_1 FILLER_36_2177 ();
 sg13g2_fill_1 FILLER_36_2201 ();
 sg13g2_fill_2 FILLER_36_2220 ();
 sg13g2_decap_8 FILLER_36_2399 ();
 sg13g2_fill_1 FILLER_36_2406 ();
 sg13g2_fill_1 FILLER_36_2436 ();
 sg13g2_fill_2 FILLER_36_2488 ();
 sg13g2_decap_4 FILLER_36_2644 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_11 ();
 sg13g2_fill_2 FILLER_37_61 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_decap_4 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_2 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_decap_4 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_decap_4 FILLER_37_401 ();
 sg13g2_fill_2 FILLER_37_436 ();
 sg13g2_fill_1 FILLER_37_438 ();
 sg13g2_fill_2 FILLER_37_512 ();
 sg13g2_fill_2 FILLER_37_544 ();
 sg13g2_fill_2 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_565 ();
 sg13g2_decap_4 FILLER_37_592 ();
 sg13g2_fill_1 FILLER_37_596 ();
 sg13g2_fill_2 FILLER_37_605 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_1 FILLER_37_675 ();
 sg13g2_fill_1 FILLER_37_682 ();
 sg13g2_fill_1 FILLER_37_691 ();
 sg13g2_fill_1 FILLER_37_717 ();
 sg13g2_fill_1 FILLER_37_724 ();
 sg13g2_decap_4 FILLER_37_733 ();
 sg13g2_fill_2 FILLER_37_737 ();
 sg13g2_fill_1 FILLER_37_743 ();
 sg13g2_fill_2 FILLER_37_748 ();
 sg13g2_fill_1 FILLER_37_772 ();
 sg13g2_fill_2 FILLER_37_786 ();
 sg13g2_fill_2 FILLER_37_837 ();
 sg13g2_fill_1 FILLER_37_839 ();
 sg13g2_fill_1 FILLER_37_846 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_1 FILLER_37_875 ();
 sg13g2_fill_2 FILLER_37_889 ();
 sg13g2_fill_1 FILLER_37_891 ();
 sg13g2_fill_1 FILLER_37_962 ();
 sg13g2_fill_2 FILLER_37_969 ();
 sg13g2_fill_1 FILLER_37_971 ();
 sg13g2_decap_4 FILLER_37_977 ();
 sg13g2_fill_1 FILLER_37_1001 ();
 sg13g2_fill_2 FILLER_37_1011 ();
 sg13g2_fill_2 FILLER_37_1023 ();
 sg13g2_fill_1 FILLER_37_1037 ();
 sg13g2_fill_2 FILLER_37_1084 ();
 sg13g2_fill_1 FILLER_37_1086 ();
 sg13g2_fill_2 FILLER_37_1124 ();
 sg13g2_fill_2 FILLER_37_1137 ();
 sg13g2_decap_4 FILLER_37_1233 ();
 sg13g2_fill_1 FILLER_37_1266 ();
 sg13g2_fill_2 FILLER_37_1298 ();
 sg13g2_fill_1 FILLER_37_1300 ();
 sg13g2_fill_1 FILLER_37_1315 ();
 sg13g2_fill_2 FILLER_37_1406 ();
 sg13g2_fill_1 FILLER_37_1414 ();
 sg13g2_fill_1 FILLER_37_1420 ();
 sg13g2_decap_8 FILLER_37_1446 ();
 sg13g2_decap_8 FILLER_37_1462 ();
 sg13g2_decap_8 FILLER_37_1469 ();
 sg13g2_fill_2 FILLER_37_1516 ();
 sg13g2_fill_1 FILLER_37_1518 ();
 sg13g2_fill_1 FILLER_37_1528 ();
 sg13g2_fill_1 FILLER_37_1553 ();
 sg13g2_fill_1 FILLER_37_1559 ();
 sg13g2_fill_2 FILLER_37_1590 ();
 sg13g2_fill_1 FILLER_37_1592 ();
 sg13g2_fill_1 FILLER_37_1635 ();
 sg13g2_fill_2 FILLER_37_1651 ();
 sg13g2_fill_1 FILLER_37_1653 ();
 sg13g2_decap_4 FILLER_37_1727 ();
 sg13g2_fill_2 FILLER_37_1731 ();
 sg13g2_fill_1 FILLER_37_1755 ();
 sg13g2_fill_1 FILLER_37_1782 ();
 sg13g2_fill_2 FILLER_37_1803 ();
 sg13g2_fill_2 FILLER_37_1863 ();
 sg13g2_fill_2 FILLER_37_1889 ();
 sg13g2_decap_4 FILLER_37_1934 ();
 sg13g2_fill_1 FILLER_37_1938 ();
 sg13g2_fill_2 FILLER_37_1965 ();
 sg13g2_fill_2 FILLER_37_2032 ();
 sg13g2_fill_1 FILLER_37_2042 ();
 sg13g2_fill_2 FILLER_37_2052 ();
 sg13g2_fill_1 FILLER_37_2054 ();
 sg13g2_fill_1 FILLER_37_2065 ();
 sg13g2_fill_2 FILLER_37_2081 ();
 sg13g2_fill_1 FILLER_37_2083 ();
 sg13g2_fill_1 FILLER_37_2129 ();
 sg13g2_decap_4 FILLER_37_2184 ();
 sg13g2_fill_2 FILLER_37_2188 ();
 sg13g2_fill_1 FILLER_37_2242 ();
 sg13g2_fill_2 FILLER_37_2279 ();
 sg13g2_fill_1 FILLER_37_2281 ();
 sg13g2_fill_2 FILLER_37_2301 ();
 sg13g2_fill_2 FILLER_37_2388 ();
 sg13g2_fill_2 FILLER_37_2424 ();
 sg13g2_fill_1 FILLER_37_2426 ();
 sg13g2_decap_4 FILLER_37_2498 ();
 sg13g2_fill_2 FILLER_37_2502 ();
 sg13g2_fill_1 FILLER_37_2544 ();
 sg13g2_fill_2 FILLER_37_2581 ();
 sg13g2_fill_1 FILLER_37_2583 ();
 sg13g2_decap_8 FILLER_37_2610 ();
 sg13g2_decap_4 FILLER_37_2617 ();
 sg13g2_decap_4 FILLER_37_2652 ();
 sg13g2_fill_1 FILLER_37_2656 ();
 sg13g2_decap_4 FILLER_38_30 ();
 sg13g2_fill_2 FILLER_38_43 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_169 ();
 sg13g2_fill_1 FILLER_38_171 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_416 ();
 sg13g2_fill_1 FILLER_38_418 ();
 sg13g2_fill_2 FILLER_38_443 ();
 sg13g2_fill_1 FILLER_38_445 ();
 sg13g2_fill_1 FILLER_38_455 ();
 sg13g2_fill_2 FILLER_38_508 ();
 sg13g2_decap_4 FILLER_38_574 ();
 sg13g2_decap_4 FILLER_38_604 ();
 sg13g2_fill_1 FILLER_38_608 ();
 sg13g2_decap_4 FILLER_38_615 ();
 sg13g2_fill_2 FILLER_38_619 ();
 sg13g2_fill_2 FILLER_38_657 ();
 sg13g2_fill_1 FILLER_38_668 ();
 sg13g2_decap_8 FILLER_38_678 ();
 sg13g2_fill_2 FILLER_38_685 ();
 sg13g2_fill_2 FILLER_38_700 ();
 sg13g2_fill_1 FILLER_38_702 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_fill_2 FILLER_38_714 ();
 sg13g2_fill_1 FILLER_38_716 ();
 sg13g2_fill_2 FILLER_38_722 ();
 sg13g2_fill_1 FILLER_38_754 ();
 sg13g2_fill_2 FILLER_38_806 ();
 sg13g2_fill_2 FILLER_38_835 ();
 sg13g2_fill_1 FILLER_38_837 ();
 sg13g2_decap_4 FILLER_38_876 ();
 sg13g2_fill_1 FILLER_38_880 ();
 sg13g2_decap_4 FILLER_38_915 ();
 sg13g2_fill_2 FILLER_38_919 ();
 sg13g2_fill_1 FILLER_38_927 ();
 sg13g2_fill_2 FILLER_38_1002 ();
 sg13g2_fill_1 FILLER_38_1004 ();
 sg13g2_fill_2 FILLER_38_1022 ();
 sg13g2_fill_2 FILLER_38_1042 ();
 sg13g2_fill_1 FILLER_38_1068 ();
 sg13g2_fill_2 FILLER_38_1083 ();
 sg13g2_fill_2 FILLER_38_1116 ();
 sg13g2_fill_2 FILLER_38_1129 ();
 sg13g2_fill_1 FILLER_38_1131 ();
 sg13g2_fill_2 FILLER_38_1137 ();
 sg13g2_fill_1 FILLER_38_1139 ();
 sg13g2_fill_2 FILLER_38_1151 ();
 sg13g2_fill_2 FILLER_38_1158 ();
 sg13g2_fill_1 FILLER_38_1181 ();
 sg13g2_fill_2 FILLER_38_1191 ();
 sg13g2_fill_1 FILLER_38_1193 ();
 sg13g2_decap_8 FILLER_38_1234 ();
 sg13g2_fill_2 FILLER_38_1342 ();
 sg13g2_fill_1 FILLER_38_1344 ();
 sg13g2_fill_2 FILLER_38_1418 ();
 sg13g2_fill_2 FILLER_38_1443 ();
 sg13g2_fill_2 FILLER_38_1479 ();
 sg13g2_fill_1 FILLER_38_1481 ();
 sg13g2_decap_4 FILLER_38_1540 ();
 sg13g2_fill_1 FILLER_38_1544 ();
 sg13g2_decap_4 FILLER_38_1580 ();
 sg13g2_fill_2 FILLER_38_1584 ();
 sg13g2_fill_2 FILLER_38_1612 ();
 sg13g2_fill_1 FILLER_38_1614 ();
 sg13g2_fill_2 FILLER_38_1645 ();
 sg13g2_fill_1 FILLER_38_1647 ();
 sg13g2_fill_1 FILLER_38_1693 ();
 sg13g2_decap_4 FILLER_38_1719 ();
 sg13g2_fill_2 FILLER_38_1754 ();
 sg13g2_fill_2 FILLER_38_1765 ();
 sg13g2_decap_4 FILLER_38_1771 ();
 sg13g2_fill_1 FILLER_38_1775 ();
 sg13g2_fill_2 FILLER_38_1791 ();
 sg13g2_fill_1 FILLER_38_1793 ();
 sg13g2_fill_2 FILLER_38_1806 ();
 sg13g2_fill_1 FILLER_38_1818 ();
 sg13g2_fill_2 FILLER_38_1870 ();
 sg13g2_decap_4 FILLER_38_1878 ();
 sg13g2_fill_2 FILLER_38_1922 ();
 sg13g2_fill_2 FILLER_38_1934 ();
 sg13g2_fill_2 FILLER_38_1974 ();
 sg13g2_fill_2 FILLER_38_2022 ();
 sg13g2_fill_2 FILLER_38_2065 ();
 sg13g2_fill_1 FILLER_38_2067 ();
 sg13g2_fill_2 FILLER_38_2077 ();
 sg13g2_decap_4 FILLER_38_2100 ();
 sg13g2_fill_1 FILLER_38_2104 ();
 sg13g2_fill_2 FILLER_38_2151 ();
 sg13g2_fill_1 FILLER_38_2153 ();
 sg13g2_fill_2 FILLER_38_2176 ();
 sg13g2_fill_1 FILLER_38_2178 ();
 sg13g2_decap_4 FILLER_38_2188 ();
 sg13g2_fill_1 FILLER_38_2192 ();
 sg13g2_fill_2 FILLER_38_2198 ();
 sg13g2_decap_8 FILLER_38_2204 ();
 sg13g2_fill_2 FILLER_38_2234 ();
 sg13g2_fill_1 FILLER_38_2236 ();
 sg13g2_fill_1 FILLER_38_2267 ();
 sg13g2_fill_2 FILLER_38_2323 ();
 sg13g2_fill_2 FILLER_38_2361 ();
 sg13g2_fill_2 FILLER_38_2399 ();
 sg13g2_fill_1 FILLER_38_2401 ();
 sg13g2_fill_2 FILLER_38_2436 ();
 sg13g2_fill_1 FILLER_38_2438 ();
 sg13g2_decap_4 FILLER_38_2465 ();
 sg13g2_fill_2 FILLER_38_2469 ();
 sg13g2_fill_1 FILLER_38_2503 ();
 sg13g2_decap_4 FILLER_38_2549 ();
 sg13g2_fill_2 FILLER_38_2570 ();
 sg13g2_fill_1 FILLER_38_2572 ();
 sg13g2_fill_2 FILLER_38_2592 ();
 sg13g2_decap_8 FILLER_38_2630 ();
 sg13g2_fill_1 FILLER_38_2647 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_fill_1 FILLER_39_66 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_fill_1 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_205 ();
 sg13g2_fill_2 FILLER_39_228 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_293 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_418 ();
 sg13g2_fill_2 FILLER_39_436 ();
 sg13g2_fill_1 FILLER_39_438 ();
 sg13g2_fill_2 FILLER_39_517 ();
 sg13g2_decap_4 FILLER_39_553 ();
 sg13g2_fill_2 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_576 ();
 sg13g2_decap_4 FILLER_39_583 ();
 sg13g2_fill_2 FILLER_39_587 ();
 sg13g2_decap_4 FILLER_39_593 ();
 sg13g2_fill_2 FILLER_39_597 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_fill_2 FILLER_39_623 ();
 sg13g2_fill_1 FILLER_39_625 ();
 sg13g2_decap_4 FILLER_39_631 ();
 sg13g2_fill_2 FILLER_39_657 ();
 sg13g2_fill_1 FILLER_39_659 ();
 sg13g2_fill_2 FILLER_39_728 ();
 sg13g2_fill_1 FILLER_39_730 ();
 sg13g2_fill_1 FILLER_39_779 ();
 sg13g2_fill_2 FILLER_39_846 ();
 sg13g2_fill_1 FILLER_39_848 ();
 sg13g2_decap_4 FILLER_39_857 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_fill_1 FILLER_39_875 ();
 sg13g2_fill_1 FILLER_39_931 ();
 sg13g2_fill_2 FILLER_39_937 ();
 sg13g2_fill_1 FILLER_39_939 ();
 sg13g2_fill_2 FILLER_39_974 ();
 sg13g2_fill_1 FILLER_39_985 ();
 sg13g2_fill_1 FILLER_39_1004 ();
 sg13g2_decap_4 FILLER_39_1010 ();
 sg13g2_decap_4 FILLER_39_1030 ();
 sg13g2_fill_1 FILLER_39_1034 ();
 sg13g2_fill_2 FILLER_39_1075 ();
 sg13g2_fill_1 FILLER_39_1111 ();
 sg13g2_fill_1 FILLER_39_1126 ();
 sg13g2_fill_2 FILLER_39_1153 ();
 sg13g2_fill_1 FILLER_39_1155 ();
 sg13g2_fill_1 FILLER_39_1165 ();
 sg13g2_fill_2 FILLER_39_1180 ();
 sg13g2_fill_1 FILLER_39_1182 ();
 sg13g2_decap_8 FILLER_39_1209 ();
 sg13g2_fill_2 FILLER_39_1216 ();
 sg13g2_fill_1 FILLER_39_1218 ();
 sg13g2_fill_1 FILLER_39_1223 ();
 sg13g2_decap_4 FILLER_39_1230 ();
 sg13g2_fill_2 FILLER_39_1272 ();
 sg13g2_fill_1 FILLER_39_1274 ();
 sg13g2_fill_1 FILLER_39_1283 ();
 sg13g2_fill_1 FILLER_39_1336 ();
 sg13g2_decap_4 FILLER_39_1363 ();
 sg13g2_fill_2 FILLER_39_1367 ();
 sg13g2_fill_1 FILLER_39_1389 ();
 sg13g2_decap_4 FILLER_39_1410 ();
 sg13g2_decap_4 FILLER_39_1424 ();
 sg13g2_fill_1 FILLER_39_1463 ();
 sg13g2_decap_4 FILLER_39_1498 ();
 sg13g2_fill_1 FILLER_39_1528 ();
 sg13g2_fill_1 FILLER_39_1532 ();
 sg13g2_decap_4 FILLER_39_1538 ();
 sg13g2_fill_1 FILLER_39_1546 ();
 sg13g2_decap_4 FILLER_39_1562 ();
 sg13g2_fill_1 FILLER_39_1566 ();
 sg13g2_decap_4 FILLER_39_1575 ();
 sg13g2_decap_4 FILLER_39_1593 ();
 sg13g2_decap_4 FILLER_39_1601 ();
 sg13g2_fill_1 FILLER_39_1605 ();
 sg13g2_fill_1 FILLER_39_1642 ();
 sg13g2_decap_4 FILLER_39_1674 ();
 sg13g2_fill_1 FILLER_39_1678 ();
 sg13g2_fill_1 FILLER_39_1705 ();
 sg13g2_fill_2 FILLER_39_1776 ();
 sg13g2_fill_1 FILLER_39_1778 ();
 sg13g2_fill_2 FILLER_39_1801 ();
 sg13g2_fill_2 FILLER_39_1843 ();
 sg13g2_fill_2 FILLER_39_1881 ();
 sg13g2_fill_1 FILLER_39_1883 ();
 sg13g2_fill_1 FILLER_39_1915 ();
 sg13g2_fill_2 FILLER_39_2019 ();
 sg13g2_fill_1 FILLER_39_2031 ();
 sg13g2_fill_2 FILLER_39_2094 ();
 sg13g2_fill_2 FILLER_39_2131 ();
 sg13g2_fill_2 FILLER_39_2143 ();
 sg13g2_fill_1 FILLER_39_2145 ();
 sg13g2_fill_1 FILLER_39_2172 ();
 sg13g2_decap_8 FILLER_39_2198 ();
 sg13g2_decap_4 FILLER_39_2205 ();
 sg13g2_fill_2 FILLER_39_2285 ();
 sg13g2_fill_1 FILLER_39_2287 ();
 sg13g2_fill_1 FILLER_39_2324 ();
 sg13g2_fill_1 FILLER_39_2382 ();
 sg13g2_fill_1 FILLER_39_2392 ();
 sg13g2_fill_2 FILLER_39_2411 ();
 sg13g2_fill_1 FILLER_39_2413 ();
 sg13g2_fill_2 FILLER_39_2430 ();
 sg13g2_fill_1 FILLER_39_2432 ();
 sg13g2_fill_2 FILLER_39_2457 ();
 sg13g2_fill_2 FILLER_39_2490 ();
 sg13g2_fill_2 FILLER_39_2554 ();
 sg13g2_fill_1 FILLER_39_2556 ();
 sg13g2_fill_2 FILLER_39_2607 ();
 sg13g2_fill_1 FILLER_39_2609 ();
 sg13g2_fill_2 FILLER_39_2623 ();
 sg13g2_fill_2 FILLER_39_2640 ();
 sg13g2_fill_1 FILLER_39_2642 ();
 sg13g2_fill_1 FILLER_39_2673 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_fill_2 FILLER_40_9 ();
 sg13g2_decap_4 FILLER_40_15 ();
 sg13g2_fill_2 FILLER_40_19 ();
 sg13g2_decap_4 FILLER_40_145 ();
 sg13g2_fill_2 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_decap_4 FILLER_40_304 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_399 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_412 ();
 sg13g2_fill_2 FILLER_40_445 ();
 sg13g2_fill_1 FILLER_40_479 ();
 sg13g2_fill_2 FILLER_40_485 ();
 sg13g2_fill_1 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_496 ();
 sg13g2_fill_2 FILLER_40_502 ();
 sg13g2_fill_1 FILLER_40_504 ();
 sg13g2_fill_1 FILLER_40_529 ();
 sg13g2_fill_2 FILLER_40_575 ();
 sg13g2_fill_2 FILLER_40_608 ();
 sg13g2_fill_1 FILLER_40_610 ();
 sg13g2_fill_2 FILLER_40_628 ();
 sg13g2_fill_2 FILLER_40_643 ();
 sg13g2_fill_1 FILLER_40_645 ();
 sg13g2_decap_8 FILLER_40_656 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_fill_2 FILLER_40_684 ();
 sg13g2_fill_2 FILLER_40_696 ();
 sg13g2_fill_2 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_fill_2 FILLER_40_776 ();
 sg13g2_fill_2 FILLER_40_791 ();
 sg13g2_fill_2 FILLER_40_887 ();
 sg13g2_fill_1 FILLER_40_910 ();
 sg13g2_fill_1 FILLER_40_929 ();
 sg13g2_fill_2 FILLER_40_961 ();
 sg13g2_fill_1 FILLER_40_978 ();
 sg13g2_fill_1 FILLER_40_1025 ();
 sg13g2_fill_2 FILLER_40_1040 ();
 sg13g2_fill_1 FILLER_40_1060 ();
 sg13g2_fill_2 FILLER_40_1092 ();
 sg13g2_fill_2 FILLER_40_1175 ();
 sg13g2_fill_1 FILLER_40_1177 ();
 sg13g2_fill_1 FILLER_40_1199 ();
 sg13g2_decap_4 FILLER_40_1217 ();
 sg13g2_fill_1 FILLER_40_1221 ();
 sg13g2_fill_1 FILLER_40_1356 ();
 sg13g2_decap_4 FILLER_40_1377 ();
 sg13g2_fill_1 FILLER_40_1381 ();
 sg13g2_fill_2 FILLER_40_1385 ();
 sg13g2_fill_1 FILLER_40_1397 ();
 sg13g2_fill_1 FILLER_40_1403 ();
 sg13g2_decap_4 FILLER_40_1409 ();
 sg13g2_fill_2 FILLER_40_1466 ();
 sg13g2_fill_1 FILLER_40_1477 ();
 sg13g2_fill_2 FILLER_40_1482 ();
 sg13g2_fill_1 FILLER_40_1484 ();
 sg13g2_decap_4 FILLER_40_1493 ();
 sg13g2_fill_1 FILLER_40_1497 ();
 sg13g2_fill_2 FILLER_40_1529 ();
 sg13g2_fill_1 FILLER_40_1582 ();
 sg13g2_decap_8 FILLER_40_1609 ();
 sg13g2_fill_2 FILLER_40_1620 ();
 sg13g2_fill_1 FILLER_40_1737 ();
 sg13g2_decap_4 FILLER_40_1768 ();
 sg13g2_fill_1 FILLER_40_1798 ();
 sg13g2_decap_8 FILLER_40_1803 ();
 sg13g2_fill_2 FILLER_40_1810 ();
 sg13g2_decap_4 FILLER_40_1825 ();
 sg13g2_fill_1 FILLER_40_1829 ();
 sg13g2_fill_2 FILLER_40_1849 ();
 sg13g2_fill_2 FILLER_40_1874 ();
 sg13g2_fill_2 FILLER_40_1899 ();
 sg13g2_fill_1 FILLER_40_1901 ();
 sg13g2_decap_8 FILLER_40_1936 ();
 sg13g2_fill_1 FILLER_40_1943 ();
 sg13g2_fill_1 FILLER_40_1961 ();
 sg13g2_decap_4 FILLER_40_2024 ();
 sg13g2_fill_1 FILLER_40_2028 ();
 sg13g2_fill_1 FILLER_40_2055 ();
 sg13g2_fill_2 FILLER_40_2087 ();
 sg13g2_fill_1 FILLER_40_2089 ();
 sg13g2_fill_1 FILLER_40_2165 ();
 sg13g2_fill_2 FILLER_40_2241 ();
 sg13g2_fill_1 FILLER_40_2243 ();
 sg13g2_fill_1 FILLER_40_2263 ();
 sg13g2_fill_1 FILLER_40_2290 ();
 sg13g2_decap_4 FILLER_40_2321 ();
 sg13g2_fill_2 FILLER_40_2325 ();
 sg13g2_fill_1 FILLER_40_2341 ();
 sg13g2_fill_1 FILLER_40_2378 ();
 sg13g2_fill_1 FILLER_40_2383 ();
 sg13g2_decap_4 FILLER_40_2430 ();
 sg13g2_fill_2 FILLER_40_2434 ();
 sg13g2_decap_4 FILLER_40_2471 ();
 sg13g2_fill_2 FILLER_40_2475 ();
 sg13g2_fill_2 FILLER_40_2515 ();
 sg13g2_fill_2 FILLER_40_2557 ();
 sg13g2_fill_1 FILLER_40_2559 ();
 sg13g2_fill_1 FILLER_40_2578 ();
 sg13g2_decap_8 FILLER_40_2626 ();
 sg13g2_fill_2 FILLER_40_2633 ();
 sg13g2_fill_1 FILLER_40_2635 ();
 sg13g2_fill_2 FILLER_40_2646 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_fill_2 FILLER_41_136 ();
 sg13g2_decap_8 FILLER_41_144 ();
 sg13g2_fill_2 FILLER_41_151 ();
 sg13g2_fill_2 FILLER_41_158 ();
 sg13g2_fill_2 FILLER_41_168 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_fill_2 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_246 ();
 sg13g2_decap_4 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_2 FILLER_41_313 ();
 sg13g2_fill_1 FILLER_41_315 ();
 sg13g2_fill_2 FILLER_41_342 ();
 sg13g2_fill_2 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_fill_2 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_421 ();
 sg13g2_fill_1 FILLER_41_427 ();
 sg13g2_fill_1 FILLER_41_453 ();
 sg13g2_fill_2 FILLER_41_459 ();
 sg13g2_fill_2 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_fill_1 FILLER_41_531 ();
 sg13g2_decap_4 FILLER_41_547 ();
 sg13g2_fill_2 FILLER_41_555 ();
 sg13g2_fill_2 FILLER_41_566 ();
 sg13g2_decap_4 FILLER_41_576 ();
 sg13g2_decap_8 FILLER_41_592 ();
 sg13g2_decap_4 FILLER_41_599 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_693 ();
 sg13g2_fill_2 FILLER_41_714 ();
 sg13g2_decap_4 FILLER_41_724 ();
 sg13g2_fill_2 FILLER_41_762 ();
 sg13g2_fill_2 FILLER_41_833 ();
 sg13g2_fill_1 FILLER_41_835 ();
 sg13g2_fill_2 FILLER_41_855 ();
 sg13g2_fill_2 FILLER_41_871 ();
 sg13g2_fill_2 FILLER_41_917 ();
 sg13g2_fill_1 FILLER_41_919 ();
 sg13g2_fill_2 FILLER_41_940 ();
 sg13g2_fill_2 FILLER_41_950 ();
 sg13g2_fill_1 FILLER_41_972 ();
 sg13g2_fill_2 FILLER_41_982 ();
 sg13g2_fill_1 FILLER_41_984 ();
 sg13g2_fill_2 FILLER_41_999 ();
 sg13g2_fill_2 FILLER_41_1015 ();
 sg13g2_fill_1 FILLER_41_1017 ();
 sg13g2_fill_2 FILLER_41_1074 ();
 sg13g2_fill_1 FILLER_41_1076 ();
 sg13g2_fill_2 FILLER_41_1126 ();
 sg13g2_fill_1 FILLER_41_1159 ();
 sg13g2_decap_4 FILLER_41_1198 ();
 sg13g2_fill_2 FILLER_41_1202 ();
 sg13g2_fill_1 FILLER_41_1234 ();
 sg13g2_fill_2 FILLER_41_1241 ();
 sg13g2_fill_1 FILLER_41_1243 ();
 sg13g2_fill_2 FILLER_41_1312 ();
 sg13g2_fill_2 FILLER_41_1327 ();
 sg13g2_fill_2 FILLER_41_1444 ();
 sg13g2_fill_1 FILLER_41_1472 ();
 sg13g2_fill_2 FILLER_41_1547 ();
 sg13g2_fill_2 FILLER_41_1566 ();
 sg13g2_fill_2 FILLER_41_1574 ();
 sg13g2_fill_1 FILLER_41_1576 ();
 sg13g2_fill_2 FILLER_41_1591 ();
 sg13g2_fill_1 FILLER_41_1593 ();
 sg13g2_fill_1 FILLER_41_1598 ();
 sg13g2_decap_4 FILLER_41_1642 ();
 sg13g2_fill_2 FILLER_41_1672 ();
 sg13g2_fill_1 FILLER_41_1674 ();
 sg13g2_fill_2 FILLER_41_1701 ();
 sg13g2_fill_2 FILLER_41_1757 ();
 sg13g2_fill_1 FILLER_41_1759 ();
 sg13g2_fill_1 FILLER_41_1786 ();
 sg13g2_fill_1 FILLER_41_1807 ();
 sg13g2_decap_8 FILLER_41_2015 ();
 sg13g2_fill_1 FILLER_41_2022 ();
 sg13g2_fill_1 FILLER_41_2053 ();
 sg13g2_fill_2 FILLER_41_2068 ();
 sg13g2_fill_2 FILLER_41_2093 ();
 sg13g2_fill_1 FILLER_41_2095 ();
 sg13g2_fill_2 FILLER_41_2122 ();
 sg13g2_fill_1 FILLER_41_2124 ();
 sg13g2_fill_2 FILLER_41_2138 ();
 sg13g2_fill_2 FILLER_41_2149 ();
 sg13g2_fill_1 FILLER_41_2151 ();
 sg13g2_fill_1 FILLER_41_2274 ();
 sg13g2_decap_4 FILLER_41_2322 ();
 sg13g2_fill_2 FILLER_41_2336 ();
 sg13g2_fill_2 FILLER_41_2365 ();
 sg13g2_fill_1 FILLER_41_2367 ();
 sg13g2_fill_1 FILLER_41_2423 ();
 sg13g2_decap_8 FILLER_41_2430 ();
 sg13g2_fill_1 FILLER_41_2437 ();
 sg13g2_fill_1 FILLER_41_2451 ();
 sg13g2_fill_2 FILLER_41_2488 ();
 sg13g2_fill_2 FILLER_41_2526 ();
 sg13g2_fill_2 FILLER_41_2532 ();
 sg13g2_fill_2 FILLER_41_2544 ();
 sg13g2_fill_1 FILLER_41_2598 ();
 sg13g2_fill_1 FILLER_41_2608 ();
 sg13g2_fill_2 FILLER_41_2671 ();
 sg13g2_fill_1 FILLER_41_2673 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_11 ();
 sg13g2_decap_4 FILLER_42_16 ();
 sg13g2_fill_1 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_116 ();
 sg13g2_decap_4 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_fill_2 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_207 ();
 sg13g2_fill_1 FILLER_42_216 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_fill_2 FILLER_42_297 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_335 ();
 sg13g2_fill_2 FILLER_42_367 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_fill_2 FILLER_42_390 ();
 sg13g2_fill_2 FILLER_42_444 ();
 sg13g2_fill_2 FILLER_42_476 ();
 sg13g2_fill_1 FILLER_42_478 ();
 sg13g2_fill_1 FILLER_42_500 ();
 sg13g2_fill_2 FILLER_42_520 ();
 sg13g2_fill_1 FILLER_42_522 ();
 sg13g2_fill_2 FILLER_42_527 ();
 sg13g2_fill_1 FILLER_42_529 ();
 sg13g2_fill_2 FILLER_42_566 ();
 sg13g2_fill_1 FILLER_42_568 ();
 sg13g2_decap_4 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_621 ();
 sg13g2_decap_4 FILLER_42_628 ();
 sg13g2_fill_2 FILLER_42_632 ();
 sg13g2_decap_4 FILLER_42_662 ();
 sg13g2_fill_1 FILLER_42_690 ();
 sg13g2_fill_2 FILLER_42_697 ();
 sg13g2_decap_4 FILLER_42_718 ();
 sg13g2_fill_2 FILLER_42_730 ();
 sg13g2_fill_1 FILLER_42_740 ();
 sg13g2_decap_8 FILLER_42_751 ();
 sg13g2_decap_4 FILLER_42_758 ();
 sg13g2_fill_1 FILLER_42_762 ();
 sg13g2_fill_1 FILLER_42_773 ();
 sg13g2_fill_2 FILLER_42_818 ();
 sg13g2_fill_2 FILLER_42_865 ();
 sg13g2_fill_1 FILLER_42_867 ();
 sg13g2_fill_1 FILLER_42_899 ();
 sg13g2_fill_2 FILLER_42_961 ();
 sg13g2_fill_1 FILLER_42_963 ();
 sg13g2_fill_2 FILLER_42_974 ();
 sg13g2_decap_4 FILLER_42_990 ();
 sg13g2_decap_4 FILLER_42_1010 ();
 sg13g2_fill_2 FILLER_42_1040 ();
 sg13g2_fill_2 FILLER_42_1055 ();
 sg13g2_fill_1 FILLER_42_1057 ();
 sg13g2_fill_2 FILLER_42_1067 ();
 sg13g2_fill_1 FILLER_42_1069 ();
 sg13g2_fill_2 FILLER_42_1096 ();
 sg13g2_fill_1 FILLER_42_1108 ();
 sg13g2_fill_2 FILLER_42_1141 ();
 sg13g2_fill_2 FILLER_42_1169 ();
 sg13g2_fill_1 FILLER_42_1171 ();
 sg13g2_fill_2 FILLER_42_1177 ();
 sg13g2_fill_1 FILLER_42_1213 ();
 sg13g2_fill_2 FILLER_42_1289 ();
 sg13g2_fill_2 FILLER_42_1298 ();
 sg13g2_fill_1 FILLER_42_1336 ();
 sg13g2_decap_4 FILLER_42_1380 ();
 sg13g2_fill_1 FILLER_42_1384 ();
 sg13g2_fill_1 FILLER_42_1393 ();
 sg13g2_decap_4 FILLER_42_1404 ();
 sg13g2_fill_1 FILLER_42_1408 ();
 sg13g2_fill_1 FILLER_42_1414 ();
 sg13g2_fill_2 FILLER_42_1439 ();
 sg13g2_fill_1 FILLER_42_1441 ();
 sg13g2_fill_1 FILLER_42_1460 ();
 sg13g2_fill_1 FILLER_42_1555 ();
 sg13g2_fill_2 FILLER_42_1607 ();
 sg13g2_fill_1 FILLER_42_1641 ();
 sg13g2_fill_1 FILLER_42_1652 ();
 sg13g2_fill_2 FILLER_42_1696 ();
 sg13g2_fill_1 FILLER_42_1698 ();
 sg13g2_fill_2 FILLER_42_1736 ();
 sg13g2_fill_1 FILLER_42_1738 ();
 sg13g2_fill_1 FILLER_42_1769 ();
 sg13g2_decap_4 FILLER_42_1774 ();
 sg13g2_fill_2 FILLER_42_1835 ();
 sg13g2_fill_2 FILLER_42_1867 ();
 sg13g2_fill_1 FILLER_42_1869 ();
 sg13g2_decap_8 FILLER_42_1878 ();
 sg13g2_fill_1 FILLER_42_1885 ();
 sg13g2_fill_1 FILLER_42_1896 ();
 sg13g2_fill_1 FILLER_42_1907 ();
 sg13g2_fill_1 FILLER_42_1957 ();
 sg13g2_fill_2 FILLER_42_1968 ();
 sg13g2_fill_2 FILLER_42_2010 ();
 sg13g2_decap_8 FILLER_42_2038 ();
 sg13g2_fill_2 FILLER_42_2081 ();
 sg13g2_fill_1 FILLER_42_2083 ();
 sg13g2_fill_2 FILLER_42_2114 ();
 sg13g2_fill_1 FILLER_42_2116 ();
 sg13g2_fill_1 FILLER_42_2161 ();
 sg13g2_decap_4 FILLER_42_2208 ();
 sg13g2_fill_2 FILLER_42_2216 ();
 sg13g2_fill_2 FILLER_42_2226 ();
 sg13g2_fill_1 FILLER_42_2228 ();
 sg13g2_fill_2 FILLER_42_2248 ();
 sg13g2_decap_4 FILLER_42_2369 ();
 sg13g2_fill_1 FILLER_42_2373 ();
 sg13g2_fill_1 FILLER_42_2414 ();
 sg13g2_fill_1 FILLER_42_2469 ();
 sg13g2_fill_2 FILLER_42_2491 ();
 sg13g2_fill_2 FILLER_42_2506 ();
 sg13g2_fill_1 FILLER_42_2588 ();
 sg13g2_decap_4 FILLER_42_2668 ();
 sg13g2_fill_2 FILLER_42_2672 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_75 ();
 sg13g2_fill_1 FILLER_43_86 ();
 sg13g2_decap_4 FILLER_43_110 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_1 FILLER_43_127 ();
 sg13g2_decap_4 FILLER_43_141 ();
 sg13g2_decap_4 FILLER_43_159 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_280 ();
 sg13g2_fill_1 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_375 ();
 sg13g2_fill_1 FILLER_43_444 ();
 sg13g2_fill_2 FILLER_43_458 ();
 sg13g2_fill_1 FILLER_43_460 ();
 sg13g2_fill_2 FILLER_43_494 ();
 sg13g2_fill_2 FILLER_43_505 ();
 sg13g2_fill_1 FILLER_43_538 ();
 sg13g2_fill_1 FILLER_43_548 ();
 sg13g2_decap_8 FILLER_43_570 ();
 sg13g2_fill_1 FILLER_43_577 ();
 sg13g2_fill_2 FILLER_43_592 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_fill_2 FILLER_43_620 ();
 sg13g2_decap_4 FILLER_43_649 ();
 sg13g2_decap_4 FILLER_43_664 ();
 sg13g2_fill_1 FILLER_43_694 ();
 sg13g2_fill_2 FILLER_43_709 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_731 ();
 sg13g2_decap_4 FILLER_43_737 ();
 sg13g2_decap_8 FILLER_43_751 ();
 sg13g2_fill_1 FILLER_43_789 ();
 sg13g2_fill_2 FILLER_43_805 ();
 sg13g2_fill_1 FILLER_43_831 ();
 sg13g2_fill_2 FILLER_43_867 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_fill_2 FILLER_43_917 ();
 sg13g2_fill_2 FILLER_43_923 ();
 sg13g2_decap_4 FILLER_43_935 ();
 sg13g2_fill_2 FILLER_43_975 ();
 sg13g2_fill_2 FILLER_43_985 ();
 sg13g2_fill_1 FILLER_43_987 ();
 sg13g2_fill_2 FILLER_43_1019 ();
 sg13g2_fill_1 FILLER_43_1034 ();
 sg13g2_fill_1 FILLER_43_1078 ();
 sg13g2_fill_1 FILLER_43_1104 ();
 sg13g2_decap_4 FILLER_43_1115 ();
 sg13g2_fill_1 FILLER_43_1119 ();
 sg13g2_fill_1 FILLER_43_1135 ();
 sg13g2_fill_1 FILLER_43_1149 ();
 sg13g2_fill_1 FILLER_43_1160 ();
 sg13g2_decap_4 FILLER_43_1202 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_fill_2 FILLER_43_1277 ();
 sg13g2_fill_2 FILLER_43_1287 ();
 sg13g2_fill_1 FILLER_43_1328 ();
 sg13g2_decap_4 FILLER_43_1334 ();
 sg13g2_fill_1 FILLER_43_1352 ();
 sg13g2_fill_1 FILLER_43_1362 ();
 sg13g2_fill_2 FILLER_43_1398 ();
 sg13g2_fill_2 FILLER_43_1522 ();
 sg13g2_fill_2 FILLER_43_1568 ();
 sg13g2_fill_1 FILLER_43_1570 ();
 sg13g2_fill_2 FILLER_43_1606 ();
 sg13g2_decap_4 FILLER_43_1634 ();
 sg13g2_fill_2 FILLER_43_1638 ();
 sg13g2_decap_8 FILLER_43_1666 ();
 sg13g2_fill_2 FILLER_43_1768 ();
 sg13g2_fill_2 FILLER_43_1806 ();
 sg13g2_decap_4 FILLER_43_1844 ();
 sg13g2_fill_2 FILLER_43_1848 ();
 sg13g2_decap_4 FILLER_43_1886 ();
 sg13g2_fill_1 FILLER_43_1959 ();
 sg13g2_fill_2 FILLER_43_1975 ();
 sg13g2_fill_2 FILLER_43_1995 ();
 sg13g2_fill_2 FILLER_43_2054 ();
 sg13g2_fill_1 FILLER_43_2070 ();
 sg13g2_fill_1 FILLER_43_2108 ();
 sg13g2_decap_4 FILLER_43_2139 ();
 sg13g2_fill_2 FILLER_43_2175 ();
 sg13g2_fill_1 FILLER_43_2177 ();
 sg13g2_fill_1 FILLER_43_2237 ();
 sg13g2_fill_1 FILLER_43_2270 ();
 sg13g2_fill_2 FILLER_43_2284 ();
 sg13g2_fill_1 FILLER_43_2286 ();
 sg13g2_fill_1 FILLER_43_2313 ();
 sg13g2_fill_2 FILLER_43_2323 ();
 sg13g2_fill_1 FILLER_43_2325 ();
 sg13g2_decap_4 FILLER_43_2344 ();
 sg13g2_fill_1 FILLER_43_2388 ();
 sg13g2_fill_1 FILLER_43_2399 ();
 sg13g2_fill_2 FILLER_43_2442 ();
 sg13g2_fill_2 FILLER_43_2510 ();
 sg13g2_fill_1 FILLER_43_2512 ();
 sg13g2_fill_2 FILLER_43_2534 ();
 sg13g2_fill_2 FILLER_43_2581 ();
 sg13g2_fill_1 FILLER_43_2583 ();
 sg13g2_fill_2 FILLER_43_2619 ();
 sg13g2_fill_1 FILLER_43_2621 ();
 sg13g2_decap_8 FILLER_43_2658 ();
 sg13g2_decap_8 FILLER_43_2665 ();
 sg13g2_fill_2 FILLER_43_2672 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_fill_1 FILLER_44_29 ();
 sg13g2_decap_8 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_99 ();
 sg13g2_fill_2 FILLER_44_109 ();
 sg13g2_fill_1 FILLER_44_111 ();
 sg13g2_fill_1 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_131 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_152 ();
 sg13g2_fill_1 FILLER_44_172 ();
 sg13g2_decap_4 FILLER_44_178 ();
 sg13g2_fill_1 FILLER_44_182 ();
 sg13g2_fill_2 FILLER_44_189 ();
 sg13g2_fill_1 FILLER_44_191 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_231 ();
 sg13g2_fill_1 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_261 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_305 ();
 sg13g2_fill_1 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_344 ();
 sg13g2_fill_2 FILLER_44_364 ();
 sg13g2_fill_2 FILLER_44_396 ();
 sg13g2_fill_1 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_413 ();
 sg13g2_fill_2 FILLER_44_431 ();
 sg13g2_fill_1 FILLER_44_442 ();
 sg13g2_fill_2 FILLER_44_457 ();
 sg13g2_fill_1 FILLER_44_478 ();
 sg13g2_fill_2 FILLER_44_516 ();
 sg13g2_decap_4 FILLER_44_602 ();
 sg13g2_fill_2 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_618 ();
 sg13g2_fill_1 FILLER_44_625 ();
 sg13g2_fill_2 FILLER_44_646 ();
 sg13g2_fill_1 FILLER_44_652 ();
 sg13g2_fill_1 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_664 ();
 sg13g2_fill_2 FILLER_44_671 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_691 ();
 sg13g2_decap_4 FILLER_44_698 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_fill_1 FILLER_44_774 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_fill_2 FILLER_44_892 ();
 sg13g2_fill_1 FILLER_44_894 ();
 sg13g2_fill_2 FILLER_44_947 ();
 sg13g2_fill_1 FILLER_44_949 ();
 sg13g2_decap_4 FILLER_44_984 ();
 sg13g2_fill_2 FILLER_44_988 ();
 sg13g2_fill_2 FILLER_44_1007 ();
 sg13g2_fill_1 FILLER_44_1009 ();
 sg13g2_decap_4 FILLER_44_1021 ();
 sg13g2_fill_2 FILLER_44_1025 ();
 sg13g2_fill_2 FILLER_44_1031 ();
 sg13g2_fill_1 FILLER_44_1044 ();
 sg13g2_fill_1 FILLER_44_1065 ();
 sg13g2_fill_2 FILLER_44_1076 ();
 sg13g2_fill_1 FILLER_44_1083 ();
 sg13g2_fill_2 FILLER_44_1154 ();
 sg13g2_fill_1 FILLER_44_1156 ();
 sg13g2_fill_2 FILLER_44_1162 ();
 sg13g2_fill_1 FILLER_44_1178 ();
 sg13g2_fill_1 FILLER_44_1200 ();
 sg13g2_fill_1 FILLER_44_1234 ();
 sg13g2_fill_2 FILLER_44_1245 ();
 sg13g2_fill_1 FILLER_44_1288 ();
 sg13g2_fill_1 FILLER_44_1304 ();
 sg13g2_fill_1 FILLER_44_1323 ();
 sg13g2_decap_4 FILLER_44_1368 ();
 sg13g2_fill_2 FILLER_44_1377 ();
 sg13g2_fill_1 FILLER_44_1379 ();
 sg13g2_decap_8 FILLER_44_1383 ();
 sg13g2_decap_8 FILLER_44_1390 ();
 sg13g2_fill_2 FILLER_44_1400 ();
 sg13g2_fill_2 FILLER_44_1407 ();
 sg13g2_fill_1 FILLER_44_1446 ();
 sg13g2_fill_2 FILLER_44_1451 ();
 sg13g2_fill_1 FILLER_44_1453 ();
 sg13g2_decap_4 FILLER_44_1466 ();
 sg13g2_fill_1 FILLER_44_1470 ();
 sg13g2_fill_2 FILLER_44_1491 ();
 sg13g2_fill_1 FILLER_44_1493 ();
 sg13g2_fill_1 FILLER_44_1499 ();
 sg13g2_fill_2 FILLER_44_1507 ();
 sg13g2_fill_1 FILLER_44_1509 ();
 sg13g2_fill_2 FILLER_44_1531 ();
 sg13g2_fill_1 FILLER_44_1580 ();
 sg13g2_decap_4 FILLER_44_1664 ();
 sg13g2_fill_1 FILLER_44_1678 ();
 sg13g2_fill_2 FILLER_44_1702 ();
 sg13g2_fill_1 FILLER_44_1704 ();
 sg13g2_fill_2 FILLER_44_1851 ();
 sg13g2_fill_1 FILLER_44_1853 ();
 sg13g2_fill_1 FILLER_44_1872 ();
 sg13g2_fill_2 FILLER_44_1888 ();
 sg13g2_fill_1 FILLER_44_1905 ();
 sg13g2_fill_1 FILLER_44_1946 ();
 sg13g2_fill_2 FILLER_44_1973 ();
 sg13g2_fill_2 FILLER_44_2010 ();
 sg13g2_decap_4 FILLER_44_2039 ();
 sg13g2_fill_2 FILLER_44_2043 ();
 sg13g2_fill_2 FILLER_44_2081 ();
 sg13g2_fill_1 FILLER_44_2083 ();
 sg13g2_fill_2 FILLER_44_2119 ();
 sg13g2_decap_4 FILLER_44_2294 ();
 sg13g2_fill_2 FILLER_44_2298 ();
 sg13g2_fill_2 FILLER_44_2367 ();
 sg13g2_fill_2 FILLER_44_2388 ();
 sg13g2_fill_2 FILLER_44_2435 ();
 sg13g2_fill_1 FILLER_44_2437 ();
 sg13g2_decap_4 FILLER_44_2457 ();
 sg13g2_decap_8 FILLER_44_2469 ();
 sg13g2_fill_1 FILLER_44_2476 ();
 sg13g2_fill_2 FILLER_44_2487 ();
 sg13g2_fill_1 FILLER_44_2489 ();
 sg13g2_fill_2 FILLER_44_2503 ();
 sg13g2_decap_4 FILLER_44_2546 ();
 sg13g2_fill_2 FILLER_44_2576 ();
 sg13g2_fill_1 FILLER_44_2578 ();
 sg13g2_fill_2 FILLER_44_2589 ();
 sg13g2_fill_1 FILLER_44_2609 ();
 sg13g2_decap_8 FILLER_44_2659 ();
 sg13g2_decap_8 FILLER_44_2666 ();
 sg13g2_fill_1 FILLER_44_2673 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_59 ();
 sg13g2_fill_2 FILLER_45_65 ();
 sg13g2_decap_4 FILLER_45_84 ();
 sg13g2_fill_1 FILLER_45_88 ();
 sg13g2_fill_1 FILLER_45_101 ();
 sg13g2_decap_4 FILLER_45_116 ();
 sg13g2_fill_1 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_fill_1 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_174 ();
 sg13g2_fill_2 FILLER_45_191 ();
 sg13g2_fill_1 FILLER_45_193 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_fill_2 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_2 FILLER_45_440 ();
 sg13g2_fill_1 FILLER_45_442 ();
 sg13g2_fill_1 FILLER_45_486 ();
 sg13g2_fill_2 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_508 ();
 sg13g2_fill_1 FILLER_45_560 ();
 sg13g2_decap_4 FILLER_45_565 ();
 sg13g2_fill_2 FILLER_45_573 ();
 sg13g2_fill_1 FILLER_45_575 ();
 sg13g2_decap_8 FILLER_45_589 ();
 sg13g2_fill_1 FILLER_45_621 ();
 sg13g2_decap_8 FILLER_45_628 ();
 sg13g2_decap_4 FILLER_45_635 ();
 sg13g2_fill_1 FILLER_45_639 ();
 sg13g2_fill_1 FILLER_45_655 ();
 sg13g2_decap_4 FILLER_45_667 ();
 sg13g2_fill_1 FILLER_45_671 ();
 sg13g2_fill_2 FILLER_45_690 ();
 sg13g2_fill_1 FILLER_45_692 ();
 sg13g2_fill_2 FILLER_45_701 ();
 sg13g2_fill_2 FILLER_45_720 ();
 sg13g2_decap_8 FILLER_45_737 ();
 sg13g2_fill_1 FILLER_45_744 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_786 ();
 sg13g2_fill_1 FILLER_45_835 ();
 sg13g2_fill_2 FILLER_45_863 ();
 sg13g2_fill_1 FILLER_45_878 ();
 sg13g2_decap_4 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_918 ();
 sg13g2_fill_1 FILLER_45_941 ();
 sg13g2_decap_4 FILLER_45_1099 ();
 sg13g2_fill_1 FILLER_45_1142 ();
 sg13g2_fill_1 FILLER_45_1148 ();
 sg13g2_fill_2 FILLER_45_1201 ();
 sg13g2_fill_1 FILLER_45_1203 ();
 sg13g2_fill_2 FILLER_45_1256 ();
 sg13g2_fill_1 FILLER_45_1279 ();
 sg13g2_fill_2 FILLER_45_1315 ();
 sg13g2_fill_1 FILLER_45_1317 ();
 sg13g2_fill_2 FILLER_45_1332 ();
 sg13g2_fill_1 FILLER_45_1347 ();
 sg13g2_fill_2 FILLER_45_1397 ();
 sg13g2_fill_1 FILLER_45_1422 ();
 sg13g2_fill_2 FILLER_45_1442 ();
 sg13g2_fill_1 FILLER_45_1444 ();
 sg13g2_fill_2 FILLER_45_1449 ();
 sg13g2_fill_1 FILLER_45_1451 ();
 sg13g2_decap_8 FILLER_45_1456 ();
 sg13g2_fill_1 FILLER_45_1503 ();
 sg13g2_fill_2 FILLER_45_1568 ();
 sg13g2_fill_2 FILLER_45_1615 ();
 sg13g2_decap_4 FILLER_45_1639 ();
 sg13g2_fill_2 FILLER_45_1643 ();
 sg13g2_fill_2 FILLER_45_1705 ();
 sg13g2_fill_1 FILLER_45_1707 ();
 sg13g2_fill_2 FILLER_45_1760 ();
 sg13g2_fill_1 FILLER_45_1762 ();
 sg13g2_decap_4 FILLER_45_1771 ();
 sg13g2_fill_1 FILLER_45_1842 ();
 sg13g2_fill_2 FILLER_45_1869 ();
 sg13g2_fill_1 FILLER_45_1871 ();
 sg13g2_fill_2 FILLER_45_1910 ();
 sg13g2_fill_1 FILLER_45_1912 ();
 sg13g2_fill_1 FILLER_45_1923 ();
 sg13g2_fill_1 FILLER_45_1950 ();
 sg13g2_fill_2 FILLER_45_1959 ();
 sg13g2_fill_2 FILLER_45_1978 ();
 sg13g2_fill_2 FILLER_45_1989 ();
 sg13g2_fill_1 FILLER_45_2016 ();
 sg13g2_fill_2 FILLER_45_2059 ();
 sg13g2_fill_2 FILLER_45_2074 ();
 sg13g2_fill_1 FILLER_45_2089 ();
 sg13g2_fill_1 FILLER_45_2112 ();
 sg13g2_fill_2 FILLER_45_2141 ();
 sg13g2_fill_1 FILLER_45_2156 ();
 sg13g2_fill_1 FILLER_45_2177 ();
 sg13g2_fill_2 FILLER_45_2186 ();
 sg13g2_fill_1 FILLER_45_2207 ();
 sg13g2_fill_1 FILLER_45_2235 ();
 sg13g2_fill_1 FILLER_45_2266 ();
 sg13g2_fill_2 FILLER_45_2279 ();
 sg13g2_fill_1 FILLER_45_2281 ();
 sg13g2_fill_1 FILLER_45_2323 ();
 sg13g2_fill_2 FILLER_45_2330 ();
 sg13g2_fill_1 FILLER_45_2332 ();
 sg13g2_fill_2 FILLER_45_2477 ();
 sg13g2_fill_1 FILLER_45_2479 ();
 sg13g2_fill_2 FILLER_45_2506 ();
 sg13g2_fill_1 FILLER_45_2508 ();
 sg13g2_fill_1 FILLER_45_2549 ();
 sg13g2_decap_8 FILLER_45_2651 ();
 sg13g2_decap_8 FILLER_45_2658 ();
 sg13g2_decap_8 FILLER_45_2665 ();
 sg13g2_fill_2 FILLER_45_2672 ();
 sg13g2_fill_2 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_74 ();
 sg13g2_decap_4 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_92 ();
 sg13g2_decap_4 FILLER_46_104 ();
 sg13g2_fill_1 FILLER_46_108 ();
 sg13g2_decap_4 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_2 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_163 ();
 sg13g2_decap_8 FILLER_46_183 ();
 sg13g2_fill_2 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_234 ();
 sg13g2_fill_1 FILLER_46_236 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_decap_4 FILLER_46_278 ();
 sg13g2_fill_1 FILLER_46_299 ();
 sg13g2_fill_2 FILLER_46_317 ();
 sg13g2_fill_1 FILLER_46_328 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_384 ();
 sg13g2_fill_2 FILLER_46_416 ();
 sg13g2_fill_1 FILLER_46_418 ();
 sg13g2_fill_2 FILLER_46_456 ();
 sg13g2_fill_1 FILLER_46_512 ();
 sg13g2_decap_4 FILLER_46_540 ();
 sg13g2_fill_1 FILLER_46_562 ();
 sg13g2_decap_4 FILLER_46_589 ();
 sg13g2_fill_1 FILLER_46_593 ();
 sg13g2_fill_1 FILLER_46_600 ();
 sg13g2_fill_2 FILLER_46_615 ();
 sg13g2_fill_1 FILLER_46_617 ();
 sg13g2_fill_1 FILLER_46_633 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_fill_2 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_682 ();
 sg13g2_fill_2 FILLER_46_709 ();
 sg13g2_fill_1 FILLER_46_711 ();
 sg13g2_fill_2 FILLER_46_719 ();
 sg13g2_fill_2 FILLER_46_759 ();
 sg13g2_fill_1 FILLER_46_761 ();
 sg13g2_fill_2 FILLER_46_772 ();
 sg13g2_fill_2 FILLER_46_778 ();
 sg13g2_fill_1 FILLER_46_815 ();
 sg13g2_decap_4 FILLER_46_835 ();
 sg13g2_fill_1 FILLER_46_889 ();
 sg13g2_fill_2 FILLER_46_907 ();
 sg13g2_fill_2 FILLER_46_935 ();
 sg13g2_fill_1 FILLER_46_937 ();
 sg13g2_fill_2 FILLER_46_974 ();
 sg13g2_fill_1 FILLER_46_976 ();
 sg13g2_fill_2 FILLER_46_1057 ();
 sg13g2_fill_1 FILLER_46_1059 ();
 sg13g2_fill_1 FILLER_46_1069 ();
 sg13g2_fill_2 FILLER_46_1075 ();
 sg13g2_fill_1 FILLER_46_1077 ();
 sg13g2_fill_2 FILLER_46_1082 ();
 sg13g2_fill_1 FILLER_46_1084 ();
 sg13g2_fill_1 FILLER_46_1130 ();
 sg13g2_fill_2 FILLER_46_1176 ();
 sg13g2_fill_1 FILLER_46_1191 ();
 sg13g2_fill_2 FILLER_46_1202 ();
 sg13g2_fill_1 FILLER_46_1204 ();
 sg13g2_decap_4 FILLER_46_1218 ();
 sg13g2_fill_1 FILLER_46_1291 ();
 sg13g2_fill_1 FILLER_46_1331 ();
 sg13g2_fill_2 FILLER_46_1366 ();
 sg13g2_fill_2 FILLER_46_1378 ();
 sg13g2_fill_1 FILLER_46_1383 ();
 sg13g2_fill_2 FILLER_46_1394 ();
 sg13g2_decap_8 FILLER_46_1404 ();
 sg13g2_decap_4 FILLER_46_1411 ();
 sg13g2_fill_1 FILLER_46_1460 ();
 sg13g2_fill_2 FILLER_46_1487 ();
 sg13g2_fill_1 FILLER_46_1489 ();
 sg13g2_fill_2 FILLER_46_1513 ();
 sg13g2_fill_2 FILLER_46_1519 ();
 sg13g2_fill_1 FILLER_46_1521 ();
 sg13g2_fill_1 FILLER_46_1529 ();
 sg13g2_fill_2 FILLER_46_1548 ();
 sg13g2_fill_1 FILLER_46_1550 ();
 sg13g2_fill_1 FILLER_46_1556 ();
 sg13g2_fill_1 FILLER_46_1571 ();
 sg13g2_fill_2 FILLER_46_1586 ();
 sg13g2_fill_1 FILLER_46_1588 ();
 sg13g2_decap_4 FILLER_46_1651 ();
 sg13g2_fill_1 FILLER_46_1668 ();
 sg13g2_fill_2 FILLER_46_1707 ();
 sg13g2_fill_2 FILLER_46_1724 ();
 sg13g2_fill_1 FILLER_46_1726 ();
 sg13g2_fill_1 FILLER_46_1755 ();
 sg13g2_fill_2 FILLER_46_1816 ();
 sg13g2_fill_2 FILLER_46_1827 ();
 sg13g2_fill_1 FILLER_46_1833 ();
 sg13g2_fill_2 FILLER_46_1840 ();
 sg13g2_decap_4 FILLER_46_1857 ();
 sg13g2_fill_2 FILLER_46_1861 ();
 sg13g2_fill_2 FILLER_46_1867 ();
 sg13g2_decap_8 FILLER_46_1880 ();
 sg13g2_fill_2 FILLER_46_1887 ();
 sg13g2_fill_1 FILLER_46_1893 ();
 sg13g2_fill_1 FILLER_46_1900 ();
 sg13g2_fill_1 FILLER_46_1905 ();
 sg13g2_fill_2 FILLER_46_1915 ();
 sg13g2_fill_1 FILLER_46_1917 ();
 sg13g2_fill_1 FILLER_46_1951 ();
 sg13g2_fill_2 FILLER_46_2022 ();
 sg13g2_decap_8 FILLER_46_2111 ();
 sg13g2_decap_4 FILLER_46_2118 ();
 sg13g2_fill_1 FILLER_46_2122 ();
 sg13g2_fill_2 FILLER_46_2200 ();
 sg13g2_fill_1 FILLER_46_2202 ();
 sg13g2_fill_2 FILLER_46_2239 ();
 sg13g2_fill_1 FILLER_46_2291 ();
 sg13g2_decap_4 FILLER_46_2302 ();
 sg13g2_fill_2 FILLER_46_2306 ();
 sg13g2_fill_2 FILLER_46_2346 ();
 sg13g2_fill_1 FILLER_46_2404 ();
 sg13g2_fill_2 FILLER_46_2470 ();
 sg13g2_decap_4 FILLER_46_2482 ();
 sg13g2_fill_2 FILLER_46_2532 ();
 sg13g2_fill_1 FILLER_46_2540 ();
 sg13g2_fill_1 FILLER_46_2557 ();
 sg13g2_decap_4 FILLER_46_2594 ();
 sg13g2_fill_2 FILLER_46_2634 ();
 sg13g2_fill_1 FILLER_46_2636 ();
 sg13g2_decap_8 FILLER_46_2663 ();
 sg13g2_decap_4 FILLER_46_2670 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_44 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_66 ();
 sg13g2_decap_4 FILLER_47_81 ();
 sg13g2_decap_8 FILLER_47_99 ();
 sg13g2_decap_4 FILLER_47_129 ();
 sg13g2_fill_2 FILLER_47_142 ();
 sg13g2_fill_2 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_156 ();
 sg13g2_fill_2 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_decap_4 FILLER_47_225 ();
 sg13g2_decap_4 FILLER_47_255 ();
 sg13g2_fill_1 FILLER_47_269 ();
 sg13g2_fill_2 FILLER_47_311 ();
 sg13g2_fill_1 FILLER_47_313 ();
 sg13g2_fill_2 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_385 ();
 sg13g2_fill_1 FILLER_47_394 ();
 sg13g2_fill_2 FILLER_47_400 ();
 sg13g2_decap_4 FILLER_47_482 ();
 sg13g2_fill_1 FILLER_47_486 ();
 sg13g2_fill_2 FILLER_47_531 ();
 sg13g2_fill_1 FILLER_47_533 ();
 sg13g2_fill_2 FILLER_47_540 ();
 sg13g2_fill_1 FILLER_47_542 ();
 sg13g2_fill_2 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_579 ();
 sg13g2_fill_1 FILLER_47_601 ();
 sg13g2_fill_1 FILLER_47_611 ();
 sg13g2_decap_4 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_636 ();
 sg13g2_fill_2 FILLER_47_642 ();
 sg13g2_fill_1 FILLER_47_644 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_fill_2 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_665 ();
 sg13g2_decap_4 FILLER_47_690 ();
 sg13g2_fill_1 FILLER_47_699 ();
 sg13g2_fill_1 FILLER_47_708 ();
 sg13g2_fill_1 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_720 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_2 FILLER_47_751 ();
 sg13g2_fill_2 FILLER_47_780 ();
 sg13g2_fill_1 FILLER_47_782 ();
 sg13g2_fill_1 FILLER_47_788 ();
 sg13g2_fill_2 FILLER_47_794 ();
 sg13g2_fill_1 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_837 ();
 sg13g2_decap_4 FILLER_47_844 ();
 sg13g2_fill_2 FILLER_47_848 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_fill_2 FILLER_47_945 ();
 sg13g2_fill_2 FILLER_47_953 ();
 sg13g2_fill_2 FILLER_47_983 ();
 sg13g2_fill_2 FILLER_47_1037 ();
 sg13g2_fill_1 FILLER_47_1039 ();
 sg13g2_fill_2 FILLER_47_1101 ();
 sg13g2_fill_2 FILLER_47_1107 ();
 sg13g2_fill_1 FILLER_47_1109 ();
 sg13g2_decap_8 FILLER_47_1132 ();
 sg13g2_fill_2 FILLER_47_1152 ();
 sg13g2_fill_1 FILLER_47_1163 ();
 sg13g2_fill_2 FILLER_47_1304 ();
 sg13g2_fill_2 FILLER_47_1311 ();
 sg13g2_fill_1 FILLER_47_1332 ();
 sg13g2_decap_8 FILLER_47_1351 ();
 sg13g2_fill_1 FILLER_47_1358 ();
 sg13g2_fill_1 FILLER_47_1371 ();
 sg13g2_fill_1 FILLER_47_1377 ();
 sg13g2_fill_2 FILLER_47_1386 ();
 sg13g2_fill_1 FILLER_47_1388 ();
 sg13g2_decap_4 FILLER_47_1394 ();
 sg13g2_fill_1 FILLER_47_1398 ();
 sg13g2_decap_4 FILLER_47_1403 ();
 sg13g2_fill_1 FILLER_47_1407 ();
 sg13g2_decap_4 FILLER_47_1423 ();
 sg13g2_fill_2 FILLER_47_1466 ();
 sg13g2_fill_1 FILLER_47_1468 ();
 sg13g2_fill_2 FILLER_47_1490 ();
 sg13g2_fill_1 FILLER_47_1492 ();
 sg13g2_fill_1 FILLER_47_1562 ();
 sg13g2_fill_1 FILLER_47_1602 ();
 sg13g2_decap_4 FILLER_47_1624 ();
 sg13g2_decap_4 FILLER_47_1632 ();
 sg13g2_fill_1 FILLER_47_1646 ();
 sg13g2_fill_2 FILLER_47_1777 ();
 sg13g2_fill_1 FILLER_47_1779 ();
 sg13g2_decap_4 FILLER_47_1804 ();
 sg13g2_fill_2 FILLER_47_1838 ();
 sg13g2_fill_1 FILLER_47_1840 ();
 sg13g2_fill_2 FILLER_47_1851 ();
 sg13g2_fill_2 FILLER_47_1884 ();
 sg13g2_fill_2 FILLER_47_1922 ();
 sg13g2_fill_1 FILLER_47_1924 ();
 sg13g2_decap_8 FILLER_47_1973 ();
 sg13g2_fill_1 FILLER_47_1980 ();
 sg13g2_fill_1 FILLER_47_1985 ();
 sg13g2_decap_4 FILLER_47_2000 ();
 sg13g2_fill_2 FILLER_47_2059 ();
 sg13g2_fill_1 FILLER_47_2061 ();
 sg13g2_fill_2 FILLER_47_2085 ();
 sg13g2_fill_1 FILLER_47_2122 ();
 sg13g2_fill_1 FILLER_47_2135 ();
 sg13g2_fill_2 FILLER_47_2157 ();
 sg13g2_fill_2 FILLER_47_2191 ();
 sg13g2_fill_1 FILLER_47_2193 ();
 sg13g2_fill_2 FILLER_47_2199 ();
 sg13g2_fill_1 FILLER_47_2201 ();
 sg13g2_decap_4 FILLER_47_2242 ();
 sg13g2_decap_4 FILLER_47_2272 ();
 sg13g2_fill_1 FILLER_47_2276 ();
 sg13g2_fill_2 FILLER_47_2313 ();
 sg13g2_fill_1 FILLER_47_2315 ();
 sg13g2_decap_8 FILLER_47_2395 ();
 sg13g2_fill_1 FILLER_47_2429 ();
 sg13g2_fill_1 FILLER_47_2528 ();
 sg13g2_fill_2 FILLER_47_2538 ();
 sg13g2_fill_1 FILLER_47_2540 ();
 sg13g2_fill_2 FILLER_47_2630 ();
 sg13g2_fill_1 FILLER_47_2632 ();
 sg13g2_fill_2 FILLER_47_2643 ();
 sg13g2_fill_2 FILLER_47_2671 ();
 sg13g2_fill_1 FILLER_47_2673 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_54 ();
 sg13g2_fill_1 FILLER_48_66 ();
 sg13g2_fill_2 FILLER_48_72 ();
 sg13g2_fill_1 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_87 ();
 sg13g2_fill_2 FILLER_48_107 ();
 sg13g2_fill_1 FILLER_48_122 ();
 sg13g2_fill_2 FILLER_48_145 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_decap_4 FILLER_48_159 ();
 sg13g2_fill_2 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_fill_2 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_fill_2 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_fill_1 FILLER_48_252 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_323 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_379 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_fill_2 FILLER_48_427 ();
 sg13g2_fill_2 FILLER_48_465 ();
 sg13g2_fill_2 FILLER_48_477 ();
 sg13g2_fill_2 FILLER_48_520 ();
 sg13g2_fill_1 FILLER_48_522 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_1 FILLER_48_531 ();
 sg13g2_fill_2 FILLER_48_551 ();
 sg13g2_fill_1 FILLER_48_553 ();
 sg13g2_fill_2 FILLER_48_604 ();
 sg13g2_fill_2 FILLER_48_649 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_decap_4 FILLER_48_683 ();
 sg13g2_fill_1 FILLER_48_687 ();
 sg13g2_decap_4 FILLER_48_696 ();
 sg13g2_fill_1 FILLER_48_700 ();
 sg13g2_fill_2 FILLER_48_712 ();
 sg13g2_fill_2 FILLER_48_754 ();
 sg13g2_fill_1 FILLER_48_756 ();
 sg13g2_fill_1 FILLER_48_834 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_fill_1 FILLER_48_954 ();
 sg13g2_fill_2 FILLER_48_984 ();
 sg13g2_fill_1 FILLER_48_1007 ();
 sg13g2_fill_2 FILLER_48_1142 ();
 sg13g2_fill_1 FILLER_48_1144 ();
 sg13g2_fill_1 FILLER_48_1171 ();
 sg13g2_fill_2 FILLER_48_1200 ();
 sg13g2_fill_1 FILLER_48_1219 ();
 sg13g2_fill_2 FILLER_48_1234 ();
 sg13g2_fill_1 FILLER_48_1274 ();
 sg13g2_fill_2 FILLER_48_1291 ();
 sg13g2_fill_1 FILLER_48_1304 ();
 sg13g2_fill_1 FILLER_48_1366 ();
 sg13g2_fill_2 FILLER_48_1418 ();
 sg13g2_fill_1 FILLER_48_1420 ();
 sg13g2_fill_2 FILLER_48_1456 ();
 sg13g2_fill_1 FILLER_48_1499 ();
 sg13g2_fill_2 FILLER_48_1511 ();
 sg13g2_fill_1 FILLER_48_1513 ();
 sg13g2_fill_1 FILLER_48_1549 ();
 sg13g2_fill_2 FILLER_48_1574 ();
 sg13g2_fill_2 FILLER_48_1602 ();
 sg13g2_fill_1 FILLER_48_1604 ();
 sg13g2_decap_8 FILLER_48_1631 ();
 sg13g2_fill_1 FILLER_48_1663 ();
 sg13g2_fill_1 FILLER_48_1668 ();
 sg13g2_fill_2 FILLER_48_1679 ();
 sg13g2_fill_1 FILLER_48_1681 ();
 sg13g2_fill_2 FILLER_48_1701 ();
 sg13g2_fill_1 FILLER_48_1703 ();
 sg13g2_fill_2 FILLER_48_1722 ();
 sg13g2_fill_1 FILLER_48_1724 ();
 sg13g2_fill_2 FILLER_48_1730 ();
 sg13g2_fill_1 FILLER_48_1751 ();
 sg13g2_fill_1 FILLER_48_1779 ();
 sg13g2_fill_2 FILLER_48_1816 ();
 sg13g2_fill_1 FILLER_48_1874 ();
 sg13g2_fill_2 FILLER_48_1915 ();
 sg13g2_fill_1 FILLER_48_1917 ();
 sg13g2_decap_8 FILLER_48_1958 ();
 sg13g2_fill_2 FILLER_48_1970 ();
 sg13g2_fill_1 FILLER_48_1998 ();
 sg13g2_fill_2 FILLER_48_2025 ();
 sg13g2_fill_1 FILLER_48_2027 ();
 sg13g2_fill_1 FILLER_48_2037 ();
 sg13g2_fill_2 FILLER_48_2051 ();
 sg13g2_decap_4 FILLER_48_2139 ();
 sg13g2_fill_1 FILLER_48_2143 ();
 sg13g2_fill_2 FILLER_48_2208 ();
 sg13g2_fill_2 FILLER_48_2220 ();
 sg13g2_fill_1 FILLER_48_2222 ();
 sg13g2_decap_8 FILLER_48_2273 ();
 sg13g2_fill_2 FILLER_48_2285 ();
 sg13g2_fill_1 FILLER_48_2287 ();
 sg13g2_fill_1 FILLER_48_2353 ();
 sg13g2_decap_4 FILLER_48_2359 ();
 sg13g2_fill_1 FILLER_48_2450 ();
 sg13g2_decap_8 FILLER_48_2455 ();
 sg13g2_fill_1 FILLER_48_2462 ();
 sg13g2_fill_2 FILLER_48_2506 ();
 sg13g2_fill_1 FILLER_48_2508 ();
 sg13g2_fill_2 FILLER_48_2545 ();
 sg13g2_decap_4 FILLER_48_2636 ();
 sg13g2_fill_2 FILLER_48_2640 ();
 sg13g2_fill_2 FILLER_48_2672 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_4 ();
 sg13g2_fill_2 FILLER_49_9 ();
 sg13g2_fill_2 FILLER_49_59 ();
 sg13g2_fill_1 FILLER_49_61 ();
 sg13g2_decap_4 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_181 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_decap_4 FILLER_49_194 ();
 sg13g2_fill_2 FILLER_49_198 ();
 sg13g2_decap_8 FILLER_49_205 ();
 sg13g2_fill_1 FILLER_49_212 ();
 sg13g2_fill_2 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_309 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_369 ();
 sg13g2_fill_1 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_49_381 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_405 ();
 sg13g2_fill_2 FILLER_49_508 ();
 sg13g2_fill_1 FILLER_49_510 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_fill_1 FILLER_49_616 ();
 sg13g2_fill_2 FILLER_49_626 ();
 sg13g2_fill_1 FILLER_49_628 ();
 sg13g2_fill_2 FILLER_49_637 ();
 sg13g2_fill_1 FILLER_49_639 ();
 sg13g2_fill_2 FILLER_49_646 ();
 sg13g2_decap_4 FILLER_49_658 ();
 sg13g2_fill_1 FILLER_49_662 ();
 sg13g2_fill_1 FILLER_49_699 ();
 sg13g2_fill_2 FILLER_49_742 ();
 sg13g2_fill_2 FILLER_49_750 ();
 sg13g2_fill_1 FILLER_49_777 ();
 sg13g2_fill_2 FILLER_49_845 ();
 sg13g2_fill_1 FILLER_49_847 ();
 sg13g2_fill_1 FILLER_49_878 ();
 sg13g2_fill_2 FILLER_49_937 ();
 sg13g2_fill_1 FILLER_49_939 ();
 sg13g2_fill_1 FILLER_49_995 ();
 sg13g2_fill_1 FILLER_49_1015 ();
 sg13g2_fill_2 FILLER_49_1056 ();
 sg13g2_fill_2 FILLER_49_1115 ();
 sg13g2_fill_1 FILLER_49_1117 ();
 sg13g2_fill_1 FILLER_49_1134 ();
 sg13g2_fill_1 FILLER_49_1145 ();
 sg13g2_fill_2 FILLER_49_1166 ();
 sg13g2_fill_1 FILLER_49_1168 ();
 sg13g2_fill_1 FILLER_49_1199 ();
 sg13g2_fill_2 FILLER_49_1252 ();
 sg13g2_fill_2 FILLER_49_1313 ();
 sg13g2_fill_2 FILLER_49_1325 ();
 sg13g2_fill_2 FILLER_49_1336 ();
 sg13g2_fill_2 FILLER_49_1376 ();
 sg13g2_fill_2 FILLER_49_1386 ();
 sg13g2_decap_4 FILLER_49_1398 ();
 sg13g2_fill_2 FILLER_49_1402 ();
 sg13g2_fill_2 FILLER_49_1465 ();
 sg13g2_fill_1 FILLER_49_1476 ();
 sg13g2_fill_1 FILLER_49_1560 ();
 sg13g2_decap_4 FILLER_49_1605 ();
 sg13g2_decap_4 FILLER_49_1649 ();
 sg13g2_decap_4 FILLER_49_1697 ();
 sg13g2_fill_1 FILLER_49_1737 ();
 sg13g2_decap_4 FILLER_49_1751 ();
 sg13g2_fill_2 FILLER_49_1755 ();
 sg13g2_decap_4 FILLER_49_1764 ();
 sg13g2_fill_2 FILLER_49_1768 ();
 sg13g2_fill_1 FILLER_49_1794 ();
 sg13g2_fill_2 FILLER_49_1820 ();
 sg13g2_fill_1 FILLER_49_1822 ();
 sg13g2_fill_2 FILLER_49_1836 ();
 sg13g2_fill_1 FILLER_49_1838 ();
 sg13g2_fill_1 FILLER_49_1849 ();
 sg13g2_fill_2 FILLER_49_1909 ();
 sg13g2_fill_1 FILLER_49_1911 ();
 sg13g2_fill_1 FILLER_49_1937 ();
 sg13g2_fill_2 FILLER_49_1947 ();
 sg13g2_decap_4 FILLER_49_2001 ();
 sg13g2_fill_1 FILLER_49_2005 ();
 sg13g2_fill_1 FILLER_49_2060 ();
 sg13g2_fill_2 FILLER_49_2075 ();
 sg13g2_fill_1 FILLER_49_2077 ();
 sg13g2_fill_2 FILLER_49_2087 ();
 sg13g2_fill_2 FILLER_49_2108 ();
 sg13g2_fill_1 FILLER_49_2110 ();
 sg13g2_fill_1 FILLER_49_2126 ();
 sg13g2_fill_2 FILLER_49_2136 ();
 sg13g2_fill_1 FILLER_49_2138 ();
 sg13g2_fill_2 FILLER_49_2171 ();
 sg13g2_fill_2 FILLER_49_2240 ();
 sg13g2_fill_2 FILLER_49_2349 ();
 sg13g2_decap_4 FILLER_49_2360 ();
 sg13g2_fill_1 FILLER_49_2368 ();
 sg13g2_decap_8 FILLER_49_2387 ();
 sg13g2_decap_4 FILLER_49_2394 ();
 sg13g2_fill_1 FILLER_49_2398 ();
 sg13g2_fill_1 FILLER_49_2403 ();
 sg13g2_fill_1 FILLER_49_2413 ();
 sg13g2_fill_2 FILLER_49_2427 ();
 sg13g2_fill_1 FILLER_49_2429 ();
 sg13g2_fill_2 FILLER_49_2492 ();
 sg13g2_fill_1 FILLER_49_2494 ();
 sg13g2_fill_1 FILLER_49_2570 ();
 sg13g2_decap_4 FILLER_49_2631 ();
 sg13g2_fill_1 FILLER_49_2645 ();
 sg13g2_fill_2 FILLER_49_2672 ();
 sg13g2_fill_2 FILLER_50_36 ();
 sg13g2_decap_8 FILLER_50_85 ();
 sg13g2_fill_1 FILLER_50_92 ();
 sg13g2_fill_2 FILLER_50_105 ();
 sg13g2_decap_4 FILLER_50_159 ();
 sg13g2_fill_2 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_188 ();
 sg13g2_fill_1 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_234 ();
 sg13g2_fill_2 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_fill_1 FILLER_50_293 ();
 sg13g2_fill_1 FILLER_50_312 ();
 sg13g2_fill_2 FILLER_50_360 ();
 sg13g2_fill_2 FILLER_50_399 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_462 ();
 sg13g2_fill_2 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_532 ();
 sg13g2_fill_1 FILLER_50_543 ();
 sg13g2_fill_2 FILLER_50_561 ();
 sg13g2_fill_2 FILLER_50_573 ();
 sg13g2_fill_2 FILLER_50_627 ();
 sg13g2_decap_4 FILLER_50_635 ();
 sg13g2_fill_2 FILLER_50_680 ();
 sg13g2_fill_1 FILLER_50_682 ();
 sg13g2_fill_2 FILLER_50_697 ();
 sg13g2_fill_2 FILLER_50_705 ();
 sg13g2_fill_1 FILLER_50_707 ();
 sg13g2_fill_1 FILLER_50_713 ();
 sg13g2_fill_1 FILLER_50_720 ();
 sg13g2_fill_2 FILLER_50_836 ();
 sg13g2_fill_1 FILLER_50_838 ();
 sg13g2_fill_2 FILLER_50_877 ();
 sg13g2_fill_1 FILLER_50_891 ();
 sg13g2_fill_2 FILLER_50_937 ();
 sg13g2_fill_1 FILLER_50_939 ();
 sg13g2_fill_1 FILLER_50_954 ();
 sg13g2_fill_2 FILLER_50_963 ();
 sg13g2_fill_1 FILLER_50_965 ();
 sg13g2_fill_2 FILLER_50_1035 ();
 sg13g2_fill_1 FILLER_50_1037 ();
 sg13g2_fill_2 FILLER_50_1097 ();
 sg13g2_fill_1 FILLER_50_1099 ();
 sg13g2_fill_2 FILLER_50_1117 ();
 sg13g2_fill_1 FILLER_50_1124 ();
 sg13g2_fill_2 FILLER_50_1142 ();
 sg13g2_fill_1 FILLER_50_1149 ();
 sg13g2_fill_1 FILLER_50_1269 ();
 sg13g2_fill_1 FILLER_50_1297 ();
 sg13g2_fill_2 FILLER_50_1303 ();
 sg13g2_fill_1 FILLER_50_1305 ();
 sg13g2_fill_1 FILLER_50_1341 ();
 sg13g2_fill_2 FILLER_50_1350 ();
 sg13g2_fill_1 FILLER_50_1396 ();
 sg13g2_decap_4 FILLER_50_1413 ();
 sg13g2_fill_2 FILLER_50_1478 ();
 sg13g2_fill_1 FILLER_50_1527 ();
 sg13g2_fill_2 FILLER_50_1580 ();
 sg13g2_fill_1 FILLER_50_1582 ();
 sg13g2_fill_2 FILLER_50_1610 ();
 sg13g2_fill_2 FILLER_50_1616 ();
 sg13g2_fill_1 FILLER_50_1618 ();
 sg13g2_decap_8 FILLER_50_1663 ();
 sg13g2_fill_2 FILLER_50_1670 ();
 sg13g2_fill_1 FILLER_50_1708 ();
 sg13g2_fill_1 FILLER_50_1788 ();
 sg13g2_fill_1 FILLER_50_1838 ();
 sg13g2_fill_1 FILLER_50_1868 ();
 sg13g2_fill_2 FILLER_50_1874 ();
 sg13g2_fill_1 FILLER_50_1898 ();
 sg13g2_fill_2 FILLER_50_1935 ();
 sg13g2_fill_2 FILLER_50_1957 ();
 sg13g2_fill_1 FILLER_50_1981 ();
 sg13g2_fill_2 FILLER_50_2007 ();
 sg13g2_fill_1 FILLER_50_2009 ();
 sg13g2_fill_2 FILLER_50_2024 ();
 sg13g2_fill_1 FILLER_50_2026 ();
 sg13g2_fill_2 FILLER_50_2054 ();
 sg13g2_fill_2 FILLER_50_2082 ();
 sg13g2_fill_2 FILLER_50_2139 ();
 sg13g2_decap_8 FILLER_50_2174 ();
 sg13g2_fill_2 FILLER_50_2219 ();
 sg13g2_fill_1 FILLER_50_2221 ();
 sg13g2_fill_2 FILLER_50_2240 ();
 sg13g2_fill_2 FILLER_50_2264 ();
 sg13g2_fill_2 FILLER_50_2286 ();
 sg13g2_fill_2 FILLER_50_2333 ();
 sg13g2_fill_1 FILLER_50_2379 ();
 sg13g2_fill_2 FILLER_50_2420 ();
 sg13g2_fill_1 FILLER_50_2422 ();
 sg13g2_fill_1 FILLER_50_2468 ();
 sg13g2_fill_1 FILLER_50_2488 ();
 sg13g2_fill_1 FILLER_50_2508 ();
 sg13g2_fill_1 FILLER_50_2563 ();
 sg13g2_decap_4 FILLER_50_2610 ();
 sg13g2_fill_1 FILLER_50_2614 ();
 sg13g2_fill_2 FILLER_50_2671 ();
 sg13g2_fill_1 FILLER_50_2673 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_15 ();
 sg13g2_fill_1 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_70 ();
 sg13g2_fill_2 FILLER_51_127 ();
 sg13g2_fill_1 FILLER_51_129 ();
 sg13g2_decap_4 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_155 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_decap_4 FILLER_51_170 ();
 sg13g2_decap_4 FILLER_51_189 ();
 sg13g2_fill_2 FILLER_51_208 ();
 sg13g2_fill_1 FILLER_51_210 ();
 sg13g2_decap_4 FILLER_51_221 ();
 sg13g2_decap_8 FILLER_51_230 ();
 sg13g2_fill_2 FILLER_51_237 ();
 sg13g2_decap_8 FILLER_51_244 ();
 sg13g2_decap_8 FILLER_51_255 ();
 sg13g2_decap_8 FILLER_51_262 ();
 sg13g2_fill_2 FILLER_51_269 ();
 sg13g2_fill_1 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_376 ();
 sg13g2_fill_1 FILLER_51_424 ();
 sg13g2_fill_2 FILLER_51_490 ();
 sg13g2_fill_2 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_607 ();
 sg13g2_decap_8 FILLER_51_638 ();
 sg13g2_fill_1 FILLER_51_645 ();
 sg13g2_fill_2 FILLER_51_674 ();
 sg13g2_fill_1 FILLER_51_676 ();
 sg13g2_fill_2 FILLER_51_682 ();
 sg13g2_fill_1 FILLER_51_684 ();
 sg13g2_fill_1 FILLER_51_712 ();
 sg13g2_fill_2 FILLER_51_722 ();
 sg13g2_fill_1 FILLER_51_724 ();
 sg13g2_fill_2 FILLER_51_751 ();
 sg13g2_fill_2 FILLER_51_770 ();
 sg13g2_fill_1 FILLER_51_772 ();
 sg13g2_fill_1 FILLER_51_791 ();
 sg13g2_fill_1 FILLER_51_801 ();
 sg13g2_fill_1 FILLER_51_867 ();
 sg13g2_fill_2 FILLER_51_891 ();
 sg13g2_fill_2 FILLER_51_928 ();
 sg13g2_fill_2 FILLER_51_956 ();
 sg13g2_fill_1 FILLER_51_958 ();
 sg13g2_fill_2 FILLER_51_986 ();
 sg13g2_fill_1 FILLER_51_988 ();
 sg13g2_fill_1 FILLER_51_1028 ();
 sg13g2_fill_2 FILLER_51_1094 ();
 sg13g2_fill_1 FILLER_51_1096 ();
 sg13g2_fill_2 FILLER_51_1111 ();
 sg13g2_fill_2 FILLER_51_1165 ();
 sg13g2_fill_1 FILLER_51_1167 ();
 sg13g2_fill_2 FILLER_51_1171 ();
 sg13g2_fill_1 FILLER_51_1173 ();
 sg13g2_fill_2 FILLER_51_1299 ();
 sg13g2_fill_2 FILLER_51_1306 ();
 sg13g2_decap_4 FILLER_51_1318 ();
 sg13g2_fill_1 FILLER_51_1357 ();
 sg13g2_fill_1 FILLER_51_1401 ();
 sg13g2_fill_2 FILLER_51_1418 ();
 sg13g2_fill_1 FILLER_51_1448 ();
 sg13g2_fill_2 FILLER_51_1569 ();
 sg13g2_fill_1 FILLER_51_1571 ();
 sg13g2_fill_2 FILLER_51_1589 ();
 sg13g2_fill_2 FILLER_51_1605 ();
 sg13g2_fill_2 FILLER_51_1627 ();
 sg13g2_fill_1 FILLER_51_1629 ();
 sg13g2_fill_1 FILLER_51_1720 ();
 sg13g2_fill_2 FILLER_51_1747 ();
 sg13g2_fill_1 FILLER_51_1764 ();
 sg13g2_fill_2 FILLER_51_1798 ();
 sg13g2_fill_2 FILLER_51_1866 ();
 sg13g2_fill_1 FILLER_51_1868 ();
 sg13g2_fill_2 FILLER_51_1879 ();
 sg13g2_fill_1 FILLER_51_1881 ();
 sg13g2_fill_2 FILLER_51_1908 ();
 sg13g2_fill_1 FILLER_51_1910 ();
 sg13g2_fill_2 FILLER_51_1942 ();
 sg13g2_fill_2 FILLER_51_1958 ();
 sg13g2_fill_1 FILLER_51_1960 ();
 sg13g2_fill_2 FILLER_51_1970 ();
 sg13g2_fill_1 FILLER_51_1972 ();
 sg13g2_fill_1 FILLER_51_1977 ();
 sg13g2_fill_2 FILLER_51_1982 ();
 sg13g2_fill_1 FILLER_51_1984 ();
 sg13g2_fill_2 FILLER_51_1995 ();
 sg13g2_fill_1 FILLER_51_1997 ();
 sg13g2_fill_2 FILLER_51_2003 ();
 sg13g2_fill_1 FILLER_51_2052 ();
 sg13g2_fill_2 FILLER_51_2070 ();
 sg13g2_fill_1 FILLER_51_2072 ();
 sg13g2_fill_2 FILLER_51_2090 ();
 sg13g2_fill_1 FILLER_51_2092 ();
 sg13g2_fill_2 FILLER_51_2106 ();
 sg13g2_fill_1 FILLER_51_2108 ();
 sg13g2_fill_1 FILLER_51_2115 ();
 sg13g2_fill_2 FILLER_51_2121 ();
 sg13g2_fill_1 FILLER_51_2123 ();
 sg13g2_fill_2 FILLER_51_2133 ();
 sg13g2_fill_1 FILLER_51_2135 ();
 sg13g2_fill_2 FILLER_51_2186 ();
 sg13g2_fill_1 FILLER_51_2205 ();
 sg13g2_decap_4 FILLER_51_2302 ();
 sg13g2_fill_2 FILLER_51_2306 ();
 sg13g2_decap_4 FILLER_51_2365 ();
 sg13g2_fill_1 FILLER_51_2369 ();
 sg13g2_fill_2 FILLER_51_2405 ();
 sg13g2_fill_1 FILLER_51_2407 ();
 sg13g2_fill_2 FILLER_51_2527 ();
 sg13g2_fill_1 FILLER_51_2552 ();
 sg13g2_fill_1 FILLER_51_2569 ();
 sg13g2_fill_2 FILLER_51_2585 ();
 sg13g2_fill_2 FILLER_51_2592 ();
 sg13g2_decap_4 FILLER_51_2607 ();
 sg13g2_fill_2 FILLER_51_2621 ();
 sg13g2_fill_1 FILLER_51_2623 ();
 sg13g2_decap_8 FILLER_51_2637 ();
 sg13g2_decap_4 FILLER_51_2644 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_35 ();
 sg13g2_fill_1 FILLER_52_86 ();
 sg13g2_fill_1 FILLER_52_104 ();
 sg13g2_fill_2 FILLER_52_111 ();
 sg13g2_fill_1 FILLER_52_113 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_172 ();
 sg13g2_decap_4 FILLER_52_179 ();
 sg13g2_decap_8 FILLER_52_187 ();
 sg13g2_fill_2 FILLER_52_249 ();
 sg13g2_fill_2 FILLER_52_286 ();
 sg13g2_fill_2 FILLER_52_302 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_2 FILLER_52_353 ();
 sg13g2_fill_1 FILLER_52_416 ();
 sg13g2_fill_2 FILLER_52_447 ();
 sg13g2_fill_1 FILLER_52_449 ();
 sg13g2_fill_1 FILLER_52_464 ();
 sg13g2_fill_1 FILLER_52_483 ();
 sg13g2_fill_2 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_566 ();
 sg13g2_fill_2 FILLER_52_597 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_fill_1 FILLER_52_735 ();
 sg13g2_fill_1 FILLER_52_745 ();
 sg13g2_fill_2 FILLER_52_781 ();
 sg13g2_fill_1 FILLER_52_807 ();
 sg13g2_fill_1 FILLER_52_817 ();
 sg13g2_fill_1 FILLER_52_830 ();
 sg13g2_fill_2 FILLER_52_857 ();
 sg13g2_fill_2 FILLER_52_916 ();
 sg13g2_fill_1 FILLER_52_918 ();
 sg13g2_fill_2 FILLER_52_942 ();
 sg13g2_fill_1 FILLER_52_944 ();
 sg13g2_fill_2 FILLER_52_979 ();
 sg13g2_fill_2 FILLER_52_1123 ();
 sg13g2_fill_1 FILLER_52_1125 ();
 sg13g2_fill_2 FILLER_52_1136 ();
 sg13g2_fill_1 FILLER_52_1138 ();
 sg13g2_fill_2 FILLER_52_1152 ();
 sg13g2_fill_1 FILLER_52_1181 ();
 sg13g2_fill_1 FILLER_52_1203 ();
 sg13g2_fill_2 FILLER_52_1232 ();
 sg13g2_fill_1 FILLER_52_1312 ();
 sg13g2_fill_2 FILLER_52_1331 ();
 sg13g2_decap_8 FILLER_52_1367 ();
 sg13g2_decap_8 FILLER_52_1374 ();
 sg13g2_fill_2 FILLER_52_1381 ();
 sg13g2_decap_4 FILLER_52_1387 ();
 sg13g2_fill_2 FILLER_52_1391 ();
 sg13g2_fill_1 FILLER_52_1402 ();
 sg13g2_fill_2 FILLER_52_1458 ();
 sg13g2_fill_2 FILLER_52_1490 ();
 sg13g2_fill_2 FILLER_52_1537 ();
 sg13g2_fill_1 FILLER_52_1539 ();
 sg13g2_fill_2 FILLER_52_1554 ();
 sg13g2_fill_1 FILLER_52_1626 ();
 sg13g2_fill_1 FILLER_52_1632 ();
 sg13g2_fill_2 FILLER_52_1654 ();
 sg13g2_decap_4 FILLER_52_1708 ();
 sg13g2_fill_1 FILLER_52_1731 ();
 sg13g2_fill_2 FILLER_52_1747 ();
 sg13g2_fill_1 FILLER_52_1749 ();
 sg13g2_fill_1 FILLER_52_1776 ();
 sg13g2_fill_1 FILLER_52_1802 ();
 sg13g2_fill_1 FILLER_52_1903 ();
 sg13g2_fill_2 FILLER_52_1909 ();
 sg13g2_fill_2 FILLER_52_1972 ();
 sg13g2_fill_1 FILLER_52_1974 ();
 sg13g2_fill_2 FILLER_52_1994 ();
 sg13g2_fill_2 FILLER_52_2032 ();
 sg13g2_fill_2 FILLER_52_2071 ();
 sg13g2_fill_2 FILLER_52_2107 ();
 sg13g2_fill_1 FILLER_52_2129 ();
 sg13g2_fill_1 FILLER_52_2145 ();
 sg13g2_decap_4 FILLER_52_2167 ();
 sg13g2_fill_2 FILLER_52_2175 ();
 sg13g2_fill_1 FILLER_52_2177 ();
 sg13g2_fill_2 FILLER_52_2259 ();
 sg13g2_fill_1 FILLER_52_2261 ();
 sg13g2_decap_4 FILLER_52_2275 ();
 sg13g2_decap_4 FILLER_52_2289 ();
 sg13g2_fill_2 FILLER_52_2303 ();
 sg13g2_fill_2 FILLER_52_2322 ();
 sg13g2_fill_1 FILLER_52_2324 ();
 sg13g2_decap_4 FILLER_52_2364 ();
 sg13g2_decap_4 FILLER_52_2381 ();
 sg13g2_fill_1 FILLER_52_2395 ();
 sg13g2_fill_1 FILLER_52_2464 ();
 sg13g2_fill_1 FILLER_52_2479 ();
 sg13g2_fill_2 FILLER_52_2561 ();
 sg13g2_fill_2 FILLER_52_2597 ();
 sg13g2_fill_1 FILLER_52_2599 ();
 sg13g2_fill_1 FILLER_52_2608 ();
 sg13g2_decap_4 FILLER_52_2619 ();
 sg13g2_fill_2 FILLER_52_2646 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_fill_1 FILLER_53_29 ();
 sg13g2_fill_2 FILLER_53_83 ();
 sg13g2_fill_1 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_decap_4 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_144 ();
 sg13g2_fill_1 FILLER_53_156 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_decap_4 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_202 ();
 sg13g2_decap_4 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_216 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_278 ();
 sg13g2_fill_1 FILLER_53_280 ();
 sg13g2_fill_2 FILLER_53_285 ();
 sg13g2_fill_1 FILLER_53_287 ();
 sg13g2_fill_2 FILLER_53_302 ();
 sg13g2_fill_1 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_311 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_fill_1 FILLER_53_361 ();
 sg13g2_fill_1 FILLER_53_440 ();
 sg13g2_fill_2 FILLER_53_451 ();
 sg13g2_fill_2 FILLER_53_466 ();
 sg13g2_fill_2 FILLER_53_472 ();
 sg13g2_fill_2 FILLER_53_489 ();
 sg13g2_fill_1 FILLER_53_501 ();
 sg13g2_fill_2 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_536 ();
 sg13g2_fill_1 FILLER_53_557 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_fill_1 FILLER_53_606 ();
 sg13g2_fill_1 FILLER_53_616 ();
 sg13g2_fill_1 FILLER_53_646 ();
 sg13g2_fill_2 FILLER_53_657 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_1 FILLER_53_759 ();
 sg13g2_fill_2 FILLER_53_822 ();
 sg13g2_fill_1 FILLER_53_839 ();
 sg13g2_fill_1 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_fill_2 FILLER_53_888 ();
 sg13g2_fill_1 FILLER_53_908 ();
 sg13g2_fill_1 FILLER_53_919 ();
 sg13g2_fill_2 FILLER_53_925 ();
 sg13g2_fill_2 FILLER_53_965 ();
 sg13g2_fill_2 FILLER_53_977 ();
 sg13g2_fill_1 FILLER_53_991 ();
 sg13g2_fill_1 FILLER_53_1010 ();
 sg13g2_fill_2 FILLER_53_1016 ();
 sg13g2_fill_1 FILLER_53_1086 ();
 sg13g2_fill_2 FILLER_53_1092 ();
 sg13g2_fill_1 FILLER_53_1094 ();
 sg13g2_decap_4 FILLER_53_1157 ();
 sg13g2_fill_2 FILLER_53_1166 ();
 sg13g2_fill_2 FILLER_53_1247 ();
 sg13g2_fill_1 FILLER_53_1249 ();
 sg13g2_fill_1 FILLER_53_1302 ();
 sg13g2_fill_1 FILLER_53_1371 ();
 sg13g2_fill_1 FILLER_53_1398 ();
 sg13g2_fill_2 FILLER_53_1455 ();
 sg13g2_fill_1 FILLER_53_1457 ();
 sg13g2_decap_8 FILLER_53_1463 ();
 sg13g2_fill_1 FILLER_53_1470 ();
 sg13g2_fill_2 FILLER_53_1479 ();
 sg13g2_fill_2 FILLER_53_1524 ();
 sg13g2_fill_1 FILLER_53_1574 ();
 sg13g2_fill_2 FILLER_53_1589 ();
 sg13g2_fill_2 FILLER_53_1619 ();
 sg13g2_fill_1 FILLER_53_1629 ();
 sg13g2_fill_1 FILLER_53_1649 ();
 sg13g2_fill_2 FILLER_53_1667 ();
 sg13g2_fill_1 FILLER_53_1669 ();
 sg13g2_fill_1 FILLER_53_1692 ();
 sg13g2_fill_2 FILLER_53_1721 ();
 sg13g2_decap_4 FILLER_53_1806 ();
 sg13g2_fill_1 FILLER_53_1884 ();
 sg13g2_fill_2 FILLER_53_1958 ();
 sg13g2_decap_4 FILLER_53_1990 ();
 sg13g2_fill_1 FILLER_53_1994 ();
 sg13g2_decap_8 FILLER_53_2000 ();
 sg13g2_fill_2 FILLER_53_2007 ();
 sg13g2_fill_2 FILLER_53_2015 ();
 sg13g2_fill_1 FILLER_53_2017 ();
 sg13g2_fill_1 FILLER_53_2040 ();
 sg13g2_fill_2 FILLER_53_2054 ();
 sg13g2_fill_2 FILLER_53_2068 ();
 sg13g2_fill_1 FILLER_53_2070 ();
 sg13g2_fill_2 FILLER_53_2079 ();
 sg13g2_fill_2 FILLER_53_2086 ();
 sg13g2_fill_1 FILLER_53_2088 ();
 sg13g2_fill_1 FILLER_53_2137 ();
 sg13g2_fill_2 FILLER_53_2195 ();
 sg13g2_fill_1 FILLER_53_2197 ();
 sg13g2_fill_2 FILLER_53_2221 ();
 sg13g2_fill_2 FILLER_53_2339 ();
 sg13g2_fill_1 FILLER_53_2341 ();
 sg13g2_fill_2 FILLER_53_2472 ();
 sg13g2_fill_2 FILLER_53_2507 ();
 sg13g2_fill_1 FILLER_53_2509 ();
 sg13g2_fill_2 FILLER_53_2546 ();
 sg13g2_fill_1 FILLER_53_2548 ();
 sg13g2_fill_1 FILLER_53_2673 ();
 sg13g2_fill_2 FILLER_54_73 ();
 sg13g2_fill_2 FILLER_54_124 ();
 sg13g2_fill_1 FILLER_54_131 ();
 sg13g2_fill_1 FILLER_54_137 ();
 sg13g2_decap_4 FILLER_54_142 ();
 sg13g2_decap_4 FILLER_54_202 ();
 sg13g2_fill_2 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_297 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_2 FILLER_54_323 ();
 sg13g2_fill_1 FILLER_54_358 ();
 sg13g2_fill_2 FILLER_54_440 ();
 sg13g2_fill_1 FILLER_54_442 ();
 sg13g2_fill_2 FILLER_54_534 ();
 sg13g2_fill_2 FILLER_54_588 ();
 sg13g2_fill_1 FILLER_54_590 ();
 sg13g2_fill_1 FILLER_54_630 ();
 sg13g2_fill_2 FILLER_54_666 ();
 sg13g2_fill_2 FILLER_54_702 ();
 sg13g2_fill_1 FILLER_54_740 ();
 sg13g2_fill_2 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_807 ();
 sg13g2_fill_2 FILLER_54_850 ();
 sg13g2_fill_2 FILLER_54_878 ();
 sg13g2_fill_2 FILLER_54_994 ();
 sg13g2_fill_2 FILLER_54_1038 ();
 sg13g2_fill_2 FILLER_54_1089 ();
 sg13g2_fill_1 FILLER_54_1091 ();
 sg13g2_fill_1 FILLER_54_1146 ();
 sg13g2_fill_1 FILLER_54_1198 ();
 sg13g2_fill_2 FILLER_54_1207 ();
 sg13g2_fill_1 FILLER_54_1237 ();
 sg13g2_fill_1 FILLER_54_1286 ();
 sg13g2_fill_2 FILLER_54_1295 ();
 sg13g2_fill_2 FILLER_54_1337 ();
 sg13g2_fill_1 FILLER_54_1339 ();
 sg13g2_fill_2 FILLER_54_1346 ();
 sg13g2_fill_1 FILLER_54_1348 ();
 sg13g2_fill_1 FILLER_54_1354 ();
 sg13g2_fill_2 FILLER_54_1396 ();
 sg13g2_fill_1 FILLER_54_1398 ();
 sg13g2_fill_2 FILLER_54_1419 ();
 sg13g2_fill_1 FILLER_54_1421 ();
 sg13g2_fill_1 FILLER_54_1432 ();
 sg13g2_fill_1 FILLER_54_1464 ();
 sg13g2_fill_2 FILLER_54_1503 ();
 sg13g2_fill_2 FILLER_54_1597 ();
 sg13g2_fill_1 FILLER_54_1607 ();
 sg13g2_fill_2 FILLER_54_1620 ();
 sg13g2_decap_4 FILLER_54_1635 ();
 sg13g2_decap_8 FILLER_54_1652 ();
 sg13g2_fill_2 FILLER_54_1710 ();
 sg13g2_fill_2 FILLER_54_1715 ();
 sg13g2_fill_1 FILLER_54_1726 ();
 sg13g2_fill_2 FILLER_54_1737 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_fill_1 FILLER_54_1768 ();
 sg13g2_decap_8 FILLER_54_1783 ();
 sg13g2_fill_1 FILLER_54_1910 ();
 sg13g2_fill_2 FILLER_54_1942 ();
 sg13g2_fill_1 FILLER_54_1944 ();
 sg13g2_fill_1 FILLER_54_1975 ();
 sg13g2_fill_2 FILLER_54_1985 ();
 sg13g2_fill_1 FILLER_54_1987 ();
 sg13g2_decap_8 FILLER_54_2024 ();
 sg13g2_fill_2 FILLER_54_2040 ();
 sg13g2_fill_1 FILLER_54_2042 ();
 sg13g2_decap_4 FILLER_54_2065 ();
 sg13g2_fill_1 FILLER_54_2069 ();
 sg13g2_fill_2 FILLER_54_2095 ();
 sg13g2_fill_1 FILLER_54_2097 ();
 sg13g2_fill_2 FILLER_54_2107 ();
 sg13g2_fill_1 FILLER_54_2109 ();
 sg13g2_fill_2 FILLER_54_2176 ();
 sg13g2_fill_1 FILLER_54_2178 ();
 sg13g2_fill_2 FILLER_54_2266 ();
 sg13g2_fill_1 FILLER_54_2287 ();
 sg13g2_fill_2 FILLER_54_2298 ();
 sg13g2_fill_1 FILLER_54_2300 ();
 sg13g2_fill_1 FILLER_54_2314 ();
 sg13g2_decap_4 FILLER_54_2364 ();
 sg13g2_fill_1 FILLER_54_2378 ();
 sg13g2_fill_1 FILLER_54_2403 ();
 sg13g2_fill_1 FILLER_54_2427 ();
 sg13g2_fill_2 FILLER_54_2440 ();
 sg13g2_fill_1 FILLER_54_2442 ();
 sg13g2_fill_2 FILLER_54_2545 ();
 sg13g2_fill_2 FILLER_54_2613 ();
 sg13g2_fill_1 FILLER_54_2615 ();
 sg13g2_fill_2 FILLER_54_2622 ();
 sg13g2_fill_1 FILLER_54_2624 ();
 sg13g2_fill_2 FILLER_54_2645 ();
 sg13g2_fill_1 FILLER_54_2647 ();
 sg13g2_fill_1 FILLER_55_71 ();
 sg13g2_fill_2 FILLER_55_90 ();
 sg13g2_fill_1 FILLER_55_92 ();
 sg13g2_decap_4 FILLER_55_107 ();
 sg13g2_fill_2 FILLER_55_111 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_fill_2 FILLER_55_146 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_fill_2 FILLER_55_192 ();
 sg13g2_fill_1 FILLER_55_204 ();
 sg13g2_fill_2 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_226 ();
 sg13g2_fill_1 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_276 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_fill_2 FILLER_55_368 ();
 sg13g2_fill_1 FILLER_55_370 ();
 sg13g2_fill_1 FILLER_55_445 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_2 FILLER_55_469 ();
 sg13g2_fill_1 FILLER_55_471 ();
 sg13g2_fill_2 FILLER_55_481 ();
 sg13g2_fill_1 FILLER_55_504 ();
 sg13g2_fill_2 FILLER_55_584 ();
 sg13g2_fill_1 FILLER_55_586 ();
 sg13g2_fill_2 FILLER_55_606 ();
 sg13g2_fill_2 FILLER_55_638 ();
 sg13g2_fill_1 FILLER_55_640 ();
 sg13g2_fill_2 FILLER_55_664 ();
 sg13g2_fill_1 FILLER_55_676 ();
 sg13g2_fill_1 FILLER_55_696 ();
 sg13g2_fill_1 FILLER_55_701 ();
 sg13g2_fill_1 FILLER_55_768 ();
 sg13g2_fill_1 FILLER_55_777 ();
 sg13g2_fill_2 FILLER_55_804 ();
 sg13g2_fill_1 FILLER_55_806 ();
 sg13g2_fill_2 FILLER_55_838 ();
 sg13g2_fill_2 FILLER_55_849 ();
 sg13g2_fill_1 FILLER_55_851 ();
 sg13g2_fill_2 FILLER_55_895 ();
 sg13g2_fill_1 FILLER_55_897 ();
 sg13g2_fill_2 FILLER_55_924 ();
 sg13g2_fill_1 FILLER_55_926 ();
 sg13g2_fill_2 FILLER_55_949 ();
 sg13g2_fill_2 FILLER_55_1064 ();
 sg13g2_fill_1 FILLER_55_1066 ();
 sg13g2_fill_1 FILLER_55_1083 ();
 sg13g2_fill_1 FILLER_55_1110 ();
 sg13g2_fill_2 FILLER_55_1152 ();
 sg13g2_fill_1 FILLER_55_1154 ();
 sg13g2_fill_2 FILLER_55_1161 ();
 sg13g2_fill_1 FILLER_55_1189 ();
 sg13g2_fill_2 FILLER_55_1295 ();
 sg13g2_fill_2 FILLER_55_1355 ();
 sg13g2_fill_1 FILLER_55_1357 ();
 sg13g2_fill_1 FILLER_55_1402 ();
 sg13g2_fill_2 FILLER_55_1422 ();
 sg13g2_fill_2 FILLER_55_1437 ();
 sg13g2_fill_2 FILLER_55_1482 ();
 sg13g2_fill_2 FILLER_55_1635 ();
 sg13g2_decap_4 FILLER_55_1657 ();
 sg13g2_decap_4 FILLER_55_1756 ();
 sg13g2_fill_2 FILLER_55_1822 ();
 sg13g2_fill_1 FILLER_55_1828 ();
 sg13g2_fill_1 FILLER_55_1924 ();
 sg13g2_fill_2 FILLER_55_1939 ();
 sg13g2_fill_1 FILLER_55_1941 ();
 sg13g2_fill_2 FILLER_55_1957 ();
 sg13g2_fill_1 FILLER_55_1978 ();
 sg13g2_fill_2 FILLER_55_1987 ();
 sg13g2_fill_1 FILLER_55_1995 ();
 sg13g2_fill_2 FILLER_55_2002 ();
 sg13g2_fill_1 FILLER_55_2004 ();
 sg13g2_fill_2 FILLER_55_2025 ();
 sg13g2_decap_4 FILLER_55_2040 ();
 sg13g2_decap_4 FILLER_55_2052 ();
 sg13g2_fill_1 FILLER_55_2080 ();
 sg13g2_fill_1 FILLER_55_2139 ();
 sg13g2_fill_1 FILLER_55_2144 ();
 sg13g2_fill_1 FILLER_55_2163 ();
 sg13g2_fill_2 FILLER_55_2178 ();
 sg13g2_fill_1 FILLER_55_2180 ();
 sg13g2_fill_2 FILLER_55_2218 ();
 sg13g2_fill_1 FILLER_55_2220 ();
 sg13g2_fill_2 FILLER_55_2238 ();
 sg13g2_fill_1 FILLER_55_2274 ();
 sg13g2_fill_2 FILLER_55_2289 ();
 sg13g2_fill_1 FILLER_55_2327 ();
 sg13g2_fill_1 FILLER_55_2434 ();
 sg13g2_fill_1 FILLER_55_2491 ();
 sg13g2_fill_1 FILLER_55_2543 ();
 sg13g2_fill_1 FILLER_55_2585 ();
 sg13g2_fill_1 FILLER_55_2642 ();
 sg13g2_fill_1 FILLER_55_2673 ();
 sg13g2_fill_2 FILLER_56_64 ();
 sg13g2_decap_4 FILLER_56_79 ();
 sg13g2_fill_2 FILLER_56_83 ();
 sg13g2_decap_4 FILLER_56_105 ();
 sg13g2_decap_4 FILLER_56_149 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_fill_2 FILLER_56_169 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_182 ();
 sg13g2_fill_1 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_194 ();
 sg13g2_fill_2 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_206 ();
 sg13g2_fill_1 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_fill_2 FILLER_56_352 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_fill_1 FILLER_56_501 ();
 sg13g2_fill_1 FILLER_56_507 ();
 sg13g2_fill_2 FILLER_56_603 ();
 sg13g2_fill_1 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_611 ();
 sg13g2_fill_2 FILLER_56_621 ();
 sg13g2_fill_2 FILLER_56_627 ();
 sg13g2_fill_1 FILLER_56_635 ();
 sg13g2_fill_1 FILLER_56_667 ();
 sg13g2_fill_2 FILLER_56_694 ();
 sg13g2_fill_1 FILLER_56_696 ();
 sg13g2_fill_1 FILLER_56_728 ();
 sg13g2_fill_2 FILLER_56_756 ();
 sg13g2_fill_1 FILLER_56_758 ();
 sg13g2_fill_2 FILLER_56_775 ();
 sg13g2_fill_2 FILLER_56_801 ();
 sg13g2_fill_1 FILLER_56_803 ();
 sg13g2_fill_1 FILLER_56_808 ();
 sg13g2_fill_2 FILLER_56_830 ();
 sg13g2_fill_2 FILLER_56_841 ();
 sg13g2_fill_1 FILLER_56_852 ();
 sg13g2_fill_2 FILLER_56_880 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_fill_1 FILLER_56_892 ();
 sg13g2_fill_2 FILLER_56_898 ();
 sg13g2_fill_2 FILLER_56_942 ();
 sg13g2_fill_1 FILLER_56_1003 ();
 sg13g2_fill_2 FILLER_56_1027 ();
 sg13g2_fill_1 FILLER_56_1034 ();
 sg13g2_fill_2 FILLER_56_1040 ();
 sg13g2_fill_1 FILLER_56_1042 ();
 sg13g2_fill_1 FILLER_56_1092 ();
 sg13g2_fill_2 FILLER_56_1102 ();
 sg13g2_fill_1 FILLER_56_1114 ();
 sg13g2_fill_2 FILLER_56_1138 ();
 sg13g2_fill_1 FILLER_56_1140 ();
 sg13g2_fill_1 FILLER_56_1184 ();
 sg13g2_fill_2 FILLER_56_1220 ();
 sg13g2_fill_2 FILLER_56_1247 ();
 sg13g2_fill_1 FILLER_56_1249 ();
 sg13g2_decap_4 FILLER_56_1324 ();
 sg13g2_fill_1 FILLER_56_1336 ();
 sg13g2_decap_4 FILLER_56_1354 ();
 sg13g2_fill_2 FILLER_56_1358 ();
 sg13g2_fill_1 FILLER_56_1365 ();
 sg13g2_fill_1 FILLER_56_1373 ();
 sg13g2_fill_1 FILLER_56_1419 ();
 sg13g2_fill_2 FILLER_56_1437 ();
 sg13g2_fill_2 FILLER_56_1465 ();
 sg13g2_fill_1 FILLER_56_1467 ();
 sg13g2_fill_1 FILLER_56_1538 ();
 sg13g2_fill_2 FILLER_56_1545 ();
 sg13g2_fill_1 FILLER_56_1547 ();
 sg13g2_fill_1 FILLER_56_1557 ();
 sg13g2_fill_1 FILLER_56_1577 ();
 sg13g2_fill_2 FILLER_56_1586 ();
 sg13g2_fill_2 FILLER_56_1596 ();
 sg13g2_fill_1 FILLER_56_1598 ();
 sg13g2_decap_4 FILLER_56_1641 ();
 sg13g2_decap_8 FILLER_56_1661 ();
 sg13g2_fill_1 FILLER_56_1668 ();
 sg13g2_fill_2 FILLER_56_1712 ();
 sg13g2_fill_1 FILLER_56_1768 ();
 sg13g2_fill_1 FILLER_56_1782 ();
 sg13g2_fill_1 FILLER_56_1870 ();
 sg13g2_fill_1 FILLER_56_1892 ();
 sg13g2_fill_2 FILLER_56_1923 ();
 sg13g2_fill_2 FILLER_56_1946 ();
 sg13g2_fill_1 FILLER_56_1948 ();
 sg13g2_fill_1 FILLER_56_1970 ();
 sg13g2_fill_1 FILLER_56_1983 ();
 sg13g2_fill_1 FILLER_56_2042 ();
 sg13g2_fill_1 FILLER_56_2068 ();
 sg13g2_fill_2 FILLER_56_2107 ();
 sg13g2_fill_2 FILLER_56_2156 ();
 sg13g2_fill_1 FILLER_56_2219 ();
 sg13g2_decap_4 FILLER_56_2265 ();
 sg13g2_fill_1 FILLER_56_2269 ();
 sg13g2_fill_2 FILLER_56_2332 ();
 sg13g2_decap_4 FILLER_56_2340 ();
 sg13g2_fill_1 FILLER_56_2344 ();
 sg13g2_fill_2 FILLER_56_2377 ();
 sg13g2_fill_1 FILLER_56_2379 ();
 sg13g2_fill_2 FILLER_56_2451 ();
 sg13g2_fill_1 FILLER_56_2453 ();
 sg13g2_fill_2 FILLER_56_2463 ();
 sg13g2_fill_2 FILLER_56_2474 ();
 sg13g2_fill_1 FILLER_56_2476 ();
 sg13g2_fill_1 FILLER_56_2549 ();
 sg13g2_decap_8 FILLER_56_2585 ();
 sg13g2_fill_2 FILLER_56_2592 ();
 sg13g2_fill_2 FILLER_56_2626 ();
 sg13g2_fill_2 FILLER_56_2649 ();
 sg13g2_fill_1 FILLER_56_2651 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_41 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_2 FILLER_57_120 ();
 sg13g2_fill_1 FILLER_57_145 ();
 sg13g2_fill_1 FILLER_57_154 ();
 sg13g2_fill_2 FILLER_57_192 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_222 ();
 sg13g2_fill_2 FILLER_57_254 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_278 ();
 sg13g2_fill_2 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_376 ();
 sg13g2_fill_2 FILLER_57_392 ();
 sg13g2_fill_2 FILLER_57_418 ();
 sg13g2_fill_1 FILLER_57_420 ();
 sg13g2_fill_2 FILLER_57_434 ();
 sg13g2_fill_1 FILLER_57_436 ();
 sg13g2_fill_2 FILLER_57_442 ();
 sg13g2_fill_2 FILLER_57_453 ();
 sg13g2_fill_1 FILLER_57_455 ();
 sg13g2_fill_2 FILLER_57_473 ();
 sg13g2_fill_1 FILLER_57_475 ();
 sg13g2_fill_2 FILLER_57_485 ();
 sg13g2_fill_1 FILLER_57_487 ();
 sg13g2_fill_2 FILLER_57_493 ();
 sg13g2_fill_2 FILLER_57_510 ();
 sg13g2_fill_1 FILLER_57_534 ();
 sg13g2_fill_2 FILLER_57_565 ();
 sg13g2_fill_1 FILLER_57_576 ();
 sg13g2_fill_2 FILLER_57_600 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_649 ();
 sg13g2_fill_1 FILLER_57_662 ();
 sg13g2_fill_2 FILLER_57_681 ();
 sg13g2_fill_1 FILLER_57_683 ();
 sg13g2_fill_1 FILLER_57_690 ();
 sg13g2_fill_2 FILLER_57_816 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_fill_1 FILLER_57_854 ();
 sg13g2_fill_2 FILLER_57_887 ();
 sg13g2_fill_2 FILLER_57_941 ();
 sg13g2_fill_1 FILLER_57_960 ();
 sg13g2_fill_1 FILLER_57_981 ();
 sg13g2_fill_2 FILLER_57_1026 ();
 sg13g2_fill_1 FILLER_57_1063 ();
 sg13g2_fill_2 FILLER_57_1087 ();
 sg13g2_fill_1 FILLER_57_1089 ();
 sg13g2_fill_2 FILLER_57_1131 ();
 sg13g2_fill_1 FILLER_57_1159 ();
 sg13g2_fill_2 FILLER_57_1177 ();
 sg13g2_fill_1 FILLER_57_1179 ();
 sg13g2_fill_2 FILLER_57_1230 ();
 sg13g2_fill_2 FILLER_57_1240 ();
 sg13g2_decap_8 FILLER_57_1251 ();
 sg13g2_fill_2 FILLER_57_1258 ();
 sg13g2_fill_1 FILLER_57_1260 ();
 sg13g2_fill_1 FILLER_57_1274 ();
 sg13g2_fill_2 FILLER_57_1288 ();
 sg13g2_fill_1 FILLER_57_1290 ();
 sg13g2_fill_2 FILLER_57_1310 ();
 sg13g2_fill_1 FILLER_57_1312 ();
 sg13g2_fill_1 FILLER_57_1318 ();
 sg13g2_fill_1 FILLER_57_1360 ();
 sg13g2_fill_1 FILLER_57_1397 ();
 sg13g2_fill_2 FILLER_57_1424 ();
 sg13g2_fill_2 FILLER_57_1432 ();
 sg13g2_fill_1 FILLER_57_1434 ();
 sg13g2_fill_1 FILLER_57_1445 ();
 sg13g2_fill_1 FILLER_57_1455 ();
 sg13g2_fill_2 FILLER_57_1469 ();
 sg13g2_fill_2 FILLER_57_1480 ();
 sg13g2_fill_1 FILLER_57_1482 ();
 sg13g2_fill_2 FILLER_57_1506 ();
 sg13g2_fill_1 FILLER_57_1508 ();
 sg13g2_fill_2 FILLER_57_1573 ();
 sg13g2_fill_2 FILLER_57_1600 ();
 sg13g2_fill_1 FILLER_57_1602 ();
 sg13g2_fill_1 FILLER_57_1633 ();
 sg13g2_fill_2 FILLER_57_1646 ();
 sg13g2_decap_4 FILLER_57_1652 ();
 sg13g2_fill_2 FILLER_57_1656 ();
 sg13g2_fill_1 FILLER_57_1662 ();
 sg13g2_fill_2 FILLER_57_1693 ();
 sg13g2_fill_1 FILLER_57_1695 ();
 sg13g2_fill_1 FILLER_57_1740 ();
 sg13g2_decap_4 FILLER_57_1777 ();
 sg13g2_decap_4 FILLER_57_1808 ();
 sg13g2_fill_1 FILLER_57_1812 ();
 sg13g2_fill_2 FILLER_57_1914 ();
 sg13g2_fill_1 FILLER_57_1916 ();
 sg13g2_decap_8 FILLER_57_1926 ();
 sg13g2_fill_2 FILLER_57_1933 ();
 sg13g2_fill_2 FILLER_57_1990 ();
 sg13g2_fill_1 FILLER_57_2001 ();
 sg13g2_fill_1 FILLER_57_2015 ();
 sg13g2_fill_2 FILLER_57_2029 ();
 sg13g2_decap_4 FILLER_57_2057 ();
 sg13g2_fill_1 FILLER_57_2061 ();
 sg13g2_fill_1 FILLER_57_2068 ();
 sg13g2_fill_2 FILLER_57_2073 ();
 sg13g2_fill_1 FILLER_57_2075 ();
 sg13g2_fill_2 FILLER_57_2084 ();
 sg13g2_fill_1 FILLER_57_2086 ();
 sg13g2_fill_1 FILLER_57_2092 ();
 sg13g2_decap_8 FILLER_57_2142 ();
 sg13g2_fill_1 FILLER_57_2149 ();
 sg13g2_fill_1 FILLER_57_2266 ();
 sg13g2_fill_2 FILLER_57_2323 ();
 sg13g2_fill_1 FILLER_57_2325 ();
 sg13g2_fill_2 FILLER_57_2383 ();
 sg13g2_fill_1 FILLER_57_2385 ();
 sg13g2_fill_1 FILLER_57_2396 ();
 sg13g2_fill_1 FILLER_57_2420 ();
 sg13g2_fill_2 FILLER_57_2485 ();
 sg13g2_fill_1 FILLER_57_2487 ();
 sg13g2_fill_2 FILLER_57_2494 ();
 sg13g2_fill_1 FILLER_57_2496 ();
 sg13g2_fill_2 FILLER_57_2527 ();
 sg13g2_fill_1 FILLER_57_2529 ();
 sg13g2_decap_4 FILLER_57_2570 ();
 sg13g2_fill_1 FILLER_57_2574 ();
 sg13g2_fill_1 FILLER_57_2585 ();
 sg13g2_fill_2 FILLER_58_48 ();
 sg13g2_decap_4 FILLER_58_65 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_fill_1 FILLER_58_86 ();
 sg13g2_fill_1 FILLER_58_108 ();
 sg13g2_fill_1 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_150 ();
 sg13g2_fill_1 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_172 ();
 sg13g2_fill_1 FILLER_58_195 ();
 sg13g2_fill_1 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_302 ();
 sg13g2_fill_2 FILLER_58_374 ();
 sg13g2_fill_1 FILLER_58_416 ();
 sg13g2_fill_1 FILLER_58_436 ();
 sg13g2_fill_2 FILLER_58_442 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_fill_1 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_536 ();
 sg13g2_fill_1 FILLER_58_546 ();
 sg13g2_fill_2 FILLER_58_562 ();
 sg13g2_fill_1 FILLER_58_592 ();
 sg13g2_fill_2 FILLER_58_706 ();
 sg13g2_fill_1 FILLER_58_747 ();
 sg13g2_fill_1 FILLER_58_763 ();
 sg13g2_fill_1 FILLER_58_782 ();
 sg13g2_fill_1 FILLER_58_804 ();
 sg13g2_fill_2 FILLER_58_814 ();
 sg13g2_fill_1 FILLER_58_828 ();
 sg13g2_fill_2 FILLER_58_838 ();
 sg13g2_fill_1 FILLER_58_840 ();
 sg13g2_fill_2 FILLER_58_909 ();
 sg13g2_fill_1 FILLER_58_911 ();
 sg13g2_fill_1 FILLER_58_922 ();
 sg13g2_fill_1 FILLER_58_967 ();
 sg13g2_fill_2 FILLER_58_981 ();
 sg13g2_fill_1 FILLER_58_983 ();
 sg13g2_fill_1 FILLER_58_997 ();
 sg13g2_fill_2 FILLER_58_1016 ();
 sg13g2_fill_1 FILLER_58_1018 ();
 sg13g2_fill_2 FILLER_58_1102 ();
 sg13g2_fill_1 FILLER_58_1104 ();
 sg13g2_fill_1 FILLER_58_1153 ();
 sg13g2_fill_1 FILLER_58_1158 ();
 sg13g2_fill_2 FILLER_58_1251 ();
 sg13g2_fill_1 FILLER_58_1253 ();
 sg13g2_fill_2 FILLER_58_1282 ();
 sg13g2_fill_2 FILLER_58_1297 ();
 sg13g2_fill_1 FILLER_58_1299 ();
 sg13g2_fill_1 FILLER_58_1350 ();
 sg13g2_fill_1 FILLER_58_1371 ();
 sg13g2_fill_2 FILLER_58_1503 ();
 sg13g2_fill_1 FILLER_58_1505 ();
 sg13g2_fill_2 FILLER_58_1516 ();
 sg13g2_fill_1 FILLER_58_1534 ();
 sg13g2_fill_1 FILLER_58_1556 ();
 sg13g2_fill_2 FILLER_58_1570 ();
 sg13g2_fill_1 FILLER_58_1581 ();
 sg13g2_fill_1 FILLER_58_1593 ();
 sg13g2_fill_2 FILLER_58_1602 ();
 sg13g2_fill_1 FILLER_58_1604 ();
 sg13g2_fill_1 FILLER_58_1625 ();
 sg13g2_fill_2 FILLER_58_1643 ();
 sg13g2_decap_4 FILLER_58_1668 ();
 sg13g2_fill_2 FILLER_58_1672 ();
 sg13g2_fill_1 FILLER_58_1714 ();
 sg13g2_fill_2 FILLER_58_1751 ();
 sg13g2_fill_1 FILLER_58_1753 ();
 sg13g2_fill_2 FILLER_58_1789 ();
 sg13g2_fill_1 FILLER_58_1791 ();
 sg13g2_fill_1 FILLER_58_1852 ();
 sg13g2_decap_4 FILLER_58_1908 ();
 sg13g2_fill_2 FILLER_58_1912 ();
 sg13g2_fill_2 FILLER_58_1943 ();
 sg13g2_fill_1 FILLER_58_1945 ();
 sg13g2_fill_1 FILLER_58_1957 ();
 sg13g2_fill_2 FILLER_58_2010 ();
 sg13g2_fill_2 FILLER_58_2055 ();
 sg13g2_fill_2 FILLER_58_2063 ();
 sg13g2_fill_2 FILLER_58_2099 ();
 sg13g2_decap_4 FILLER_58_2128 ();
 sg13g2_fill_1 FILLER_58_2132 ();
 sg13g2_fill_1 FILLER_58_2225 ();
 sg13g2_decap_8 FILLER_58_2239 ();
 sg13g2_decap_4 FILLER_58_2246 ();
 sg13g2_decap_4 FILLER_58_2279 ();
 sg13g2_fill_2 FILLER_58_2283 ();
 sg13g2_fill_1 FILLER_58_2292 ();
 sg13g2_fill_1 FILLER_58_2314 ();
 sg13g2_fill_2 FILLER_58_2341 ();
 sg13g2_fill_2 FILLER_58_2371 ();
 sg13g2_fill_1 FILLER_58_2373 ();
 sg13g2_fill_2 FILLER_58_2415 ();
 sg13g2_fill_2 FILLER_58_2443 ();
 sg13g2_fill_2 FILLER_58_2547 ();
 sg13g2_fill_1 FILLER_58_2549 ();
 sg13g2_fill_2 FILLER_58_2571 ();
 sg13g2_fill_2 FILLER_58_2623 ();
 sg13g2_fill_1 FILLER_58_2625 ();
 sg13g2_fill_1 FILLER_58_2645 ();
 sg13g2_fill_2 FILLER_58_2672 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_4 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_19 ();
 sg13g2_fill_2 FILLER_59_66 ();
 sg13g2_fill_2 FILLER_59_73 ();
 sg13g2_fill_1 FILLER_59_75 ();
 sg13g2_fill_1 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_129 ();
 sg13g2_fill_2 FILLER_59_135 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_160 ();
 sg13g2_fill_2 FILLER_59_177 ();
 sg13g2_fill_2 FILLER_59_247 ();
 sg13g2_fill_2 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_312 ();
 sg13g2_fill_1 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_550 ();
 sg13g2_fill_1 FILLER_59_572 ();
 sg13g2_fill_1 FILLER_59_597 ();
 sg13g2_fill_2 FILLER_59_643 ();
 sg13g2_fill_2 FILLER_59_650 ();
 sg13g2_fill_2 FILLER_59_691 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_800 ();
 sg13g2_fill_1 FILLER_59_834 ();
 sg13g2_fill_2 FILLER_59_884 ();
 sg13g2_fill_1 FILLER_59_886 ();
 sg13g2_fill_1 FILLER_59_910 ();
 sg13g2_fill_1 FILLER_59_945 ();
 sg13g2_fill_2 FILLER_59_973 ();
 sg13g2_fill_1 FILLER_59_975 ();
 sg13g2_fill_1 FILLER_59_981 ();
 sg13g2_fill_2 FILLER_59_987 ();
 sg13g2_fill_1 FILLER_59_1002 ();
 sg13g2_fill_1 FILLER_59_1034 ();
 sg13g2_fill_2 FILLER_59_1063 ();
 sg13g2_fill_2 FILLER_59_1075 ();
 sg13g2_fill_1 FILLER_59_1077 ();
 sg13g2_fill_2 FILLER_59_1110 ();
 sg13g2_fill_2 FILLER_59_1122 ();
 sg13g2_fill_1 FILLER_59_1124 ();
 sg13g2_fill_1 FILLER_59_1188 ();
 sg13g2_fill_2 FILLER_59_1215 ();
 sg13g2_fill_2 FILLER_59_1225 ();
 sg13g2_fill_2 FILLER_59_1269 ();
 sg13g2_fill_1 FILLER_59_1316 ();
 sg13g2_fill_2 FILLER_59_1322 ();
 sg13g2_decap_8 FILLER_59_1336 ();
 sg13g2_decap_8 FILLER_59_1343 ();
 sg13g2_decap_4 FILLER_59_1350 ();
 sg13g2_fill_1 FILLER_59_1354 ();
 sg13g2_decap_4 FILLER_59_1364 ();
 sg13g2_fill_1 FILLER_59_1368 ();
 sg13g2_decap_4 FILLER_59_1384 ();
 sg13g2_fill_2 FILLER_59_1388 ();
 sg13g2_fill_2 FILLER_59_1432 ();
 sg13g2_fill_2 FILLER_59_1458 ();
 sg13g2_fill_1 FILLER_59_1460 ();
 sg13g2_fill_2 FILLER_59_1471 ();
 sg13g2_fill_2 FILLER_59_1482 ();
 sg13g2_fill_2 FILLER_59_1575 ();
 sg13g2_fill_1 FILLER_59_1577 ();
 sg13g2_fill_2 FILLER_59_1592 ();
 sg13g2_fill_1 FILLER_59_1594 ();
 sg13g2_fill_1 FILLER_59_1605 ();
 sg13g2_fill_1 FILLER_59_1633 ();
 sg13g2_fill_2 FILLER_59_1657 ();
 sg13g2_fill_2 FILLER_59_1679 ();
 sg13g2_fill_2 FILLER_59_1690 ();
 sg13g2_fill_2 FILLER_59_1749 ();
 sg13g2_fill_2 FILLER_59_1755 ();
 sg13g2_fill_1 FILLER_59_1810 ();
 sg13g2_fill_2 FILLER_59_1845 ();
 sg13g2_fill_2 FILLER_59_1873 ();
 sg13g2_fill_1 FILLER_59_1875 ();
 sg13g2_fill_2 FILLER_59_1892 ();
 sg13g2_fill_2 FILLER_59_1924 ();
 sg13g2_fill_2 FILLER_59_1944 ();
 sg13g2_fill_1 FILLER_59_1946 ();
 sg13g2_decap_8 FILLER_59_1962 ();
 sg13g2_fill_2 FILLER_59_1969 ();
 sg13g2_fill_2 FILLER_59_1990 ();
 sg13g2_decap_8 FILLER_59_1998 ();
 sg13g2_fill_1 FILLER_59_2005 ();
 sg13g2_fill_2 FILLER_59_2016 ();
 sg13g2_fill_1 FILLER_59_2018 ();
 sg13g2_decap_8 FILLER_59_2036 ();
 sg13g2_decap_4 FILLER_59_2043 ();
 sg13g2_fill_2 FILLER_59_2060 ();
 sg13g2_fill_1 FILLER_59_2079 ();
 sg13g2_fill_2 FILLER_59_2093 ();
 sg13g2_fill_2 FILLER_59_2175 ();
 sg13g2_fill_2 FILLER_59_2239 ();
 sg13g2_fill_2 FILLER_59_2307 ();
 sg13g2_fill_1 FILLER_59_2309 ();
 sg13g2_fill_2 FILLER_59_2350 ();
 sg13g2_fill_1 FILLER_59_2352 ();
 sg13g2_fill_2 FILLER_59_2451 ();
 sg13g2_fill_1 FILLER_59_2453 ();
 sg13g2_decap_4 FILLER_59_2569 ();
 sg13g2_fill_2 FILLER_59_2601 ();
 sg13g2_decap_4 FILLER_59_2628 ();
 sg13g2_fill_1 FILLER_59_2632 ();
 sg13g2_fill_2 FILLER_59_2672 ();
 sg13g2_decap_4 FILLER_60_45 ();
 sg13g2_fill_2 FILLER_60_49 ();
 sg13g2_fill_2 FILLER_60_57 ();
 sg13g2_fill_1 FILLER_60_59 ();
 sg13g2_fill_2 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_77 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_fill_2 FILLER_60_144 ();
 sg13g2_fill_2 FILLER_60_230 ();
 sg13g2_fill_2 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_fill_1 FILLER_60_379 ();
 sg13g2_fill_2 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_482 ();
 sg13g2_fill_2 FILLER_60_514 ();
 sg13g2_fill_1 FILLER_60_530 ();
 sg13g2_fill_1 FILLER_60_566 ();
 sg13g2_fill_2 FILLER_60_611 ();
 sg13g2_fill_1 FILLER_60_626 ();
 sg13g2_fill_1 FILLER_60_655 ();
 sg13g2_fill_2 FILLER_60_678 ();
 sg13g2_fill_2 FILLER_60_686 ();
 sg13g2_fill_1 FILLER_60_688 ();
 sg13g2_fill_2 FILLER_60_703 ();
 sg13g2_fill_2 FILLER_60_719 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_758 ();
 sg13g2_fill_1 FILLER_60_773 ();
 sg13g2_fill_2 FILLER_60_791 ();
 sg13g2_fill_1 FILLER_60_793 ();
 sg13g2_fill_2 FILLER_60_808 ();
 sg13g2_fill_1 FILLER_60_846 ();
 sg13g2_fill_1 FILLER_60_862 ();
 sg13g2_fill_1 FILLER_60_867 ();
 sg13g2_fill_1 FILLER_60_881 ();
 sg13g2_fill_2 FILLER_60_930 ();
 sg13g2_fill_1 FILLER_60_932 ();
 sg13g2_fill_2 FILLER_60_973 ();
 sg13g2_fill_1 FILLER_60_1011 ();
 sg13g2_fill_2 FILLER_60_1037 ();
 sg13g2_fill_1 FILLER_60_1116 ();
 sg13g2_fill_2 FILLER_60_1152 ();
 sg13g2_fill_2 FILLER_60_1237 ();
 sg13g2_fill_1 FILLER_60_1239 ();
 sg13g2_fill_1 FILLER_60_1245 ();
 sg13g2_decap_4 FILLER_60_1258 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_fill_2 FILLER_60_1302 ();
 sg13g2_fill_2 FILLER_60_1328 ();
 sg13g2_fill_2 FILLER_60_1375 ();
 sg13g2_fill_1 FILLER_60_1377 ();
 sg13g2_fill_2 FILLER_60_1412 ();
 sg13g2_fill_1 FILLER_60_1414 ();
 sg13g2_fill_2 FILLER_60_1420 ();
 sg13g2_fill_2 FILLER_60_1430 ();
 sg13g2_fill_1 FILLER_60_1432 ();
 sg13g2_fill_2 FILLER_60_1467 ();
 sg13g2_fill_1 FILLER_60_1477 ();
 sg13g2_fill_1 FILLER_60_1495 ();
 sg13g2_fill_1 FILLER_60_1505 ();
 sg13g2_fill_2 FILLER_60_1510 ();
 sg13g2_fill_1 FILLER_60_1512 ();
 sg13g2_fill_2 FILLER_60_1543 ();
 sg13g2_fill_1 FILLER_60_1545 ();
 sg13g2_fill_2 FILLER_60_1571 ();
 sg13g2_fill_2 FILLER_60_1589 ();
 sg13g2_fill_1 FILLER_60_1615 ();
 sg13g2_fill_1 FILLER_60_1635 ();
 sg13g2_fill_1 FILLER_60_1650 ();
 sg13g2_decap_4 FILLER_60_1657 ();
 sg13g2_fill_2 FILLER_60_1661 ();
 sg13g2_fill_2 FILLER_60_1667 ();
 sg13g2_fill_1 FILLER_60_1669 ();
 sg13g2_decap_4 FILLER_60_1771 ();
 sg13g2_fill_2 FILLER_60_1775 ();
 sg13g2_fill_2 FILLER_60_1813 ();
 sg13g2_fill_1 FILLER_60_1815 ();
 sg13g2_fill_2 FILLER_60_1829 ();
 sg13g2_fill_2 FILLER_60_1908 ();
 sg13g2_fill_1 FILLER_60_1910 ();
 sg13g2_fill_2 FILLER_60_1926 ();
 sg13g2_fill_2 FILLER_60_1934 ();
 sg13g2_fill_1 FILLER_60_1936 ();
 sg13g2_fill_2 FILLER_60_1946 ();
 sg13g2_fill_1 FILLER_60_1948 ();
 sg13g2_fill_2 FILLER_60_1963 ();
 sg13g2_fill_1 FILLER_60_1965 ();
 sg13g2_decap_4 FILLER_60_1970 ();
 sg13g2_fill_2 FILLER_60_1979 ();
 sg13g2_fill_1 FILLER_60_1981 ();
 sg13g2_fill_2 FILLER_60_1987 ();
 sg13g2_fill_1 FILLER_60_1989 ();
 sg13g2_fill_1 FILLER_60_2011 ();
 sg13g2_fill_1 FILLER_60_2061 ();
 sg13g2_decap_8 FILLER_60_2072 ();
 sg13g2_decap_4 FILLER_60_2079 ();
 sg13g2_fill_2 FILLER_60_2083 ();
 sg13g2_decap_8 FILLER_60_2094 ();
 sg13g2_fill_1 FILLER_60_2101 ();
 sg13g2_fill_2 FILLER_60_2151 ();
 sg13g2_fill_1 FILLER_60_2153 ();
 sg13g2_fill_2 FILLER_60_2210 ();
 sg13g2_fill_1 FILLER_60_2212 ();
 sg13g2_fill_1 FILLER_60_2237 ();
 sg13g2_fill_1 FILLER_60_2248 ();
 sg13g2_decap_8 FILLER_60_2320 ();
 sg13g2_fill_2 FILLER_60_2327 ();
 sg13g2_fill_1 FILLER_60_2329 ();
 sg13g2_fill_2 FILLER_60_2344 ();
 sg13g2_fill_2 FILLER_60_2392 ();
 sg13g2_fill_1 FILLER_60_2404 ();
 sg13g2_fill_2 FILLER_60_2438 ();
 sg13g2_fill_1 FILLER_60_2452 ();
 sg13g2_fill_2 FILLER_60_2498 ();
 sg13g2_fill_1 FILLER_60_2500 ();
 sg13g2_fill_2 FILLER_60_2518 ();
 sg13g2_fill_2 FILLER_60_2530 ();
 sg13g2_fill_1 FILLER_60_2532 ();
 sg13g2_fill_1 FILLER_60_2537 ();
 sg13g2_fill_1 FILLER_60_2547 ();
 sg13g2_fill_2 FILLER_60_2558 ();
 sg13g2_fill_1 FILLER_60_2560 ();
 sg13g2_fill_2 FILLER_60_2671 ();
 sg13g2_fill_1 FILLER_60_2673 ();
 sg13g2_fill_2 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_86 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_decap_4 FILLER_61_111 ();
 sg13g2_fill_1 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_160 ();
 sg13g2_fill_2 FILLER_61_208 ();
 sg13g2_fill_1 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_251 ();
 sg13g2_fill_1 FILLER_61_261 ();
 sg13g2_fill_1 FILLER_61_310 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_fill_2 FILLER_61_642 ();
 sg13g2_fill_1 FILLER_61_644 ();
 sg13g2_fill_2 FILLER_61_658 ();
 sg13g2_fill_2 FILLER_61_686 ();
 sg13g2_fill_1 FILLER_61_688 ();
 sg13g2_fill_2 FILLER_61_729 ();
 sg13g2_fill_1 FILLER_61_731 ();
 sg13g2_fill_1 FILLER_61_736 ();
 sg13g2_fill_1 FILLER_61_750 ();
 sg13g2_fill_2 FILLER_61_807 ();
 sg13g2_fill_1 FILLER_61_835 ();
 sg13g2_fill_2 FILLER_61_871 ();
 sg13g2_fill_2 FILLER_61_886 ();
 sg13g2_fill_1 FILLER_61_888 ();
 sg13g2_fill_1 FILLER_61_893 ();
 sg13g2_fill_1 FILLER_61_942 ();
 sg13g2_fill_1 FILLER_61_974 ();
 sg13g2_fill_1 FILLER_61_1042 ();
 sg13g2_fill_2 FILLER_61_1049 ();
 sg13g2_fill_1 FILLER_61_1051 ();
 sg13g2_fill_1 FILLER_61_1066 ();
 sg13g2_fill_2 FILLER_61_1101 ();
 sg13g2_fill_2 FILLER_61_1166 ();
 sg13g2_fill_2 FILLER_61_1183 ();
 sg13g2_fill_1 FILLER_61_1185 ();
 sg13g2_fill_2 FILLER_61_1204 ();
 sg13g2_fill_1 FILLER_61_1206 ();
 sg13g2_fill_2 FILLER_61_1247 ();
 sg13g2_fill_1 FILLER_61_1275 ();
 sg13g2_fill_1 FILLER_61_1301 ();
 sg13g2_fill_1 FILLER_61_1305 ();
 sg13g2_fill_2 FILLER_61_1319 ();
 sg13g2_decap_8 FILLER_61_1342 ();
 sg13g2_fill_2 FILLER_61_1349 ();
 sg13g2_decap_4 FILLER_61_1356 ();
 sg13g2_fill_2 FILLER_61_1360 ();
 sg13g2_fill_1 FILLER_61_1367 ();
 sg13g2_fill_1 FILLER_61_1373 ();
 sg13g2_decap_4 FILLER_61_1382 ();
 sg13g2_fill_2 FILLER_61_1391 ();
 sg13g2_decap_4 FILLER_61_1401 ();
 sg13g2_fill_1 FILLER_61_1405 ();
 sg13g2_fill_2 FILLER_61_1436 ();
 sg13g2_fill_1 FILLER_61_1447 ();
 sg13g2_fill_1 FILLER_61_1554 ();
 sg13g2_fill_1 FILLER_61_1567 ();
 sg13g2_fill_2 FILLER_61_1593 ();
 sg13g2_fill_1 FILLER_61_1595 ();
 sg13g2_fill_2 FILLER_61_1601 ();
 sg13g2_fill_2 FILLER_61_1607 ();
 sg13g2_decap_4 FILLER_61_1619 ();
 sg13g2_fill_1 FILLER_61_1623 ();
 sg13g2_decap_8 FILLER_61_1629 ();
 sg13g2_decap_8 FILLER_61_1655 ();
 sg13g2_fill_2 FILLER_61_1662 ();
 sg13g2_fill_1 FILLER_61_1664 ();
 sg13g2_fill_2 FILLER_61_1672 ();
 sg13g2_fill_2 FILLER_61_1690 ();
 sg13g2_fill_2 FILLER_61_1709 ();
 sg13g2_fill_2 FILLER_61_1732 ();
 sg13g2_fill_2 FILLER_61_1742 ();
 sg13g2_fill_1 FILLER_61_1744 ();
 sg13g2_decap_4 FILLER_61_1750 ();
 sg13g2_fill_2 FILLER_61_1791 ();
 sg13g2_decap_4 FILLER_61_1899 ();
 sg13g2_fill_1 FILLER_61_1903 ();
 sg13g2_decap_4 FILLER_61_1924 ();
 sg13g2_fill_2 FILLER_61_1932 ();
 sg13g2_fill_2 FILLER_61_1996 ();
 sg13g2_fill_1 FILLER_61_1998 ();
 sg13g2_decap_4 FILLER_61_2006 ();
 sg13g2_decap_8 FILLER_61_2021 ();
 sg13g2_fill_1 FILLER_61_2028 ();
 sg13g2_fill_2 FILLER_61_2039 ();
 sg13g2_fill_1 FILLER_61_2041 ();
 sg13g2_fill_2 FILLER_61_2064 ();
 sg13g2_fill_1 FILLER_61_2066 ();
 sg13g2_fill_2 FILLER_61_2074 ();
 sg13g2_decap_8 FILLER_61_2084 ();
 sg13g2_fill_2 FILLER_61_2091 ();
 sg13g2_fill_2 FILLER_61_2187 ();
 sg13g2_fill_2 FILLER_61_2215 ();
 sg13g2_fill_2 FILLER_61_2247 ();
 sg13g2_fill_1 FILLER_61_2249 ();
 sg13g2_fill_2 FILLER_61_2255 ();
 sg13g2_decap_8 FILLER_61_2269 ();
 sg13g2_fill_2 FILLER_61_2352 ();
 sg13g2_fill_1 FILLER_61_2354 ();
 sg13g2_decap_4 FILLER_61_2391 ();
 sg13g2_fill_2 FILLER_61_2421 ();
 sg13g2_fill_2 FILLER_61_2449 ();
 sg13g2_fill_1 FILLER_61_2451 ();
 sg13g2_fill_2 FILLER_61_2552 ();
 sg13g2_fill_1 FILLER_61_2554 ();
 sg13g2_fill_1 FILLER_61_2598 ();
 sg13g2_fill_2 FILLER_61_2609 ();
 sg13g2_fill_1 FILLER_61_2631 ();
 sg13g2_fill_1 FILLER_61_2641 ();
 sg13g2_decap_4 FILLER_61_2655 ();
 sg13g2_decap_8 FILLER_61_2663 ();
 sg13g2_decap_4 FILLER_61_2670 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_33 ();
 sg13g2_fill_1 FILLER_62_51 ();
 sg13g2_fill_1 FILLER_62_60 ();
 sg13g2_fill_2 FILLER_62_69 ();
 sg13g2_fill_2 FILLER_62_115 ();
 sg13g2_fill_1 FILLER_62_117 ();
 sg13g2_fill_1 FILLER_62_149 ();
 sg13g2_fill_1 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_298 ();
 sg13g2_fill_1 FILLER_62_338 ();
 sg13g2_fill_2 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_448 ();
 sg13g2_fill_1 FILLER_62_491 ();
 sg13g2_fill_2 FILLER_62_592 ();
 sg13g2_fill_2 FILLER_62_630 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_fill_2 FILLER_62_691 ();
 sg13g2_fill_2 FILLER_62_709 ();
 sg13g2_fill_2 FILLER_62_760 ();
 sg13g2_fill_2 FILLER_62_772 ();
 sg13g2_fill_2 FILLER_62_830 ();
 sg13g2_fill_1 FILLER_62_876 ();
 sg13g2_fill_2 FILLER_62_903 ();
 sg13g2_fill_2 FILLER_62_919 ();
 sg13g2_fill_2 FILLER_62_940 ();
 sg13g2_fill_1 FILLER_62_946 ();
 sg13g2_fill_2 FILLER_62_1011 ();
 sg13g2_fill_2 FILLER_62_1079 ();
 sg13g2_fill_1 FILLER_62_1081 ();
 sg13g2_fill_2 FILLER_62_1091 ();
 sg13g2_fill_2 FILLER_62_1110 ();
 sg13g2_fill_1 FILLER_62_1112 ();
 sg13g2_fill_1 FILLER_62_1138 ();
 sg13g2_fill_2 FILLER_62_1157 ();
 sg13g2_fill_1 FILLER_62_1211 ();
 sg13g2_fill_2 FILLER_62_1240 ();
 sg13g2_fill_1 FILLER_62_1247 ();
 sg13g2_decap_8 FILLER_62_1263 ();
 sg13g2_fill_1 FILLER_62_1281 ();
 sg13g2_fill_2 FILLER_62_1295 ();
 sg13g2_fill_1 FILLER_62_1297 ();
 sg13g2_fill_1 FILLER_62_1315 ();
 sg13g2_fill_1 FILLER_62_1320 ();
 sg13g2_decap_4 FILLER_62_1343 ();
 sg13g2_fill_1 FILLER_62_1347 ();
 sg13g2_fill_2 FILLER_62_1356 ();
 sg13g2_fill_2 FILLER_62_1366 ();
 sg13g2_fill_2 FILLER_62_1384 ();
 sg13g2_fill_1 FILLER_62_1399 ();
 sg13g2_fill_1 FILLER_62_1434 ();
 sg13g2_fill_2 FILLER_62_1454 ();
 sg13g2_fill_1 FILLER_62_1472 ();
 sg13g2_fill_2 FILLER_62_1487 ();
 sg13g2_fill_1 FILLER_62_1489 ();
 sg13g2_fill_1 FILLER_62_1495 ();
 sg13g2_fill_1 FILLER_62_1505 ();
 sg13g2_fill_2 FILLER_62_1569 ();
 sg13g2_fill_1 FILLER_62_1571 ();
 sg13g2_fill_1 FILLER_62_1577 ();
 sg13g2_fill_2 FILLER_62_1650 ();
 sg13g2_fill_2 FILLER_62_1660 ();
 sg13g2_fill_1 FILLER_62_1662 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_fill_2 FILLER_62_1686 ();
 sg13g2_fill_2 FILLER_62_1724 ();
 sg13g2_fill_1 FILLER_62_1814 ();
 sg13g2_fill_2 FILLER_62_1850 ();
 sg13g2_decap_8 FILLER_62_1897 ();
 sg13g2_fill_2 FILLER_62_1904 ();
 sg13g2_fill_1 FILLER_62_1906 ();
 sg13g2_decap_4 FILLER_62_1912 ();
 sg13g2_fill_2 FILLER_62_1916 ();
 sg13g2_decap_4 FILLER_62_1943 ();
 sg13g2_decap_4 FILLER_62_1966 ();
 sg13g2_fill_1 FILLER_62_1986 ();
 sg13g2_decap_4 FILLER_62_2001 ();
 sg13g2_fill_1 FILLER_62_2020 ();
 sg13g2_decap_8 FILLER_62_2036 ();
 sg13g2_fill_1 FILLER_62_2043 ();
 sg13g2_decap_4 FILLER_62_2052 ();
 sg13g2_decap_4 FILLER_62_2099 ();
 sg13g2_fill_1 FILLER_62_2103 ();
 sg13g2_fill_2 FILLER_62_2108 ();
 sg13g2_fill_1 FILLER_62_2110 ();
 sg13g2_fill_2 FILLER_62_2172 ();
 sg13g2_fill_1 FILLER_62_2174 ();
 sg13g2_fill_1 FILLER_62_2183 ();
 sg13g2_fill_2 FILLER_62_2240 ();
 sg13g2_fill_2 FILLER_62_2349 ();
 sg13g2_fill_1 FILLER_62_2387 ();
 sg13g2_fill_2 FILLER_62_2410 ();
 sg13g2_fill_2 FILLER_62_2437 ();
 sg13g2_fill_1 FILLER_62_2439 ();
 sg13g2_fill_2 FILLER_62_2466 ();
 sg13g2_fill_2 FILLER_62_2504 ();
 sg13g2_fill_2 FILLER_62_2563 ();
 sg13g2_fill_1 FILLER_62_2565 ();
 sg13g2_fill_1 FILLER_62_2605 ();
 sg13g2_decap_8 FILLER_62_2662 ();
 sg13g2_decap_4 FILLER_62_2669 ();
 sg13g2_fill_1 FILLER_62_2673 ();
 sg13g2_fill_2 FILLER_63_62 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_fill_1 FILLER_63_102 ();
 sg13g2_fill_2 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_fill_1 FILLER_63_174 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_369 ();
 sg13g2_fill_2 FILLER_63_386 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_2 FILLER_63_442 ();
 sg13g2_fill_2 FILLER_63_462 ();
 sg13g2_fill_2 FILLER_63_616 ();
 sg13g2_fill_2 FILLER_63_632 ();
 sg13g2_fill_1 FILLER_63_634 ();
 sg13g2_fill_2 FILLER_63_640 ();
 sg13g2_fill_1 FILLER_63_642 ();
 sg13g2_fill_2 FILLER_63_648 ();
 sg13g2_fill_1 FILLER_63_650 ();
 sg13g2_fill_2 FILLER_63_660 ();
 sg13g2_fill_2 FILLER_63_694 ();
 sg13g2_fill_1 FILLER_63_696 ();
 sg13g2_fill_2 FILLER_63_738 ();
 sg13g2_fill_1 FILLER_63_740 ();
 sg13g2_fill_2 FILLER_63_785 ();
 sg13g2_fill_2 FILLER_63_805 ();
 sg13g2_fill_2 FILLER_63_824 ();
 sg13g2_fill_1 FILLER_63_826 ();
 sg13g2_fill_2 FILLER_63_868 ();
 sg13g2_fill_1 FILLER_63_883 ();
 sg13g2_fill_1 FILLER_63_921 ();
 sg13g2_fill_1 FILLER_63_957 ();
 sg13g2_fill_2 FILLER_63_969 ();
 sg13g2_fill_1 FILLER_63_971 ();
 sg13g2_fill_1 FILLER_63_981 ();
 sg13g2_fill_2 FILLER_63_1035 ();
 sg13g2_fill_1 FILLER_63_1091 ();
 sg13g2_fill_2 FILLER_63_1172 ();
 sg13g2_fill_2 FILLER_63_1209 ();
 sg13g2_fill_1 FILLER_63_1211 ();
 sg13g2_fill_2 FILLER_63_1231 ();
 sg13g2_fill_1 FILLER_63_1233 ();
 sg13g2_fill_1 FILLER_63_1286 ();
 sg13g2_decap_8 FILLER_63_1294 ();
 sg13g2_fill_1 FILLER_63_1301 ();
 sg13g2_fill_2 FILLER_63_1310 ();
 sg13g2_fill_1 FILLER_63_1312 ();
 sg13g2_fill_1 FILLER_63_1327 ();
 sg13g2_fill_1 FILLER_63_1333 ();
 sg13g2_decap_4 FILLER_63_1339 ();
 sg13g2_fill_1 FILLER_63_1358 ();
 sg13g2_fill_1 FILLER_63_1368 ();
 sg13g2_fill_2 FILLER_63_1390 ();
 sg13g2_fill_2 FILLER_63_1401 ();
 sg13g2_fill_1 FILLER_63_1403 ();
 sg13g2_fill_2 FILLER_63_1408 ();
 sg13g2_fill_1 FILLER_63_1410 ();
 sg13g2_fill_2 FILLER_63_1438 ();
 sg13g2_fill_2 FILLER_63_1445 ();
 sg13g2_fill_1 FILLER_63_1447 ();
 sg13g2_fill_1 FILLER_63_1453 ();
 sg13g2_fill_2 FILLER_63_1485 ();
 sg13g2_fill_2 FILLER_63_1495 ();
 sg13g2_fill_2 FILLER_63_1570 ();
 sg13g2_decap_4 FILLER_63_1593 ();
 sg13g2_fill_2 FILLER_63_1597 ();
 sg13g2_decap_4 FILLER_63_1616 ();
 sg13g2_fill_1 FILLER_63_1620 ();
 sg13g2_fill_2 FILLER_63_1626 ();
 sg13g2_fill_1 FILLER_63_1628 ();
 sg13g2_fill_1 FILLER_63_1641 ();
 sg13g2_fill_2 FILLER_63_1692 ();
 sg13g2_fill_1 FILLER_63_1694 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_fill_2 FILLER_63_1813 ();
 sg13g2_fill_2 FILLER_63_1841 ();
 sg13g2_fill_1 FILLER_63_1843 ();
 sg13g2_fill_2 FILLER_63_1874 ();
 sg13g2_fill_1 FILLER_63_1876 ();
 sg13g2_fill_1 FILLER_63_1907 ();
 sg13g2_decap_4 FILLER_63_1948 ();
 sg13g2_fill_1 FILLER_63_1956 ();
 sg13g2_fill_1 FILLER_63_1966 ();
 sg13g2_decap_4 FILLER_63_1977 ();
 sg13g2_fill_2 FILLER_63_2005 ();
 sg13g2_fill_1 FILLER_63_2007 ();
 sg13g2_decap_8 FILLER_63_2018 ();
 sg13g2_decap_4 FILLER_63_2029 ();
 sg13g2_fill_2 FILLER_63_2060 ();
 sg13g2_fill_2 FILLER_63_2066 ();
 sg13g2_fill_1 FILLER_63_2078 ();
 sg13g2_fill_1 FILLER_63_2096 ();
 sg13g2_decap_4 FILLER_63_2133 ();
 sg13g2_fill_1 FILLER_63_2137 ();
 sg13g2_fill_1 FILLER_63_2224 ();
 sg13g2_fill_2 FILLER_63_2235 ();
 sg13g2_fill_1 FILLER_63_2247 ();
 sg13g2_fill_2 FILLER_63_2275 ();
 sg13g2_fill_1 FILLER_63_2277 ();
 sg13g2_decap_4 FILLER_63_2282 ();
 sg13g2_fill_2 FILLER_63_2328 ();
 sg13g2_decap_4 FILLER_63_2370 ();
 sg13g2_fill_2 FILLER_63_2374 ();
 sg13g2_decap_8 FILLER_63_2384 ();
 sg13g2_fill_2 FILLER_63_2391 ();
 sg13g2_fill_1 FILLER_63_2393 ();
 sg13g2_fill_1 FILLER_63_2425 ();
 sg13g2_fill_2 FILLER_63_2452 ();
 sg13g2_fill_2 FILLER_63_2494 ();
 sg13g2_fill_1 FILLER_63_2496 ();
 sg13g2_fill_2 FILLER_63_2516 ();
 sg13g2_fill_1 FILLER_63_2518 ();
 sg13g2_fill_2 FILLER_63_2542 ();
 sg13g2_fill_2 FILLER_63_2590 ();
 sg13g2_fill_1 FILLER_63_2592 ();
 sg13g2_fill_2 FILLER_63_2623 ();
 sg13g2_decap_4 FILLER_63_2639 ();
 sg13g2_fill_2 FILLER_63_2643 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_decap_4 FILLER_63_2669 ();
 sg13g2_fill_1 FILLER_63_2673 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_15 ();
 sg13g2_fill_2 FILLER_64_34 ();
 sg13g2_fill_1 FILLER_64_111 ();
 sg13g2_fill_2 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_132 ();
 sg13g2_fill_1 FILLER_64_226 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_244 ();
 sg13g2_fill_2 FILLER_64_258 ();
 sg13g2_fill_2 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_490 ();
 sg13g2_fill_1 FILLER_64_526 ();
 sg13g2_fill_1 FILLER_64_542 ();
 sg13g2_fill_2 FILLER_64_577 ();
 sg13g2_fill_1 FILLER_64_593 ();
 sg13g2_fill_2 FILLER_64_630 ();
 sg13g2_fill_1 FILLER_64_632 ();
 sg13g2_fill_1 FILLER_64_644 ();
 sg13g2_fill_2 FILLER_64_676 ();
 sg13g2_fill_1 FILLER_64_678 ();
 sg13g2_fill_1 FILLER_64_717 ();
 sg13g2_fill_1 FILLER_64_753 ();
 sg13g2_fill_1 FILLER_64_799 ();
 sg13g2_fill_2 FILLER_64_826 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_fill_2 FILLER_64_899 ();
 sg13g2_fill_2 FILLER_64_927 ();
 sg13g2_fill_2 FILLER_64_953 ();
 sg13g2_fill_1 FILLER_64_955 ();
 sg13g2_fill_2 FILLER_64_984 ();
 sg13g2_fill_1 FILLER_64_986 ();
 sg13g2_fill_2 FILLER_64_1001 ();
 sg13g2_fill_1 FILLER_64_1061 ();
 sg13g2_fill_2 FILLER_64_1103 ();
 sg13g2_fill_1 FILLER_64_1105 ();
 sg13g2_fill_1 FILLER_64_1142 ();
 sg13g2_fill_2 FILLER_64_1182 ();
 sg13g2_fill_2 FILLER_64_1189 ();
 sg13g2_fill_1 FILLER_64_1191 ();
 sg13g2_fill_1 FILLER_64_1258 ();
 sg13g2_fill_2 FILLER_64_1275 ();
 sg13g2_fill_1 FILLER_64_1277 ();
 sg13g2_fill_2 FILLER_64_1286 ();
 sg13g2_fill_1 FILLER_64_1288 ();
 sg13g2_decap_8 FILLER_64_1302 ();
 sg13g2_decap_4 FILLER_64_1309 ();
 sg13g2_decap_4 FILLER_64_1335 ();
 sg13g2_fill_1 FILLER_64_1339 ();
 sg13g2_fill_2 FILLER_64_1392 ();
 sg13g2_fill_1 FILLER_64_1394 ();
 sg13g2_fill_2 FILLER_64_1457 ();
 sg13g2_fill_2 FILLER_64_1464 ();
 sg13g2_fill_2 FILLER_64_1471 ();
 sg13g2_fill_1 FILLER_64_1473 ();
 sg13g2_fill_2 FILLER_64_1491 ();
 sg13g2_fill_1 FILLER_64_1493 ();
 sg13g2_fill_1 FILLER_64_1499 ();
 sg13g2_fill_2 FILLER_64_1509 ();
 sg13g2_fill_1 FILLER_64_1511 ();
 sg13g2_fill_1 FILLER_64_1529 ();
 sg13g2_fill_1 FILLER_64_1543 ();
 sg13g2_fill_1 FILLER_64_1562 ();
 sg13g2_decap_8 FILLER_64_1584 ();
 sg13g2_decap_4 FILLER_64_1603 ();
 sg13g2_fill_1 FILLER_64_1607 ();
 sg13g2_fill_2 FILLER_64_1612 ();
 sg13g2_fill_2 FILLER_64_1619 ();
 sg13g2_fill_1 FILLER_64_1621 ();
 sg13g2_decap_4 FILLER_64_1634 ();
 sg13g2_fill_2 FILLER_64_1638 ();
 sg13g2_fill_2 FILLER_64_1653 ();
 sg13g2_fill_1 FILLER_64_1655 ();
 sg13g2_fill_1 FILLER_64_1678 ();
 sg13g2_decap_4 FILLER_64_1687 ();
 sg13g2_fill_2 FILLER_64_1741 ();
 sg13g2_fill_1 FILLER_64_1743 ();
 sg13g2_fill_2 FILLER_64_1780 ();
 sg13g2_fill_2 FILLER_64_1827 ();
 sg13g2_fill_1 FILLER_64_1829 ();
 sg13g2_fill_2 FILLER_64_1866 ();
 sg13g2_fill_1 FILLER_64_1868 ();
 sg13g2_fill_2 FILLER_64_1905 ();
 sg13g2_fill_2 FILLER_64_1932 ();
 sg13g2_fill_2 FILLER_64_1938 ();
 sg13g2_fill_2 FILLER_64_1945 ();
 sg13g2_fill_2 FILLER_64_1956 ();
 sg13g2_fill_1 FILLER_64_1958 ();
 sg13g2_fill_2 FILLER_64_1973 ();
 sg13g2_fill_1 FILLER_64_1975 ();
 sg13g2_fill_1 FILLER_64_2003 ();
 sg13g2_fill_1 FILLER_64_2008 ();
 sg13g2_fill_2 FILLER_64_2016 ();
 sg13g2_fill_1 FILLER_64_2018 ();
 sg13g2_fill_2 FILLER_64_2037 ();
 sg13g2_fill_1 FILLER_64_2039 ();
 sg13g2_decap_8 FILLER_64_2050 ();
 sg13g2_fill_2 FILLER_64_2057 ();
 sg13g2_fill_1 FILLER_64_2064 ();
 sg13g2_fill_2 FILLER_64_2070 ();
 sg13g2_fill_2 FILLER_64_2081 ();
 sg13g2_fill_1 FILLER_64_2088 ();
 sg13g2_decap_4 FILLER_64_2094 ();
 sg13g2_fill_1 FILLER_64_2098 ();
 sg13g2_decap_4 FILLER_64_2134 ();
 sg13g2_decap_4 FILLER_64_2155 ();
 sg13g2_fill_2 FILLER_64_2172 ();
 sg13g2_fill_1 FILLER_64_2174 ();
 sg13g2_fill_2 FILLER_64_2194 ();
 sg13g2_fill_1 FILLER_64_2196 ();
 sg13g2_fill_2 FILLER_64_2287 ();
 sg13g2_fill_2 FILLER_64_2348 ();
 sg13g2_fill_2 FILLER_64_2399 ();
 sg13g2_fill_1 FILLER_64_2418 ();
 sg13g2_fill_2 FILLER_64_2438 ();
 sg13g2_fill_1 FILLER_64_2440 ();
 sg13g2_fill_1 FILLER_64_2545 ();
 sg13g2_decap_8 FILLER_64_2573 ();
 sg13g2_fill_2 FILLER_64_2580 ();
 sg13g2_fill_1 FILLER_64_2582 ();
 sg13g2_fill_1 FILLER_64_2632 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_8 FILLER_64_2666 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_1 FILLER_65_25 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_fill_2 FILLER_65_184 ();
 sg13g2_fill_2 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_291 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_fill_1 FILLER_65_314 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_2 FILLER_65_357 ();
 sg13g2_fill_2 FILLER_65_383 ();
 sg13g2_fill_2 FILLER_65_434 ();
 sg13g2_fill_2 FILLER_65_527 ();
 sg13g2_fill_1 FILLER_65_538 ();
 sg13g2_fill_1 FILLER_65_564 ();
 sg13g2_fill_2 FILLER_65_623 ();
 sg13g2_fill_1 FILLER_65_625 ();
 sg13g2_fill_1 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_645 ();
 sg13g2_fill_2 FILLER_65_651 ();
 sg13g2_fill_1 FILLER_65_653 ();
 sg13g2_fill_2 FILLER_65_667 ();
 sg13g2_fill_1 FILLER_65_681 ();
 sg13g2_fill_2 FILLER_65_687 ();
 sg13g2_fill_1 FILLER_65_689 ();
 sg13g2_fill_1 FILLER_65_750 ();
 sg13g2_fill_2 FILLER_65_843 ();
 sg13g2_fill_2 FILLER_65_860 ();
 sg13g2_fill_2 FILLER_65_875 ();
 sg13g2_fill_1 FILLER_65_882 ();
 sg13g2_fill_2 FILLER_65_934 ();
 sg13g2_fill_1 FILLER_65_966 ();
 sg13g2_fill_2 FILLER_65_979 ();
 sg13g2_fill_2 FILLER_65_985 ();
 sg13g2_fill_1 FILLER_65_987 ();
 sg13g2_fill_2 FILLER_65_1034 ();
 sg13g2_fill_2 FILLER_65_1118 ();
 sg13g2_fill_2 FILLER_65_1172 ();
 sg13g2_fill_1 FILLER_65_1174 ();
 sg13g2_fill_2 FILLER_65_1181 ();
 sg13g2_fill_2 FILLER_65_1188 ();
 sg13g2_fill_1 FILLER_65_1239 ();
 sg13g2_fill_2 FILLER_65_1289 ();
 sg13g2_fill_1 FILLER_65_1295 ();
 sg13g2_fill_2 FILLER_65_1308 ();
 sg13g2_fill_1 FILLER_65_1314 ();
 sg13g2_fill_1 FILLER_65_1321 ();
 sg13g2_fill_2 FILLER_65_1333 ();
 sg13g2_fill_1 FILLER_65_1335 ();
 sg13g2_fill_2 FILLER_65_1351 ();
 sg13g2_fill_2 FILLER_65_1358 ();
 sg13g2_fill_1 FILLER_65_1360 ();
 sg13g2_decap_4 FILLER_65_1366 ();
 sg13g2_fill_1 FILLER_65_1370 ();
 sg13g2_fill_1 FILLER_65_1381 ();
 sg13g2_decap_4 FILLER_65_1387 ();
 sg13g2_fill_1 FILLER_65_1426 ();
 sg13g2_fill_1 FILLER_65_1458 ();
 sg13g2_fill_1 FILLER_65_1507 ();
 sg13g2_fill_2 FILLER_65_1564 ();
 sg13g2_decap_4 FILLER_65_1580 ();
 sg13g2_fill_1 FILLER_65_1584 ();
 sg13g2_fill_2 FILLER_65_1597 ();
 sg13g2_fill_1 FILLER_65_1599 ();
 sg13g2_fill_1 FILLER_65_1645 ();
 sg13g2_fill_1 FILLER_65_1679 ();
 sg13g2_decap_8 FILLER_65_1688 ();
 sg13g2_fill_2 FILLER_65_1758 ();
 sg13g2_decap_4 FILLER_65_1777 ();
 sg13g2_fill_1 FILLER_65_1781 ();
 sg13g2_fill_1 FILLER_65_1791 ();
 sg13g2_fill_1 FILLER_65_1806 ();
 sg13g2_fill_2 FILLER_65_1828 ();
 sg13g2_fill_1 FILLER_65_1850 ();
 sg13g2_fill_2 FILLER_65_1855 ();
 sg13g2_decap_8 FILLER_65_1904 ();
 sg13g2_fill_1 FILLER_65_1911 ();
 sg13g2_fill_2 FILLER_65_1917 ();
 sg13g2_fill_2 FILLER_65_1936 ();
 sg13g2_fill_2 FILLER_65_1943 ();
 sg13g2_fill_2 FILLER_65_1952 ();
 sg13g2_fill_1 FILLER_65_1982 ();
 sg13g2_fill_1 FILLER_65_1989 ();
 sg13g2_fill_1 FILLER_65_2013 ();
 sg13g2_fill_2 FILLER_65_2049 ();
 sg13g2_fill_2 FILLER_65_2072 ();
 sg13g2_fill_1 FILLER_65_2074 ();
 sg13g2_fill_2 FILLER_65_2083 ();
 sg13g2_fill_1 FILLER_65_2085 ();
 sg13g2_decap_4 FILLER_65_2098 ();
 sg13g2_fill_2 FILLER_65_2102 ();
 sg13g2_fill_2 FILLER_65_2165 ();
 sg13g2_fill_2 FILLER_65_2237 ();
 sg13g2_fill_1 FILLER_65_2239 ();
 sg13g2_fill_2 FILLER_65_2282 ();
 sg13g2_fill_1 FILLER_65_2284 ();
 sg13g2_fill_1 FILLER_65_2306 ();
 sg13g2_fill_2 FILLER_65_2323 ();
 sg13g2_fill_1 FILLER_65_2325 ();
 sg13g2_decap_8 FILLER_65_2374 ();
 sg13g2_fill_1 FILLER_65_2381 ();
 sg13g2_fill_2 FILLER_65_2417 ();
 sg13g2_fill_1 FILLER_65_2419 ();
 sg13g2_fill_2 FILLER_65_2472 ();
 sg13g2_fill_1 FILLER_65_2518 ();
 sg13g2_decap_4 FILLER_65_2580 ();
 sg13g2_fill_1 FILLER_65_2584 ();
 sg13g2_fill_2 FILLER_65_2611 ();
 sg13g2_fill_1 FILLER_65_2613 ();
 sg13g2_decap_8 FILLER_65_2663 ();
 sg13g2_decap_4 FILLER_65_2670 ();
 sg13g2_fill_2 FILLER_66_160 ();
 sg13g2_fill_1 FILLER_66_253 ();
 sg13g2_fill_2 FILLER_66_259 ();
 sg13g2_fill_1 FILLER_66_266 ();
 sg13g2_fill_1 FILLER_66_277 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_354 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_fill_1 FILLER_66_404 ();
 sg13g2_fill_2 FILLER_66_414 ();
 sg13g2_fill_1 FILLER_66_482 ();
 sg13g2_fill_2 FILLER_66_492 ();
 sg13g2_fill_1 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_2 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_791 ();
 sg13g2_fill_2 FILLER_66_832 ();
 sg13g2_fill_1 FILLER_66_899 ();
 sg13g2_fill_2 FILLER_66_918 ();
 sg13g2_fill_2 FILLER_66_943 ();
 sg13g2_fill_1 FILLER_66_962 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_fill_2 FILLER_66_1002 ();
 sg13g2_fill_1 FILLER_66_1004 ();
 sg13g2_fill_1 FILLER_66_1017 ();
 sg13g2_fill_2 FILLER_66_1084 ();
 sg13g2_fill_1 FILLER_66_1100 ();
 sg13g2_fill_1 FILLER_66_1155 ();
 sg13g2_fill_1 FILLER_66_1288 ();
 sg13g2_decap_4 FILLER_66_1313 ();
 sg13g2_fill_1 FILLER_66_1317 ();
 sg13g2_fill_2 FILLER_66_1324 ();
 sg13g2_fill_1 FILLER_66_1326 ();
 sg13g2_fill_2 FILLER_66_1337 ();
 sg13g2_fill_2 FILLER_66_1352 ();
 sg13g2_fill_2 FILLER_66_1364 ();
 sg13g2_fill_2 FILLER_66_1378 ();
 sg13g2_fill_1 FILLER_66_1385 ();
 sg13g2_fill_1 FILLER_66_1393 ();
 sg13g2_fill_1 FILLER_66_1425 ();
 sg13g2_fill_2 FILLER_66_1431 ();
 sg13g2_fill_1 FILLER_66_1446 ();
 sg13g2_fill_2 FILLER_66_1471 ();
 sg13g2_fill_2 FILLER_66_1482 ();
 sg13g2_fill_1 FILLER_66_1484 ();
 sg13g2_fill_1 FILLER_66_1508 ();
 sg13g2_fill_1 FILLER_66_1547 ();
 sg13g2_fill_2 FILLER_66_1556 ();
 sg13g2_fill_2 FILLER_66_1583 ();
 sg13g2_fill_2 FILLER_66_1599 ();
 sg13g2_fill_1 FILLER_66_1601 ();
 sg13g2_decap_4 FILLER_66_1621 ();
 sg13g2_fill_1 FILLER_66_1625 ();
 sg13g2_fill_1 FILLER_66_1642 ();
 sg13g2_fill_2 FILLER_66_1649 ();
 sg13g2_fill_2 FILLER_66_1665 ();
 sg13g2_fill_1 FILLER_66_1667 ();
 sg13g2_fill_1 FILLER_66_1733 ();
 sg13g2_fill_1 FILLER_66_1784 ();
 sg13g2_fill_1 FILLER_66_1789 ();
 sg13g2_fill_1 FILLER_66_1842 ();
 sg13g2_fill_2 FILLER_66_1874 ();
 sg13g2_fill_2 FILLER_66_1885 ();
 sg13g2_fill_1 FILLER_66_1887 ();
 sg13g2_fill_2 FILLER_66_1892 ();
 sg13g2_fill_1 FILLER_66_1894 ();
 sg13g2_decap_4 FILLER_66_1903 ();
 sg13g2_fill_2 FILLER_66_1907 ();
 sg13g2_fill_1 FILLER_66_1919 ();
 sg13g2_fill_2 FILLER_66_1960 ();
 sg13g2_fill_2 FILLER_66_1988 ();
 sg13g2_fill_1 FILLER_66_1990 ();
 sg13g2_fill_2 FILLER_66_1996 ();
 sg13g2_fill_1 FILLER_66_1998 ();
 sg13g2_fill_2 FILLER_66_2009 ();
 sg13g2_fill_1 FILLER_66_2025 ();
 sg13g2_fill_1 FILLER_66_2038 ();
 sg13g2_fill_1 FILLER_66_2063 ();
 sg13g2_fill_2 FILLER_66_2080 ();
 sg13g2_fill_1 FILLER_66_2166 ();
 sg13g2_fill_2 FILLER_66_2175 ();
 sg13g2_fill_1 FILLER_66_2177 ();
 sg13g2_fill_1 FILLER_66_2182 ();
 sg13g2_fill_2 FILLER_66_2226 ();
 sg13g2_fill_1 FILLER_66_2228 ();
 sg13g2_fill_2 FILLER_66_2295 ();
 sg13g2_fill_1 FILLER_66_2297 ();
 sg13g2_fill_2 FILLER_66_2334 ();
 sg13g2_fill_2 FILLER_66_2350 ();
 sg13g2_fill_1 FILLER_66_2352 ();
 sg13g2_fill_2 FILLER_66_2435 ();
 sg13g2_fill_1 FILLER_66_2437 ();
 sg13g2_fill_1 FILLER_66_2456 ();
 sg13g2_fill_2 FILLER_66_2501 ();
 sg13g2_fill_1 FILLER_66_2552 ();
 sg13g2_fill_1 FILLER_66_2562 ();
 sg13g2_decap_8 FILLER_66_2591 ();
 sg13g2_decap_8 FILLER_66_2654 ();
 sg13g2_decap_8 FILLER_66_2661 ();
 sg13g2_decap_4 FILLER_66_2668 ();
 sg13g2_fill_2 FILLER_66_2672 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_59 ();
 sg13g2_fill_2 FILLER_67_66 ();
 sg13g2_fill_2 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_117 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_fill_1 FILLER_67_394 ();
 sg13g2_fill_1 FILLER_67_414 ();
 sg13g2_fill_1 FILLER_67_441 ();
 sg13g2_fill_2 FILLER_67_460 ();
 sg13g2_fill_2 FILLER_67_636 ();
 sg13g2_fill_1 FILLER_67_638 ();
 sg13g2_fill_1 FILLER_67_657 ();
 sg13g2_fill_2 FILLER_67_667 ();
 sg13g2_fill_1 FILLER_67_669 ();
 sg13g2_fill_2 FILLER_67_687 ();
 sg13g2_fill_1 FILLER_67_689 ();
 sg13g2_fill_2 FILLER_67_699 ();
 sg13g2_fill_1 FILLER_67_701 ();
 sg13g2_fill_2 FILLER_67_738 ();
 sg13g2_fill_2 FILLER_67_753 ();
 sg13g2_fill_1 FILLER_67_755 ();
 sg13g2_fill_1 FILLER_67_782 ();
 sg13g2_fill_1 FILLER_67_802 ();
 sg13g2_fill_1 FILLER_67_853 ();
 sg13g2_fill_2 FILLER_67_917 ();
 sg13g2_fill_1 FILLER_67_919 ();
 sg13g2_fill_1 FILLER_67_992 ();
 sg13g2_fill_2 FILLER_67_1005 ();
 sg13g2_fill_1 FILLER_67_1007 ();
 sg13g2_fill_1 FILLER_67_1115 ();
 sg13g2_fill_2 FILLER_67_1125 ();
 sg13g2_fill_1 FILLER_67_1149 ();
 sg13g2_fill_2 FILLER_67_1155 ();
 sg13g2_fill_1 FILLER_67_1157 ();
 sg13g2_fill_2 FILLER_67_1177 ();
 sg13g2_fill_2 FILLER_67_1210 ();
 sg13g2_fill_1 FILLER_67_1212 ();
 sg13g2_fill_1 FILLER_67_1222 ();
 sg13g2_fill_2 FILLER_67_1241 ();
 sg13g2_fill_2 FILLER_67_1253 ();
 sg13g2_fill_1 FILLER_67_1255 ();
 sg13g2_decap_8 FILLER_67_1269 ();
 sg13g2_fill_1 FILLER_67_1276 ();
 sg13g2_fill_1 FILLER_67_1296 ();
 sg13g2_fill_1 FILLER_67_1341 ();
 sg13g2_fill_1 FILLER_67_1350 ();
 sg13g2_fill_1 FILLER_67_1376 ();
 sg13g2_fill_1 FILLER_67_1403 ();
 sg13g2_fill_2 FILLER_67_1417 ();
 sg13g2_fill_1 FILLER_67_1419 ();
 sg13g2_fill_1 FILLER_67_1438 ();
 sg13g2_fill_2 FILLER_67_1460 ();
 sg13g2_fill_2 FILLER_67_1488 ();
 sg13g2_fill_1 FILLER_67_1490 ();
 sg13g2_fill_2 FILLER_67_1538 ();
 sg13g2_fill_2 FILLER_67_1553 ();
 sg13g2_fill_1 FILLER_67_1560 ();
 sg13g2_decap_8 FILLER_67_1619 ();
 sg13g2_decap_4 FILLER_67_1626 ();
 sg13g2_fill_2 FILLER_67_1642 ();
 sg13g2_fill_1 FILLER_67_1644 ();
 sg13g2_fill_1 FILLER_67_1654 ();
 sg13g2_decap_8 FILLER_67_1664 ();
 sg13g2_fill_1 FILLER_67_1671 ();
 sg13g2_fill_1 FILLER_67_1685 ();
 sg13g2_fill_2 FILLER_67_1699 ();
 sg13g2_fill_1 FILLER_67_1701 ();
 sg13g2_fill_2 FILLER_67_1744 ();
 sg13g2_fill_2 FILLER_67_1772 ();
 sg13g2_fill_1 FILLER_67_1804 ();
 sg13g2_fill_2 FILLER_67_1819 ();
 sg13g2_fill_2 FILLER_67_1856 ();
 sg13g2_fill_1 FILLER_67_1858 ();
 sg13g2_fill_2 FILLER_67_1882 ();
 sg13g2_decap_8 FILLER_67_1912 ();
 sg13g2_fill_2 FILLER_67_1928 ();
 sg13g2_fill_1 FILLER_67_1930 ();
 sg13g2_decap_8 FILLER_67_1948 ();
 sg13g2_decap_4 FILLER_67_1955 ();
 sg13g2_fill_2 FILLER_67_1975 ();
 sg13g2_fill_2 FILLER_67_1991 ();
 sg13g2_fill_2 FILLER_67_2008 ();
 sg13g2_decap_4 FILLER_67_2027 ();
 sg13g2_decap_4 FILLER_67_2049 ();
 sg13g2_fill_1 FILLER_67_2058 ();
 sg13g2_fill_1 FILLER_67_2073 ();
 sg13g2_decap_4 FILLER_67_2101 ();
 sg13g2_fill_2 FILLER_67_2105 ();
 sg13g2_fill_2 FILLER_67_2111 ();
 sg13g2_fill_1 FILLER_67_2113 ();
 sg13g2_fill_2 FILLER_67_2199 ();
 sg13g2_fill_1 FILLER_67_2201 ();
 sg13g2_fill_2 FILLER_67_2314 ();
 sg13g2_fill_1 FILLER_67_2394 ();
 sg13g2_fill_1 FILLER_67_2441 ();
 sg13g2_fill_1 FILLER_67_2468 ();
 sg13g2_fill_2 FILLER_67_2509 ();
 sg13g2_fill_1 FILLER_67_2535 ();
 sg13g2_fill_1 FILLER_67_2568 ();
 sg13g2_fill_1 FILLER_67_2634 ();
 sg13g2_decap_8 FILLER_67_2665 ();
 sg13g2_fill_2 FILLER_67_2672 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_51 ();
 sg13g2_fill_2 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_89 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_1 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_fill_1 FILLER_68_279 ();
 sg13g2_fill_2 FILLER_68_301 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_fill_2 FILLER_68_469 ();
 sg13g2_fill_1 FILLER_68_522 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_600 ();
 sg13g2_fill_2 FILLER_68_620 ();
 sg13g2_fill_2 FILLER_68_726 ();
 sg13g2_fill_2 FILLER_68_821 ();
 sg13g2_fill_1 FILLER_68_863 ();
 sg13g2_fill_2 FILLER_68_873 ();
 sg13g2_fill_2 FILLER_68_892 ();
 sg13g2_fill_2 FILLER_68_900 ();
 sg13g2_fill_2 FILLER_68_907 ();
 sg13g2_fill_1 FILLER_68_920 ();
 sg13g2_fill_1 FILLER_68_927 ();
 sg13g2_fill_1 FILLER_68_950 ();
 sg13g2_fill_2 FILLER_68_961 ();
 sg13g2_fill_1 FILLER_68_963 ();
 sg13g2_fill_1 FILLER_68_999 ();
 sg13g2_fill_1 FILLER_68_1051 ();
 sg13g2_fill_1 FILLER_68_1071 ();
 sg13g2_fill_2 FILLER_68_1097 ();
 sg13g2_fill_1 FILLER_68_1170 ();
 sg13g2_fill_1 FILLER_68_1191 ();
 sg13g2_fill_1 FILLER_68_1240 ();
 sg13g2_fill_1 FILLER_68_1250 ();
 sg13g2_decap_8 FILLER_68_1312 ();
 sg13g2_fill_2 FILLER_68_1319 ();
 sg13g2_fill_1 FILLER_68_1321 ();
 sg13g2_decap_4 FILLER_68_1335 ();
 sg13g2_fill_1 FILLER_68_1339 ();
 sg13g2_decap_8 FILLER_68_1351 ();
 sg13g2_decap_4 FILLER_68_1367 ();
 sg13g2_fill_2 FILLER_68_1371 ();
 sg13g2_fill_1 FILLER_68_1383 ();
 sg13g2_fill_2 FILLER_68_1394 ();
 sg13g2_fill_1 FILLER_68_1438 ();
 sg13g2_fill_2 FILLER_68_1460 ();
 sg13g2_fill_2 FILLER_68_1517 ();
 sg13g2_fill_2 FILLER_68_1542 ();
 sg13g2_fill_1 FILLER_68_1553 ();
 sg13g2_fill_2 FILLER_68_1571 ();
 sg13g2_fill_1 FILLER_68_1579 ();
 sg13g2_fill_2 FILLER_68_1598 ();
 sg13g2_fill_2 FILLER_68_1650 ();
 sg13g2_fill_1 FILLER_68_1652 ();
 sg13g2_fill_1 FILLER_68_1669 ();
 sg13g2_decap_8 FILLER_68_1680 ();
 sg13g2_decap_8 FILLER_68_1687 ();
 sg13g2_fill_2 FILLER_68_1694 ();
 sg13g2_fill_1 FILLER_68_1714 ();
 sg13g2_fill_2 FILLER_68_1755 ();
 sg13g2_decap_4 FILLER_68_1780 ();
 sg13g2_fill_2 FILLER_68_1784 ();
 sg13g2_fill_1 FILLER_68_1794 ();
 sg13g2_fill_2 FILLER_68_1898 ();
 sg13g2_fill_1 FILLER_68_1900 ();
 sg13g2_fill_1 FILLER_68_1934 ();
 sg13g2_fill_2 FILLER_68_1948 ();
 sg13g2_fill_2 FILLER_68_1988 ();
 sg13g2_fill_1 FILLER_68_2002 ();
 sg13g2_decap_8 FILLER_68_2093 ();
 sg13g2_decap_4 FILLER_68_2100 ();
 sg13g2_fill_1 FILLER_68_2104 ();
 sg13g2_fill_2 FILLER_68_2186 ();
 sg13g2_fill_1 FILLER_68_2188 ();
 sg13g2_fill_2 FILLER_68_2208 ();
 sg13g2_fill_1 FILLER_68_2279 ();
 sg13g2_fill_1 FILLER_68_2316 ();
 sg13g2_fill_2 FILLER_68_2359 ();
 sg13g2_fill_1 FILLER_68_2371 ();
 sg13g2_fill_1 FILLER_68_2425 ();
 sg13g2_fill_2 FILLER_68_2439 ();
 sg13g2_fill_1 FILLER_68_2441 ();
 sg13g2_fill_2 FILLER_68_2447 ();
 sg13g2_fill_1 FILLER_68_2449 ();
 sg13g2_fill_2 FILLER_68_2472 ();
 sg13g2_fill_1 FILLER_68_2474 ();
 sg13g2_fill_1 FILLER_68_2502 ();
 sg13g2_fill_1 FILLER_68_2548 ();
 sg13g2_fill_1 FILLER_68_2568 ();
 sg13g2_decap_8 FILLER_68_2658 ();
 sg13g2_decap_8 FILLER_68_2665 ();
 sg13g2_fill_2 FILLER_68_2672 ();
 sg13g2_fill_1 FILLER_69_26 ();
 sg13g2_fill_2 FILLER_69_45 ();
 sg13g2_fill_2 FILLER_69_102 ();
 sg13g2_fill_2 FILLER_69_175 ();
 sg13g2_fill_2 FILLER_69_229 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_1 FILLER_69_370 ();
 sg13g2_fill_2 FILLER_69_585 ();
 sg13g2_fill_2 FILLER_69_636 ();
 sg13g2_fill_1 FILLER_69_647 ();
 sg13g2_fill_1 FILLER_69_673 ();
 sg13g2_fill_2 FILLER_69_679 ();
 sg13g2_fill_1 FILLER_69_681 ();
 sg13g2_fill_2 FILLER_69_695 ();
 sg13g2_fill_1 FILLER_69_697 ();
 sg13g2_fill_2 FILLER_69_724 ();
 sg13g2_fill_2 FILLER_69_754 ();
 sg13g2_fill_1 FILLER_69_788 ();
 sg13g2_fill_1 FILLER_69_803 ();
 sg13g2_fill_2 FILLER_69_826 ();
 sg13g2_fill_1 FILLER_69_856 ();
 sg13g2_fill_1 FILLER_69_927 ();
 sg13g2_fill_1 FILLER_69_940 ();
 sg13g2_fill_1 FILLER_69_979 ();
 sg13g2_fill_1 FILLER_69_989 ();
 sg13g2_fill_2 FILLER_69_1000 ();
 sg13g2_fill_2 FILLER_69_1011 ();
 sg13g2_fill_1 FILLER_69_1013 ();
 sg13g2_fill_2 FILLER_69_1106 ();
 sg13g2_fill_1 FILLER_69_1108 ();
 sg13g2_fill_2 FILLER_69_1142 ();
 sg13g2_fill_1 FILLER_69_1144 ();
 sg13g2_fill_1 FILLER_69_1154 ();
 sg13g2_fill_2 FILLER_69_1185 ();
 sg13g2_fill_2 FILLER_69_1200 ();
 sg13g2_fill_1 FILLER_69_1202 ();
 sg13g2_decap_4 FILLER_69_1256 ();
 sg13g2_fill_2 FILLER_69_1260 ();
 sg13g2_fill_1 FILLER_69_1288 ();
 sg13g2_decap_4 FILLER_69_1294 ();
 sg13g2_decap_4 FILLER_69_1306 ();
 sg13g2_decap_4 FILLER_69_1318 ();
 sg13g2_fill_1 FILLER_69_1322 ();
 sg13g2_fill_2 FILLER_69_1332 ();
 sg13g2_fill_1 FILLER_69_1334 ();
 sg13g2_fill_1 FILLER_69_1355 ();
 sg13g2_decap_4 FILLER_69_1388 ();
 sg13g2_fill_2 FILLER_69_1405 ();
 sg13g2_fill_1 FILLER_69_1423 ();
 sg13g2_fill_1 FILLER_69_1446 ();
 sg13g2_fill_1 FILLER_69_1452 ();
 sg13g2_fill_2 FILLER_69_1481 ();
 sg13g2_fill_1 FILLER_69_1520 ();
 sg13g2_fill_2 FILLER_69_1600 ();
 sg13g2_decap_8 FILLER_69_1629 ();
 sg13g2_fill_1 FILLER_69_1644 ();
 sg13g2_decap_4 FILLER_69_1661 ();
 sg13g2_fill_2 FILLER_69_1665 ();
 sg13g2_fill_1 FILLER_69_1684 ();
 sg13g2_fill_2 FILLER_69_1728 ();
 sg13g2_fill_2 FILLER_69_1764 ();
 sg13g2_fill_2 FILLER_69_1770 ();
 sg13g2_fill_1 FILLER_69_1796 ();
 sg13g2_fill_2 FILLER_69_1881 ();
 sg13g2_fill_1 FILLER_69_1883 ();
 sg13g2_fill_2 FILLER_69_1903 ();
 sg13g2_fill_2 FILLER_69_1909 ();
 sg13g2_decap_4 FILLER_69_1919 ();
 sg13g2_decap_8 FILLER_69_1927 ();
 sg13g2_decap_4 FILLER_69_1934 ();
 sg13g2_fill_1 FILLER_69_1938 ();
 sg13g2_decap_8 FILLER_69_1948 ();
 sg13g2_decap_4 FILLER_69_1955 ();
 sg13g2_fill_1 FILLER_69_1959 ();
 sg13g2_fill_1 FILLER_69_1964 ();
 sg13g2_fill_1 FILLER_69_1969 ();
 sg13g2_decap_4 FILLER_69_1975 ();
 sg13g2_fill_1 FILLER_69_1979 ();
 sg13g2_fill_2 FILLER_69_1993 ();
 sg13g2_fill_1 FILLER_69_2017 ();
 sg13g2_decap_4 FILLER_69_2024 ();
 sg13g2_fill_1 FILLER_69_2028 ();
 sg13g2_decap_4 FILLER_69_2037 ();
 sg13g2_fill_1 FILLER_69_2041 ();
 sg13g2_decap_4 FILLER_69_2051 ();
 sg13g2_fill_1 FILLER_69_2055 ();
 sg13g2_fill_2 FILLER_69_2069 ();
 sg13g2_fill_1 FILLER_69_2071 ();
 sg13g2_decap_4 FILLER_69_2124 ();
 sg13g2_fill_1 FILLER_69_2154 ();
 sg13g2_fill_2 FILLER_69_2165 ();
 sg13g2_fill_1 FILLER_69_2167 ();
 sg13g2_fill_1 FILLER_69_2198 ();
 sg13g2_fill_1 FILLER_69_2323 ();
 sg13g2_fill_1 FILLER_69_2334 ();
 sg13g2_fill_2 FILLER_69_2481 ();
 sg13g2_fill_1 FILLER_69_2483 ();
 sg13g2_fill_2 FILLER_69_2510 ();
 sg13g2_fill_1 FILLER_69_2522 ();
 sg13g2_fill_1 FILLER_69_2532 ();
 sg13g2_fill_1 FILLER_69_2584 ();
 sg13g2_fill_1 FILLER_69_2635 ();
 sg13g2_decap_8 FILLER_69_2662 ();
 sg13g2_decap_4 FILLER_69_2669 ();
 sg13g2_fill_1 FILLER_69_2673 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_43 ();
 sg13g2_fill_1 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_94 ();
 sg13g2_fill_2 FILLER_70_121 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_fill_2 FILLER_70_207 ();
 sg13g2_fill_2 FILLER_70_432 ();
 sg13g2_fill_1 FILLER_70_488 ();
 sg13g2_fill_2 FILLER_70_532 ();
 sg13g2_fill_1 FILLER_70_622 ();
 sg13g2_fill_2 FILLER_70_637 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_fill_1 FILLER_70_702 ();
 sg13g2_fill_2 FILLER_70_760 ();
 sg13g2_fill_2 FILLER_70_775 ();
 sg13g2_fill_1 FILLER_70_817 ();
 sg13g2_fill_2 FILLER_70_874 ();
 sg13g2_fill_2 FILLER_70_902 ();
 sg13g2_fill_1 FILLER_70_913 ();
 sg13g2_fill_1 FILLER_70_948 ();
 sg13g2_fill_2 FILLER_70_962 ();
 sg13g2_fill_2 FILLER_70_1061 ();
 sg13g2_fill_1 FILLER_70_1102 ();
 sg13g2_decap_4 FILLER_70_1204 ();
 sg13g2_fill_2 FILLER_70_1213 ();
 sg13g2_decap_8 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1243 ();
 sg13g2_fill_2 FILLER_70_1276 ();
 sg13g2_fill_1 FILLER_70_1278 ();
 sg13g2_fill_2 FILLER_70_1287 ();
 sg13g2_fill_1 FILLER_70_1304 ();
 sg13g2_fill_2 FILLER_70_1342 ();
 sg13g2_fill_2 FILLER_70_1349 ();
 sg13g2_fill_1 FILLER_70_1355 ();
 sg13g2_fill_2 FILLER_70_1365 ();
 sg13g2_decap_4 FILLER_70_1371 ();
 sg13g2_fill_1 FILLER_70_1379 ();
 sg13g2_fill_1 FILLER_70_1397 ();
 sg13g2_fill_2 FILLER_70_1490 ();
 sg13g2_fill_1 FILLER_70_1532 ();
 sg13g2_fill_1 FILLER_70_1597 ();
 sg13g2_fill_2 FILLER_70_1618 ();
 sg13g2_fill_2 FILLER_70_1625 ();
 sg13g2_decap_8 FILLER_70_1640 ();
 sg13g2_fill_2 FILLER_70_1647 ();
 sg13g2_fill_2 FILLER_70_1706 ();
 sg13g2_fill_1 FILLER_70_1721 ();
 sg13g2_fill_1 FILLER_70_1761 ();
 sg13g2_fill_2 FILLER_70_1773 ();
 sg13g2_decap_8 FILLER_70_1780 ();
 sg13g2_fill_1 FILLER_70_1787 ();
 sg13g2_fill_2 FILLER_70_1796 ();
 sg13g2_decap_8 FILLER_70_1845 ();
 sg13g2_decap_4 FILLER_70_1852 ();
 sg13g2_fill_2 FILLER_70_1864 ();
 sg13g2_fill_1 FILLER_70_1866 ();
 sg13g2_fill_2 FILLER_70_1913 ();
 sg13g2_fill_2 FILLER_70_1949 ();
 sg13g2_fill_1 FILLER_70_1951 ();
 sg13g2_decap_8 FILLER_70_1983 ();
 sg13g2_decap_4 FILLER_70_1990 ();
 sg13g2_fill_1 FILLER_70_1994 ();
 sg13g2_decap_8 FILLER_70_2013 ();
 sg13g2_decap_8 FILLER_70_2020 ();
 sg13g2_decap_8 FILLER_70_2027 ();
 sg13g2_fill_1 FILLER_70_2034 ();
 sg13g2_decap_8 FILLER_70_2043 ();
 sg13g2_fill_2 FILLER_70_2050 ();
 sg13g2_fill_1 FILLER_70_2062 ();
 sg13g2_decap_8 FILLER_70_2066 ();
 sg13g2_fill_2 FILLER_70_2073 ();
 sg13g2_fill_2 FILLER_70_2080 ();
 sg13g2_fill_1 FILLER_70_2082 ();
 sg13g2_fill_2 FILLER_70_2100 ();
 sg13g2_fill_2 FILLER_70_2106 ();
 sg13g2_fill_2 FILLER_70_2121 ();
 sg13g2_fill_2 FILLER_70_2131 ();
 sg13g2_decap_8 FILLER_70_2201 ();
 sg13g2_fill_2 FILLER_70_2247 ();
 sg13g2_fill_1 FILLER_70_2249 ();
 sg13g2_fill_2 FILLER_70_2376 ();
 sg13g2_fill_1 FILLER_70_2378 ();
 sg13g2_fill_2 FILLER_70_2443 ();
 sg13g2_fill_1 FILLER_70_2445 ();
 sg13g2_fill_2 FILLER_70_2485 ();
 sg13g2_fill_2 FILLER_70_2513 ();
 sg13g2_fill_1 FILLER_70_2515 ();
 sg13g2_fill_2 FILLER_70_2568 ();
 sg13g2_fill_2 FILLER_70_2600 ();
 sg13g2_fill_1 FILLER_70_2635 ();
 sg13g2_decap_8 FILLER_70_2662 ();
 sg13g2_decap_4 FILLER_70_2669 ();
 sg13g2_fill_1 FILLER_70_2673 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_37 ();
 sg13g2_fill_2 FILLER_71_98 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_71_495 ();
 sg13g2_fill_1 FILLER_71_548 ();
 sg13g2_fill_1 FILLER_71_603 ();
 sg13g2_fill_1 FILLER_71_665 ();
 sg13g2_fill_2 FILLER_71_713 ();
 sg13g2_fill_1 FILLER_71_780 ();
 sg13g2_fill_2 FILLER_71_795 ();
 sg13g2_fill_1 FILLER_71_814 ();
 sg13g2_fill_2 FILLER_71_823 ();
 sg13g2_fill_1 FILLER_71_851 ();
 sg13g2_fill_2 FILLER_71_862 ();
 sg13g2_fill_1 FILLER_71_864 ();
 sg13g2_fill_2 FILLER_71_882 ();
 sg13g2_fill_1 FILLER_71_884 ();
 sg13g2_fill_2 FILLER_71_902 ();
 sg13g2_fill_1 FILLER_71_904 ();
 sg13g2_fill_2 FILLER_71_931 ();
 sg13g2_fill_1 FILLER_71_933 ();
 sg13g2_fill_1 FILLER_71_974 ();
 sg13g2_fill_2 FILLER_71_993 ();
 sg13g2_fill_1 FILLER_71_995 ();
 sg13g2_fill_1 FILLER_71_1001 ();
 sg13g2_fill_2 FILLER_71_1012 ();
 sg13g2_fill_1 FILLER_71_1014 ();
 sg13g2_fill_2 FILLER_71_1046 ();
 sg13g2_fill_2 FILLER_71_1152 ();
 sg13g2_fill_1 FILLER_71_1180 ();
 sg13g2_fill_2 FILLER_71_1206 ();
 sg13g2_decap_4 FILLER_71_1212 ();
 sg13g2_fill_1 FILLER_71_1225 ();
 sg13g2_fill_2 FILLER_71_1238 ();
 sg13g2_fill_1 FILLER_71_1240 ();
 sg13g2_fill_2 FILLER_71_1249 ();
 sg13g2_fill_1 FILLER_71_1281 ();
 sg13g2_fill_1 FILLER_71_1302 ();
 sg13g2_fill_2 FILLER_71_1316 ();
 sg13g2_fill_2 FILLER_71_1323 ();
 sg13g2_fill_2 FILLER_71_1330 ();
 sg13g2_fill_2 FILLER_71_1348 ();
 sg13g2_decap_8 FILLER_71_1392 ();
 sg13g2_decap_8 FILLER_71_1399 ();
 sg13g2_fill_2 FILLER_71_1406 ();
 sg13g2_fill_1 FILLER_71_1408 ();
 sg13g2_fill_2 FILLER_71_1436 ();
 sg13g2_fill_1 FILLER_71_1438 ();
 sg13g2_fill_1 FILLER_71_1472 ();
 sg13g2_fill_2 FILLER_71_1486 ();
 sg13g2_fill_1 FILLER_71_1513 ();
 sg13g2_fill_2 FILLER_71_1527 ();
 sg13g2_fill_1 FILLER_71_1542 ();
 sg13g2_fill_2 FILLER_71_1551 ();
 sg13g2_fill_1 FILLER_71_1609 ();
 sg13g2_decap_8 FILLER_71_1660 ();
 sg13g2_fill_2 FILLER_71_1667 ();
 sg13g2_fill_2 FILLER_71_1682 ();
 sg13g2_fill_1 FILLER_71_1684 ();
 sg13g2_fill_1 FILLER_71_1743 ();
 sg13g2_fill_1 FILLER_71_1762 ();
 sg13g2_fill_2 FILLER_71_1768 ();
 sg13g2_fill_1 FILLER_71_1770 ();
 sg13g2_decap_4 FILLER_71_1776 ();
 sg13g2_fill_1 FILLER_71_1832 ();
 sg13g2_decap_8 FILLER_71_1841 ();
 sg13g2_fill_2 FILLER_71_1859 ();
 sg13g2_fill_1 FILLER_71_1861 ();
 sg13g2_decap_4 FILLER_71_1898 ();
 sg13g2_decap_8 FILLER_71_1917 ();
 sg13g2_fill_2 FILLER_71_1924 ();
 sg13g2_fill_2 FILLER_71_1930 ();
 sg13g2_decap_4 FILLER_71_1967 ();
 sg13g2_fill_2 FILLER_71_1989 ();
 sg13g2_decap_4 FILLER_71_2026 ();
 sg13g2_fill_2 FILLER_71_2030 ();
 sg13g2_decap_4 FILLER_71_2044 ();
 sg13g2_fill_1 FILLER_71_2048 ();
 sg13g2_fill_1 FILLER_71_2078 ();
 sg13g2_fill_1 FILLER_71_2095 ();
 sg13g2_decap_8 FILLER_71_2165 ();
 sg13g2_fill_1 FILLER_71_2172 ();
 sg13g2_fill_2 FILLER_71_2225 ();
 sg13g2_fill_1 FILLER_71_2258 ();
 sg13g2_fill_2 FILLER_71_2268 ();
 sg13g2_fill_1 FILLER_71_2279 ();
 sg13g2_fill_1 FILLER_71_2309 ();
 sg13g2_fill_2 FILLER_71_2328 ();
 sg13g2_fill_2 FILLER_71_2383 ();
 sg13g2_fill_1 FILLER_71_2385 ();
 sg13g2_fill_2 FILLER_71_2405 ();
 sg13g2_fill_1 FILLER_71_2407 ();
 sg13g2_fill_2 FILLER_71_2474 ();
 sg13g2_fill_1 FILLER_71_2476 ();
 sg13g2_fill_1 FILLER_71_2496 ();
 sg13g2_fill_2 FILLER_71_2524 ();
 sg13g2_fill_2 FILLER_71_2564 ();
 sg13g2_fill_1 FILLER_71_2576 ();
 sg13g2_fill_2 FILLER_71_2617 ();
 sg13g2_fill_1 FILLER_71_2619 ();
 sg13g2_fill_2 FILLER_71_2630 ();
 sg13g2_decap_8 FILLER_71_2658 ();
 sg13g2_decap_8 FILLER_71_2665 ();
 sg13g2_fill_2 FILLER_71_2672 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_130 ();
 sg13g2_fill_1 FILLER_72_184 ();
 sg13g2_fill_2 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_363 ();
 sg13g2_fill_1 FILLER_72_411 ();
 sg13g2_fill_2 FILLER_72_494 ();
 sg13g2_fill_2 FILLER_72_535 ();
 sg13g2_fill_2 FILLER_72_546 ();
 sg13g2_fill_1 FILLER_72_564 ();
 sg13g2_fill_1 FILLER_72_570 ();
 sg13g2_fill_1 FILLER_72_619 ();
 sg13g2_fill_1 FILLER_72_647 ();
 sg13g2_fill_1 FILLER_72_657 ();
 sg13g2_fill_2 FILLER_72_696 ();
 sg13g2_fill_2 FILLER_72_721 ();
 sg13g2_fill_1 FILLER_72_756 ();
 sg13g2_fill_1 FILLER_72_837 ();
 sg13g2_fill_2 FILLER_72_864 ();
 sg13g2_fill_1 FILLER_72_871 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_fill_2 FILLER_72_921 ();
 sg13g2_fill_1 FILLER_72_943 ();
 sg13g2_fill_2 FILLER_72_957 ();
 sg13g2_fill_2 FILLER_72_969 ();
 sg13g2_fill_1 FILLER_72_1003 ();
 sg13g2_fill_1 FILLER_72_1060 ();
 sg13g2_fill_1 FILLER_72_1123 ();
 sg13g2_fill_1 FILLER_72_1134 ();
 sg13g2_fill_1 FILLER_72_1165 ();
 sg13g2_fill_2 FILLER_72_1195 ();
 sg13g2_fill_1 FILLER_72_1278 ();
 sg13g2_decap_8 FILLER_72_1292 ();
 sg13g2_fill_2 FILLER_72_1299 ();
 sg13g2_fill_1 FILLER_72_1301 ();
 sg13g2_fill_1 FILLER_72_1330 ();
 sg13g2_decap_8 FILLER_72_1349 ();
 sg13g2_fill_2 FILLER_72_1356 ();
 sg13g2_fill_1 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1373 ();
 sg13g2_fill_2 FILLER_72_1380 ();
 sg13g2_fill_1 FILLER_72_1382 ();
 sg13g2_fill_1 FILLER_72_1391 ();
 sg13g2_decap_8 FILLER_72_1400 ();
 sg13g2_fill_1 FILLER_72_1407 ();
 sg13g2_fill_1 FILLER_72_1421 ();
 sg13g2_fill_1 FILLER_72_1456 ();
 sg13g2_fill_1 FILLER_72_1501 ();
 sg13g2_fill_1 FILLER_72_1528 ();
 sg13g2_fill_1 FILLER_72_1558 ();
 sg13g2_fill_2 FILLER_72_1580 ();
 sg13g2_fill_1 FILLER_72_1582 ();
 sg13g2_fill_1 FILLER_72_1626 ();
 sg13g2_fill_2 FILLER_72_1661 ();
 sg13g2_fill_2 FILLER_72_1679 ();
 sg13g2_fill_1 FILLER_72_1681 ();
 sg13g2_fill_1 FILLER_72_1700 ();
 sg13g2_fill_2 FILLER_72_1736 ();
 sg13g2_fill_1 FILLER_72_1738 ();
 sg13g2_fill_2 FILLER_72_1753 ();
 sg13g2_fill_1 FILLER_72_1763 ();
 sg13g2_fill_1 FILLER_72_1770 ();
 sg13g2_fill_2 FILLER_72_1796 ();
 sg13g2_fill_1 FILLER_72_1798 ();
 sg13g2_fill_2 FILLER_72_1805 ();
 sg13g2_fill_2 FILLER_72_1819 ();
 sg13g2_decap_4 FILLER_72_1827 ();
 sg13g2_fill_2 FILLER_72_1831 ();
 sg13g2_decap_8 FILLER_72_1861 ();
 sg13g2_fill_2 FILLER_72_1868 ();
 sg13g2_fill_1 FILLER_72_1883 ();
 sg13g2_decap_8 FILLER_72_1892 ();
 sg13g2_decap_8 FILLER_72_1904 ();
 sg13g2_fill_2 FILLER_72_1911 ();
 sg13g2_decap_4 FILLER_72_1986 ();
 sg13g2_fill_2 FILLER_72_2053 ();
 sg13g2_decap_4 FILLER_72_2060 ();
 sg13g2_fill_2 FILLER_72_2089 ();
 sg13g2_fill_1 FILLER_72_2091 ();
 sg13g2_fill_2 FILLER_72_2182 ();
 sg13g2_fill_1 FILLER_72_2202 ();
 sg13g2_fill_2 FILLER_72_2217 ();
 sg13g2_fill_1 FILLER_72_2229 ();
 sg13g2_fill_1 FILLER_72_2282 ();
 sg13g2_fill_2 FILLER_72_2293 ();
 sg13g2_fill_1 FILLER_72_2321 ();
 sg13g2_fill_2 FILLER_72_2370 ();
 sg13g2_fill_2 FILLER_72_2413 ();
 sg13g2_fill_1 FILLER_72_2415 ();
 sg13g2_fill_2 FILLER_72_2430 ();
 sg13g2_fill_2 FILLER_72_2480 ();
 sg13g2_fill_1 FILLER_72_2503 ();
 sg13g2_decap_4 FILLER_72_2622 ();
 sg13g2_fill_1 FILLER_72_2626 ();
 sg13g2_decap_8 FILLER_72_2666 ();
 sg13g2_fill_1 FILLER_72_2673 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_16 ();
 sg13g2_fill_1 FILLER_73_30 ();
 sg13g2_fill_1 FILLER_73_39 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_fill_1 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_2 FILLER_73_173 ();
 sg13g2_fill_2 FILLER_73_201 ();
 sg13g2_fill_1 FILLER_73_218 ();
 sg13g2_fill_1 FILLER_73_297 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_2 FILLER_73_469 ();
 sg13g2_fill_2 FILLER_73_524 ();
 sg13g2_fill_2 FILLER_73_610 ();
 sg13g2_fill_1 FILLER_73_617 ();
 sg13g2_fill_1 FILLER_73_649 ();
 sg13g2_fill_2 FILLER_73_657 ();
 sg13g2_fill_1 FILLER_73_659 ();
 sg13g2_fill_1 FILLER_73_762 ();
 sg13g2_fill_2 FILLER_73_816 ();
 sg13g2_fill_1 FILLER_73_823 ();
 sg13g2_fill_1 FILLER_73_846 ();
 sg13g2_fill_1 FILLER_73_962 ();
 sg13g2_fill_2 FILLER_73_1012 ();
 sg13g2_fill_2 FILLER_73_1029 ();
 sg13g2_fill_1 FILLER_73_1052 ();
 sg13g2_fill_2 FILLER_73_1091 ();
 sg13g2_fill_2 FILLER_73_1118 ();
 sg13g2_fill_1 FILLER_73_1120 ();
 sg13g2_fill_2 FILLER_73_1151 ();
 sg13g2_fill_1 FILLER_73_1153 ();
 sg13g2_fill_1 FILLER_73_1230 ();
 sg13g2_decap_8 FILLER_73_1251 ();
 sg13g2_decap_4 FILLER_73_1258 ();
 sg13g2_fill_2 FILLER_73_1270 ();
 sg13g2_decap_4 FILLER_73_1298 ();
 sg13g2_fill_1 FILLER_73_1302 ();
 sg13g2_fill_2 FILLER_73_1317 ();
 sg13g2_decap_8 FILLER_73_1331 ();
 sg13g2_fill_1 FILLER_73_1338 ();
 sg13g2_fill_1 FILLER_73_1348 ();
 sg13g2_fill_2 FILLER_73_1354 ();
 sg13g2_fill_2 FILLER_73_1392 ();
 sg13g2_fill_1 FILLER_73_1394 ();
 sg13g2_fill_1 FILLER_73_1421 ();
 sg13g2_fill_1 FILLER_73_1427 ();
 sg13g2_fill_1 FILLER_73_1446 ();
 sg13g2_fill_1 FILLER_73_1460 ();
 sg13g2_fill_2 FILLER_73_1488 ();
 sg13g2_fill_2 FILLER_73_1503 ();
 sg13g2_fill_1 FILLER_73_1505 ();
 sg13g2_fill_1 FILLER_73_1537 ();
 sg13g2_fill_2 FILLER_73_1556 ();
 sg13g2_fill_1 FILLER_73_1558 ();
 sg13g2_fill_2 FILLER_73_1564 ();
 sg13g2_fill_1 FILLER_73_1614 ();
 sg13g2_fill_2 FILLER_73_1688 ();
 sg13g2_fill_2 FILLER_73_1713 ();
 sg13g2_fill_2 FILLER_73_1733 ();
 sg13g2_fill_1 FILLER_73_1735 ();
 sg13g2_fill_2 FILLER_73_1748 ();
 sg13g2_fill_1 FILLER_73_1771 ();
 sg13g2_fill_1 FILLER_73_1777 ();
 sg13g2_decap_4 FILLER_73_1792 ();
 sg13g2_fill_1 FILLER_73_1796 ();
 sg13g2_decap_8 FILLER_73_1809 ();
 sg13g2_fill_1 FILLER_73_1816 ();
 sg13g2_decap_8 FILLER_73_1825 ();
 sg13g2_decap_4 FILLER_73_1832 ();
 sg13g2_decap_4 FILLER_73_1930 ();
 sg13g2_decap_4 FILLER_73_1942 ();
 sg13g2_fill_1 FILLER_73_1946 ();
 sg13g2_fill_2 FILLER_73_1952 ();
 sg13g2_decap_8 FILLER_73_1958 ();
 sg13g2_fill_1 FILLER_73_1965 ();
 sg13g2_decap_4 FILLER_73_1969 ();
 sg13g2_fill_1 FILLER_73_1973 ();
 sg13g2_decap_8 FILLER_73_1986 ();
 sg13g2_fill_2 FILLER_73_1993 ();
 sg13g2_fill_1 FILLER_73_1995 ();
 sg13g2_decap_8 FILLER_73_2001 ();
 sg13g2_fill_2 FILLER_73_2012 ();
 sg13g2_decap_8 FILLER_73_2022 ();
 sg13g2_decap_4 FILLER_73_2079 ();
 sg13g2_fill_2 FILLER_73_2083 ();
 sg13g2_fill_1 FILLER_73_2093 ();
 sg13g2_fill_1 FILLER_73_2098 ();
 sg13g2_fill_1 FILLER_73_2103 ();
 sg13g2_fill_2 FILLER_73_2174 ();
 sg13g2_fill_1 FILLER_73_2176 ();
 sg13g2_fill_2 FILLER_73_2207 ();
 sg13g2_fill_1 FILLER_73_2232 ();
 sg13g2_fill_2 FILLER_73_2304 ();
 sg13g2_fill_2 FILLER_73_2315 ();
 sg13g2_fill_1 FILLER_73_2317 ();
 sg13g2_fill_2 FILLER_73_2337 ();
 sg13g2_fill_1 FILLER_73_2339 ();
 sg13g2_fill_2 FILLER_73_2381 ();
 sg13g2_fill_1 FILLER_73_2393 ();
 sg13g2_fill_1 FILLER_73_2403 ();
 sg13g2_fill_2 FILLER_73_2501 ();
 sg13g2_fill_1 FILLER_73_2524 ();
 sg13g2_fill_2 FILLER_73_2613 ();
 sg13g2_fill_1 FILLER_73_2615 ();
 sg13g2_decap_8 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2659 ();
 sg13g2_decap_8 FILLER_73_2666 ();
 sg13g2_fill_1 FILLER_73_2673 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_14 ();
 sg13g2_fill_1 FILLER_74_16 ();
 sg13g2_fill_2 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_147 ();
 sg13g2_fill_1 FILLER_74_189 ();
 sg13g2_fill_2 FILLER_74_199 ();
 sg13g2_fill_2 FILLER_74_210 ();
 sg13g2_fill_1 FILLER_74_262 ();
 sg13g2_fill_2 FILLER_74_302 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_390 ();
 sg13g2_fill_2 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_426 ();
 sg13g2_fill_2 FILLER_74_535 ();
 sg13g2_fill_2 FILLER_74_551 ();
 sg13g2_fill_2 FILLER_74_584 ();
 sg13g2_fill_2 FILLER_74_595 ();
 sg13g2_fill_1 FILLER_74_597 ();
 sg13g2_fill_2 FILLER_74_607 ();
 sg13g2_fill_2 FILLER_74_628 ();
 sg13g2_fill_1 FILLER_74_630 ();
 sg13g2_fill_2 FILLER_74_663 ();
 sg13g2_fill_1 FILLER_74_665 ();
 sg13g2_fill_2 FILLER_74_742 ();
 sg13g2_fill_2 FILLER_74_749 ();
 sg13g2_fill_1 FILLER_74_756 ();
 sg13g2_fill_2 FILLER_74_783 ();
 sg13g2_fill_1 FILLER_74_828 ();
 sg13g2_fill_1 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_883 ();
 sg13g2_fill_1 FILLER_74_885 ();
 sg13g2_fill_2 FILLER_74_917 ();
 sg13g2_fill_1 FILLER_74_919 ();
 sg13g2_fill_2 FILLER_74_935 ();
 sg13g2_fill_1 FILLER_74_937 ();
 sg13g2_fill_2 FILLER_74_966 ();
 sg13g2_fill_1 FILLER_74_1011 ();
 sg13g2_fill_2 FILLER_74_1106 ();
 sg13g2_fill_1 FILLER_74_1116 ();
 sg13g2_fill_2 FILLER_74_1131 ();
 sg13g2_fill_1 FILLER_74_1133 ();
 sg13g2_fill_1 FILLER_74_1160 ();
 sg13g2_fill_2 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1236 ();
 sg13g2_fill_2 FILLER_74_1243 ();
 sg13g2_fill_1 FILLER_74_1245 ();
 sg13g2_fill_2 FILLER_74_1275 ();
 sg13g2_fill_1 FILLER_74_1277 ();
 sg13g2_fill_1 FILLER_74_1282 ();
 sg13g2_fill_2 FILLER_74_1287 ();
 sg13g2_decap_8 FILLER_74_1293 ();
 sg13g2_fill_2 FILLER_74_1300 ();
 sg13g2_fill_1 FILLER_74_1302 ();
 sg13g2_fill_2 FILLER_74_1335 ();
 sg13g2_fill_1 FILLER_74_1337 ();
 sg13g2_decap_8 FILLER_74_1360 ();
 sg13g2_decap_8 FILLER_74_1367 ();
 sg13g2_fill_2 FILLER_74_1374 ();
 sg13g2_fill_1 FILLER_74_1397 ();
 sg13g2_fill_1 FILLER_74_1415 ();
 sg13g2_fill_2 FILLER_74_1433 ();
 sg13g2_fill_2 FILLER_74_1490 ();
 sg13g2_fill_2 FILLER_74_1505 ();
 sg13g2_fill_1 FILLER_74_1585 ();
 sg13g2_fill_2 FILLER_74_1600 ();
 sg13g2_fill_1 FILLER_74_1665 ();
 sg13g2_fill_2 FILLER_74_1705 ();
 sg13g2_fill_1 FILLER_74_1707 ();
 sg13g2_fill_2 FILLER_74_1791 ();
 sg13g2_fill_1 FILLER_74_1793 ();
 sg13g2_fill_1 FILLER_74_1814 ();
 sg13g2_fill_2 FILLER_74_1856 ();
 sg13g2_decap_4 FILLER_74_1881 ();
 sg13g2_fill_2 FILLER_74_1885 ();
 sg13g2_fill_2 FILLER_74_1891 ();
 sg13g2_fill_1 FILLER_74_1910 ();
 sg13g2_fill_1 FILLER_74_1929 ();
 sg13g2_fill_1 FILLER_74_1966 ();
 sg13g2_fill_1 FILLER_74_1981 ();
 sg13g2_fill_2 FILLER_74_2008 ();
 sg13g2_fill_1 FILLER_74_2010 ();
 sg13g2_fill_1 FILLER_74_2016 ();
 sg13g2_fill_2 FILLER_74_2031 ();
 sg13g2_fill_1 FILLER_74_2033 ();
 sg13g2_fill_1 FILLER_74_2038 ();
 sg13g2_decap_8 FILLER_74_2044 ();
 sg13g2_fill_2 FILLER_74_2051 ();
 sg13g2_fill_1 FILLER_74_2053 ();
 sg13g2_fill_2 FILLER_74_2066 ();
 sg13g2_decap_8 FILLER_74_2072 ();
 sg13g2_decap_4 FILLER_74_2079 ();
 sg13g2_fill_1 FILLER_74_2109 ();
 sg13g2_fill_1 FILLER_74_2130 ();
 sg13g2_fill_2 FILLER_74_2210 ();
 sg13g2_fill_1 FILLER_74_2212 ();
 sg13g2_fill_2 FILLER_74_2239 ();
 sg13g2_fill_2 FILLER_74_2267 ();
 sg13g2_fill_2 FILLER_74_2373 ();
 sg13g2_fill_2 FILLER_74_2422 ();
 sg13g2_fill_1 FILLER_74_2459 ();
 sg13g2_fill_2 FILLER_74_2567 ();
 sg13g2_fill_1 FILLER_74_2579 ();
 sg13g2_fill_1 FILLER_74_2599 ();
 sg13g2_decap_8 FILLER_74_2649 ();
 sg13g2_decap_8 FILLER_74_2656 ();
 sg13g2_decap_8 FILLER_74_2663 ();
 sg13g2_decap_4 FILLER_74_2670 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_18 ();
 sg13g2_fill_2 FILLER_75_118 ();
 sg13g2_fill_1 FILLER_75_151 ();
 sg13g2_fill_2 FILLER_75_160 ();
 sg13g2_fill_1 FILLER_75_220 ();
 sg13g2_fill_2 FILLER_75_226 ();
 sg13g2_fill_1 FILLER_75_237 ();
 sg13g2_fill_2 FILLER_75_253 ();
 sg13g2_fill_1 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_309 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_454 ();
 sg13g2_fill_2 FILLER_75_476 ();
 sg13g2_fill_2 FILLER_75_555 ();
 sg13g2_fill_2 FILLER_75_575 ();
 sg13g2_fill_1 FILLER_75_603 ();
 sg13g2_fill_1 FILLER_75_610 ();
 sg13g2_fill_2 FILLER_75_620 ();
 sg13g2_fill_1 FILLER_75_622 ();
 sg13g2_fill_2 FILLER_75_629 ();
 sg13g2_fill_1 FILLER_75_631 ();
 sg13g2_fill_1 FILLER_75_728 ();
 sg13g2_fill_2 FILLER_75_759 ();
 sg13g2_fill_2 FILLER_75_797 ();
 sg13g2_fill_2 FILLER_75_808 ();
 sg13g2_fill_2 FILLER_75_862 ();
 sg13g2_fill_1 FILLER_75_864 ();
 sg13g2_fill_2 FILLER_75_874 ();
 sg13g2_fill_2 FILLER_75_881 ();
 sg13g2_fill_1 FILLER_75_901 ();
 sg13g2_fill_2 FILLER_75_928 ();
 sg13g2_fill_1 FILLER_75_930 ();
 sg13g2_fill_2 FILLER_75_990 ();
 sg13g2_fill_1 FILLER_75_1006 ();
 sg13g2_fill_2 FILLER_75_1020 ();
 sg13g2_fill_1 FILLER_75_1039 ();
 sg13g2_fill_2 FILLER_75_1045 ();
 sg13g2_fill_1 FILLER_75_1064 ();
 sg13g2_fill_1 FILLER_75_1075 ();
 sg13g2_fill_1 FILLER_75_1097 ();
 sg13g2_fill_1 FILLER_75_1106 ();
 sg13g2_fill_2 FILLER_75_1131 ();
 sg13g2_fill_2 FILLER_75_1147 ();
 sg13g2_fill_1 FILLER_75_1149 ();
 sg13g2_fill_2 FILLER_75_1176 ();
 sg13g2_fill_1 FILLER_75_1178 ();
 sg13g2_fill_2 FILLER_75_1188 ();
 sg13g2_fill_2 FILLER_75_1204 ();
 sg13g2_fill_1 FILLER_75_1245 ();
 sg13g2_fill_1 FILLER_75_1309 ();
 sg13g2_fill_2 FILLER_75_1318 ();
 sg13g2_fill_1 FILLER_75_1320 ();
 sg13g2_fill_2 FILLER_75_1347 ();
 sg13g2_decap_8 FILLER_75_1354 ();
 sg13g2_decap_4 FILLER_75_1361 ();
 sg13g2_fill_1 FILLER_75_1386 ();
 sg13g2_decap_4 FILLER_75_1392 ();
 sg13g2_fill_2 FILLER_75_1396 ();
 sg13g2_fill_2 FILLER_75_1424 ();
 sg13g2_fill_2 FILLER_75_1435 ();
 sg13g2_fill_2 FILLER_75_1459 ();
 sg13g2_fill_1 FILLER_75_1461 ();
 sg13g2_fill_1 FILLER_75_1477 ();
 sg13g2_fill_2 FILLER_75_1530 ();
 sg13g2_fill_2 FILLER_75_1592 ();
 sg13g2_fill_2 FILLER_75_1707 ();
 sg13g2_fill_1 FILLER_75_1719 ();
 sg13g2_decap_4 FILLER_75_1732 ();
 sg13g2_fill_2 FILLER_75_1736 ();
 sg13g2_decap_4 FILLER_75_1752 ();
 sg13g2_decap_8 FILLER_75_1769 ();
 sg13g2_fill_2 FILLER_75_1776 ();
 sg13g2_fill_1 FILLER_75_1778 ();
 sg13g2_fill_2 FILLER_75_1792 ();
 sg13g2_fill_2 FILLER_75_1810 ();
 sg13g2_fill_1 FILLER_75_1812 ();
 sg13g2_decap_8 FILLER_75_1828 ();
 sg13g2_fill_1 FILLER_75_1835 ();
 sg13g2_decap_4 FILLER_75_1857 ();
 sg13g2_fill_1 FILLER_75_1861 ();
 sg13g2_fill_1 FILLER_75_1872 ();
 sg13g2_decap_4 FILLER_75_1881 ();
 sg13g2_fill_1 FILLER_75_1885 ();
 sg13g2_fill_2 FILLER_75_1921 ();
 sg13g2_fill_2 FILLER_75_1931 ();
 sg13g2_fill_2 FILLER_75_1983 ();
 sg13g2_fill_1 FILLER_75_1985 ();
 sg13g2_fill_2 FILLER_75_1990 ();
 sg13g2_fill_1 FILLER_75_1992 ();
 sg13g2_decap_4 FILLER_75_2003 ();
 sg13g2_fill_1 FILLER_75_2015 ();
 sg13g2_fill_1 FILLER_75_2022 ();
 sg13g2_fill_2 FILLER_75_2053 ();
 sg13g2_fill_2 FILLER_75_2060 ();
 sg13g2_decap_8 FILLER_75_2066 ();
 sg13g2_fill_2 FILLER_75_2073 ();
 sg13g2_fill_1 FILLER_75_2075 ();
 sg13g2_fill_2 FILLER_75_2116 ();
 sg13g2_fill_2 FILLER_75_2189 ();
 sg13g2_fill_1 FILLER_75_2225 ();
 sg13g2_fill_2 FILLER_75_2241 ();
 sg13g2_fill_2 FILLER_75_2266 ();
 sg13g2_fill_2 FILLER_75_2313 ();
 sg13g2_fill_1 FILLER_75_2315 ();
 sg13g2_fill_1 FILLER_75_2347 ();
 sg13g2_fill_2 FILLER_75_2490 ();
 sg13g2_fill_1 FILLER_75_2492 ();
 sg13g2_fill_1 FILLER_75_2502 ();
 sg13g2_fill_1 FILLER_75_2536 ();
 sg13g2_fill_2 FILLER_75_2584 ();
 sg13g2_fill_2 FILLER_75_2621 ();
 sg13g2_fill_1 FILLER_75_2623 ();
 sg13g2_decap_8 FILLER_75_2650 ();
 sg13g2_decap_8 FILLER_75_2657 ();
 sg13g2_decap_8 FILLER_75_2664 ();
 sg13g2_fill_2 FILLER_75_2671 ();
 sg13g2_fill_1 FILLER_75_2673 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_2 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_16 ();
 sg13g2_fill_2 FILLER_76_85 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_285 ();
 sg13g2_fill_1 FILLER_76_444 ();
 sg13g2_fill_1 FILLER_76_463 ();
 sg13g2_fill_1 FILLER_76_530 ();
 sg13g2_fill_2 FILLER_76_549 ();
 sg13g2_fill_1 FILLER_76_562 ();
 sg13g2_fill_2 FILLER_76_586 ();
 sg13g2_fill_1 FILLER_76_588 ();
 sg13g2_fill_2 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_601 ();
 sg13g2_fill_1 FILLER_76_665 ();
 sg13g2_fill_1 FILLER_76_729 ();
 sg13g2_fill_2 FILLER_76_780 ();
 sg13g2_fill_1 FILLER_76_788 ();
 sg13g2_fill_2 FILLER_76_882 ();
 sg13g2_fill_1 FILLER_76_884 ();
 sg13g2_fill_2 FILLER_76_896 ();
 sg13g2_fill_2 FILLER_76_912 ();
 sg13g2_fill_1 FILLER_76_943 ();
 sg13g2_fill_1 FILLER_76_991 ();
 sg13g2_fill_1 FILLER_76_1028 ();
 sg13g2_fill_2 FILLER_76_1039 ();
 sg13g2_fill_1 FILLER_76_1041 ();
 sg13g2_fill_2 FILLER_76_1051 ();
 sg13g2_fill_1 FILLER_76_1053 ();
 sg13g2_fill_1 FILLER_76_1094 ();
 sg13g2_fill_1 FILLER_76_1101 ();
 sg13g2_fill_2 FILLER_76_1132 ();
 sg13g2_fill_1 FILLER_76_1134 ();
 sg13g2_fill_2 FILLER_76_1153 ();
 sg13g2_fill_1 FILLER_76_1155 ();
 sg13g2_fill_2 FILLER_76_1216 ();
 sg13g2_fill_2 FILLER_76_1269 ();
 sg13g2_fill_2 FILLER_76_1283 ();
 sg13g2_decap_8 FILLER_76_1293 ();
 sg13g2_decap_4 FILLER_76_1300 ();
 sg13g2_fill_2 FILLER_76_1358 ();
 sg13g2_fill_1 FILLER_76_1360 ();
 sg13g2_decap_4 FILLER_76_1376 ();
 sg13g2_fill_2 FILLER_76_1388 ();
 sg13g2_decap_4 FILLER_76_1398 ();
 sg13g2_fill_2 FILLER_76_1402 ();
 sg13g2_fill_2 FILLER_76_1455 ();
 sg13g2_fill_1 FILLER_76_1457 ();
 sg13g2_fill_2 FILLER_76_1532 ();
 sg13g2_fill_2 FILLER_76_1554 ();
 sg13g2_fill_2 FILLER_76_1570 ();
 sg13g2_fill_1 FILLER_76_1701 ();
 sg13g2_decap_8 FILLER_76_1723 ();
 sg13g2_decap_8 FILLER_76_1730 ();
 sg13g2_decap_8 FILLER_76_1737 ();
 sg13g2_decap_4 FILLER_76_1744 ();
 sg13g2_fill_2 FILLER_76_1779 ();
 sg13g2_fill_1 FILLER_76_1781 ();
 sg13g2_fill_2 FILLER_76_1800 ();
 sg13g2_fill_1 FILLER_76_1802 ();
 sg13g2_fill_2 FILLER_76_1812 ();
 sg13g2_fill_1 FILLER_76_1865 ();
 sg13g2_fill_1 FILLER_76_1870 ();
 sg13g2_fill_2 FILLER_76_1885 ();
 sg13g2_fill_1 FILLER_76_1887 ();
 sg13g2_fill_2 FILLER_76_1905 ();
 sg13g2_fill_1 FILLER_76_1954 ();
 sg13g2_decap_4 FILLER_76_1961 ();
 sg13g2_fill_2 FILLER_76_1973 ();
 sg13g2_fill_2 FILLER_76_2013 ();
 sg13g2_fill_1 FILLER_76_2015 ();
 sg13g2_fill_2 FILLER_76_2020 ();
 sg13g2_fill_2 FILLER_76_2027 ();
 sg13g2_fill_2 FILLER_76_2048 ();
 sg13g2_fill_2 FILLER_76_2090 ();
 sg13g2_fill_2 FILLER_76_2127 ();
 sg13g2_fill_1 FILLER_76_2129 ();
 sg13g2_fill_1 FILLER_76_2161 ();
 sg13g2_fill_2 FILLER_76_2198 ();
 sg13g2_fill_1 FILLER_76_2200 ();
 sg13g2_fill_2 FILLER_76_2246 ();
 sg13g2_fill_2 FILLER_76_2324 ();
 sg13g2_fill_1 FILLER_76_2326 ();
 sg13g2_fill_2 FILLER_76_2337 ();
 sg13g2_fill_2 FILLER_76_2378 ();
 sg13g2_fill_1 FILLER_76_2380 ();
 sg13g2_fill_2 FILLER_76_2436 ();
 sg13g2_fill_1 FILLER_76_2438 ();
 sg13g2_fill_2 FILLER_76_2463 ();
 sg13g2_fill_2 FILLER_76_2501 ();
 sg13g2_fill_1 FILLER_76_2503 ();
 sg13g2_fill_2 FILLER_76_2534 ();
 sg13g2_fill_1 FILLER_76_2566 ();
 sg13g2_fill_2 FILLER_76_2585 ();
 sg13g2_fill_2 FILLER_76_2596 ();
 sg13g2_fill_2 FILLER_76_2634 ();
 sg13g2_fill_1 FILLER_76_2636 ();
 sg13g2_decap_8 FILLER_76_2646 ();
 sg13g2_decap_8 FILLER_76_2653 ();
 sg13g2_decap_8 FILLER_76_2660 ();
 sg13g2_decap_8 FILLER_76_2667 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_16 ();
 sg13g2_fill_1 FILLER_77_95 ();
 sg13g2_fill_2 FILLER_77_111 ();
 sg13g2_fill_1 FILLER_77_127 ();
 sg13g2_fill_2 FILLER_77_135 ();
 sg13g2_fill_1 FILLER_77_232 ();
 sg13g2_fill_2 FILLER_77_273 ();
 sg13g2_fill_2 FILLER_77_344 ();
 sg13g2_fill_1 FILLER_77_365 ();
 sg13g2_fill_1 FILLER_77_411 ();
 sg13g2_fill_2 FILLER_77_438 ();
 sg13g2_fill_2 FILLER_77_551 ();
 sg13g2_fill_1 FILLER_77_563 ();
 sg13g2_fill_2 FILLER_77_660 ();
 sg13g2_fill_1 FILLER_77_679 ();
 sg13g2_fill_2 FILLER_77_689 ();
 sg13g2_fill_1 FILLER_77_755 ();
 sg13g2_fill_1 FILLER_77_763 ();
 sg13g2_fill_2 FILLER_77_779 ();
 sg13g2_fill_2 FILLER_77_853 ();
 sg13g2_fill_1 FILLER_77_868 ();
 sg13g2_fill_1 FILLER_77_966 ();
 sg13g2_fill_1 FILLER_77_993 ();
 sg13g2_fill_2 FILLER_77_1014 ();
 sg13g2_fill_1 FILLER_77_1072 ();
 sg13g2_fill_1 FILLER_77_1078 ();
 sg13g2_fill_1 FILLER_77_1096 ();
 sg13g2_fill_2 FILLER_77_1123 ();
 sg13g2_fill_1 FILLER_77_1125 ();
 sg13g2_fill_2 FILLER_77_1210 ();
 sg13g2_fill_1 FILLER_77_1212 ();
 sg13g2_fill_1 FILLER_77_1220 ();
 sg13g2_fill_2 FILLER_77_1247 ();
 sg13g2_decap_4 FILLER_77_1281 ();
 sg13g2_decap_8 FILLER_77_1289 ();
 sg13g2_decap_8 FILLER_77_1296 ();
 sg13g2_fill_1 FILLER_77_1303 ();
 sg13g2_decap_4 FILLER_77_1340 ();
 sg13g2_fill_2 FILLER_77_1344 ();
 sg13g2_decap_8 FILLER_77_1351 ();
 sg13g2_decap_4 FILLER_77_1358 ();
 sg13g2_decap_4 FILLER_77_1375 ();
 sg13g2_fill_1 FILLER_77_1379 ();
 sg13g2_decap_4 FILLER_77_1390 ();
 sg13g2_fill_2 FILLER_77_1420 ();
 sg13g2_fill_1 FILLER_77_1422 ();
 sg13g2_fill_2 FILLER_77_1469 ();
 sg13g2_fill_1 FILLER_77_1499 ();
 sg13g2_fill_2 FILLER_77_1574 ();
 sg13g2_fill_2 FILLER_77_1602 ();
 sg13g2_fill_1 FILLER_77_1657 ();
 sg13g2_decap_8 FILLER_77_1728 ();
 sg13g2_decap_8 FILLER_77_1735 ();
 sg13g2_decap_8 FILLER_77_1742 ();
 sg13g2_decap_8 FILLER_77_1749 ();
 sg13g2_decap_4 FILLER_77_1756 ();
 sg13g2_fill_2 FILLER_77_1760 ();
 sg13g2_fill_1 FILLER_77_1766 ();
 sg13g2_decap_4 FILLER_77_1787 ();
 sg13g2_fill_2 FILLER_77_1798 ();
 sg13g2_fill_1 FILLER_77_1824 ();
 sg13g2_fill_1 FILLER_77_1833 ();
 sg13g2_decap_8 FILLER_77_1839 ();
 sg13g2_fill_1 FILLER_77_1846 ();
 sg13g2_decap_4 FILLER_77_1865 ();
 sg13g2_fill_2 FILLER_77_1869 ();
 sg13g2_decap_4 FILLER_77_1892 ();
 sg13g2_fill_1 FILLER_77_1896 ();
 sg13g2_fill_2 FILLER_77_1909 ();
 sg13g2_decap_4 FILLER_77_1916 ();
 sg13g2_fill_2 FILLER_77_1928 ();
 sg13g2_fill_1 FILLER_77_1930 ();
 sg13g2_fill_1 FILLER_77_1957 ();
 sg13g2_decap_8 FILLER_77_1986 ();
 sg13g2_decap_4 FILLER_77_1993 ();
 sg13g2_decap_8 FILLER_77_2018 ();
 sg13g2_fill_1 FILLER_77_2025 ();
 sg13g2_fill_2 FILLER_77_2049 ();
 sg13g2_fill_1 FILLER_77_2055 ();
 sg13g2_fill_1 FILLER_77_2061 ();
 sg13g2_fill_2 FILLER_77_2079 ();
 sg13g2_fill_1 FILLER_77_2081 ();
 sg13g2_fill_2 FILLER_77_2087 ();
 sg13g2_fill_1 FILLER_77_2089 ();
 sg13g2_fill_2 FILLER_77_2179 ();
 sg13g2_fill_1 FILLER_77_2181 ();
 sg13g2_fill_2 FILLER_77_2218 ();
 sg13g2_fill_1 FILLER_77_2220 ();
 sg13g2_fill_2 FILLER_77_2278 ();
 sg13g2_fill_1 FILLER_77_2280 ();
 sg13g2_fill_2 FILLER_77_2312 ();
 sg13g2_fill_1 FILLER_77_2327 ();
 sg13g2_fill_1 FILLER_77_2338 ();
 sg13g2_fill_1 FILLER_77_2391 ();
 sg13g2_fill_1 FILLER_77_2440 ();
 sg13g2_fill_1 FILLER_77_2512 ();
 sg13g2_fill_2 FILLER_77_2604 ();
 sg13g2_decap_8 FILLER_77_2627 ();
 sg13g2_fill_1 FILLER_77_2634 ();
 sg13g2_decap_8 FILLER_77_2639 ();
 sg13g2_decap_8 FILLER_77_2646 ();
 sg13g2_decap_8 FILLER_77_2653 ();
 sg13g2_decap_8 FILLER_77_2660 ();
 sg13g2_decap_8 FILLER_77_2667 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_114 ();
 sg13g2_fill_2 FILLER_78_139 ();
 sg13g2_fill_1 FILLER_78_158 ();
 sg13g2_fill_1 FILLER_78_172 ();
 sg13g2_fill_1 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_318 ();
 sg13g2_fill_2 FILLER_78_327 ();
 sg13g2_fill_2 FILLER_78_534 ();
 sg13g2_fill_1 FILLER_78_555 ();
 sg13g2_fill_2 FILLER_78_643 ();
 sg13g2_fill_1 FILLER_78_715 ();
 sg13g2_fill_2 FILLER_78_768 ();
 sg13g2_fill_1 FILLER_78_779 ();
 sg13g2_fill_2 FILLER_78_852 ();
 sg13g2_fill_1 FILLER_78_854 ();
 sg13g2_fill_2 FILLER_78_884 ();
 sg13g2_fill_1 FILLER_78_899 ();
 sg13g2_fill_2 FILLER_78_914 ();
 sg13g2_fill_1 FILLER_78_916 ();
 sg13g2_fill_2 FILLER_78_922 ();
 sg13g2_fill_2 FILLER_78_938 ();
 sg13g2_fill_1 FILLER_78_940 ();
 sg13g2_fill_2 FILLER_78_972 ();
 sg13g2_fill_1 FILLER_78_974 ();
 sg13g2_fill_2 FILLER_78_988 ();
 sg13g2_fill_1 FILLER_78_990 ();
 sg13g2_fill_2 FILLER_78_1040 ();
 sg13g2_fill_1 FILLER_78_1042 ();
 sg13g2_fill_1 FILLER_78_1052 ();
 sg13g2_fill_1 FILLER_78_1058 ();
 sg13g2_fill_2 FILLER_78_1074 ();
 sg13g2_fill_2 FILLER_78_1119 ();
 sg13g2_fill_1 FILLER_78_1121 ();
 sg13g2_fill_2 FILLER_78_1130 ();
 sg13g2_fill_1 FILLER_78_1144 ();
 sg13g2_fill_2 FILLER_78_1149 ();
 sg13g2_fill_1 FILLER_78_1151 ();
 sg13g2_fill_1 FILLER_78_1229 ();
 sg13g2_fill_2 FILLER_78_1243 ();
 sg13g2_fill_2 FILLER_78_1275 ();
 sg13g2_fill_1 FILLER_78_1277 ();
 sg13g2_fill_2 FILLER_78_1298 ();
 sg13g2_fill_2 FILLER_78_1317 ();
 sg13g2_fill_1 FILLER_78_1319 ();
 sg13g2_fill_1 FILLER_78_1374 ();
 sg13g2_fill_1 FILLER_78_1401 ();
 sg13g2_fill_1 FILLER_78_1428 ();
 sg13g2_fill_1 FILLER_78_1453 ();
 sg13g2_fill_1 FILLER_78_1462 ();
 sg13g2_fill_1 FILLER_78_1493 ();
 sg13g2_fill_1 FILLER_78_1518 ();
 sg13g2_fill_2 FILLER_78_1551 ();
 sg13g2_fill_1 FILLER_78_1584 ();
 sg13g2_fill_2 FILLER_78_1634 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_4 FILLER_78_1800 ();
 sg13g2_decap_4 FILLER_78_1818 ();
 sg13g2_fill_2 FILLER_78_1830 ();
 sg13g2_decap_8 FILLER_78_1850 ();
 sg13g2_fill_2 FILLER_78_1857 ();
 sg13g2_fill_2 FILLER_78_1864 ();
 sg13g2_fill_1 FILLER_78_1871 ();
 sg13g2_fill_2 FILLER_78_1877 ();
 sg13g2_decap_8 FILLER_78_1884 ();
 sg13g2_decap_8 FILLER_78_1891 ();
 sg13g2_fill_1 FILLER_78_1898 ();
 sg13g2_fill_2 FILLER_78_1912 ();
 sg13g2_fill_2 FILLER_78_1922 ();
 sg13g2_decap_4 FILLER_78_1936 ();
 sg13g2_fill_2 FILLER_78_1940 ();
 sg13g2_decap_8 FILLER_78_1951 ();
 sg13g2_decap_8 FILLER_78_1958 ();
 sg13g2_fill_2 FILLER_78_1984 ();
 sg13g2_decap_4 FILLER_78_1994 ();
 sg13g2_fill_2 FILLER_78_1998 ();
 sg13g2_fill_2 FILLER_78_2017 ();
 sg13g2_fill_1 FILLER_78_2019 ();
 sg13g2_fill_1 FILLER_78_2032 ();
 sg13g2_fill_1 FILLER_78_2051 ();
 sg13g2_fill_2 FILLER_78_2060 ();
 sg13g2_fill_2 FILLER_78_2098 ();
 sg13g2_fill_2 FILLER_78_2133 ();
 sg13g2_fill_1 FILLER_78_2171 ();
 sg13g2_fill_1 FILLER_78_2211 ();
 sg13g2_fill_2 FILLER_78_2292 ();
 sg13g2_fill_1 FILLER_78_2360 ();
 sg13g2_fill_1 FILLER_78_2387 ();
 sg13g2_fill_2 FILLER_78_2397 ();
 sg13g2_fill_1 FILLER_78_2399 ();
 sg13g2_fill_2 FILLER_78_2452 ();
 sg13g2_fill_2 FILLER_78_2484 ();
 sg13g2_fill_1 FILLER_78_2486 ();
 sg13g2_fill_2 FILLER_78_2517 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_4 FILLER_78_2670 ();
 sg13g2_decap_4 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_fill_1 FILLER_79_148 ();
 sg13g2_fill_2 FILLER_79_179 ();
 sg13g2_fill_1 FILLER_79_297 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_fill_2 FILLER_79_402 ();
 sg13g2_fill_1 FILLER_79_550 ();
 sg13g2_fill_1 FILLER_79_569 ();
 sg13g2_fill_1 FILLER_79_584 ();
 sg13g2_fill_1 FILLER_79_691 ();
 sg13g2_fill_2 FILLER_79_700 ();
 sg13g2_fill_2 FILLER_79_720 ();
 sg13g2_fill_2 FILLER_79_762 ();
 sg13g2_fill_1 FILLER_79_860 ();
 sg13g2_fill_2 FILLER_79_908 ();
 sg13g2_fill_1 FILLER_79_910 ();
 sg13g2_fill_1 FILLER_79_951 ();
 sg13g2_fill_2 FILLER_79_1058 ();
 sg13g2_decap_8 FILLER_79_1134 ();
 sg13g2_decap_8 FILLER_79_1145 ();
 sg13g2_fill_2 FILLER_79_1152 ();
 sg13g2_fill_1 FILLER_79_1154 ();
 sg13g2_fill_2 FILLER_79_1307 ();
 sg13g2_fill_2 FILLER_79_1351 ();
 sg13g2_fill_1 FILLER_79_1376 ();
 sg13g2_decap_4 FILLER_79_1390 ();
 sg13g2_fill_2 FILLER_79_1394 ();
 sg13g2_fill_2 FILLER_79_1477 ();
 sg13g2_fill_2 FILLER_79_1492 ();
 sg13g2_fill_2 FILLER_79_1548 ();
 sg13g2_decap_8 FILLER_79_1725 ();
 sg13g2_decap_8 FILLER_79_1732 ();
 sg13g2_decap_8 FILLER_79_1739 ();
 sg13g2_decap_4 FILLER_79_1746 ();
 sg13g2_fill_2 FILLER_79_1750 ();
 sg13g2_fill_2 FILLER_79_1779 ();
 sg13g2_fill_1 FILLER_79_1781 ();
 sg13g2_fill_1 FILLER_79_1839 ();
 sg13g2_fill_1 FILLER_79_1844 ();
 sg13g2_decap_8 FILLER_79_1884 ();
 sg13g2_fill_1 FILLER_79_1891 ();
 sg13g2_fill_2 FILLER_79_1971 ();
 sg13g2_fill_1 FILLER_79_1973 ();
 sg13g2_fill_2 FILLER_79_1982 ();
 sg13g2_fill_1 FILLER_79_2016 ();
 sg13g2_fill_1 FILLER_79_2035 ();
 sg13g2_decap_4 FILLER_79_2040 ();
 sg13g2_fill_2 FILLER_79_2044 ();
 sg13g2_fill_2 FILLER_79_2050 ();
 sg13g2_fill_2 FILLER_79_2056 ();
 sg13g2_fill_1 FILLER_79_2058 ();
 sg13g2_fill_2 FILLER_79_2069 ();
 sg13g2_fill_2 FILLER_79_2110 ();
 sg13g2_fill_2 FILLER_79_2117 ();
 sg13g2_fill_1 FILLER_79_2119 ();
 sg13g2_fill_1 FILLER_79_2146 ();
 sg13g2_fill_1 FILLER_79_2166 ();
 sg13g2_fill_2 FILLER_79_2204 ();
 sg13g2_fill_1 FILLER_79_2206 ();
 sg13g2_fill_2 FILLER_79_2269 ();
 sg13g2_fill_2 FILLER_79_2311 ();
 sg13g2_fill_2 FILLER_79_2371 ();
 sg13g2_fill_2 FILLER_79_2413 ();
 sg13g2_fill_1 FILLER_79_2415 ();
 sg13g2_fill_2 FILLER_79_2433 ();
 sg13g2_fill_2 FILLER_79_2468 ();
 sg13g2_fill_2 FILLER_79_2499 ();
 sg13g2_fill_1 FILLER_79_2501 ();
 sg13g2_fill_2 FILLER_79_2543 ();
 sg13g2_fill_1 FILLER_79_2545 ();
 sg13g2_fill_2 FILLER_79_2566 ();
 sg13g2_decap_8 FILLER_79_2598 ();
 sg13g2_decap_8 FILLER_79_2605 ();
 sg13g2_decap_8 FILLER_79_2612 ();
 sg13g2_decap_8 FILLER_79_2619 ();
 sg13g2_decap_8 FILLER_79_2626 ();
 sg13g2_decap_8 FILLER_79_2633 ();
 sg13g2_decap_8 FILLER_79_2640 ();
 sg13g2_decap_8 FILLER_79_2647 ();
 sg13g2_decap_8 FILLER_79_2654 ();
 sg13g2_decap_8 FILLER_79_2661 ();
 sg13g2_decap_4 FILLER_79_2668 ();
 sg13g2_fill_2 FILLER_79_2672 ();
 sg13g2_fill_2 FILLER_80_105 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_2 FILLER_80_150 ();
 sg13g2_fill_2 FILLER_80_247 ();
 sg13g2_fill_2 FILLER_80_323 ();
 sg13g2_fill_2 FILLER_80_338 ();
 sg13g2_fill_1 FILLER_80_446 ();
 sg13g2_fill_1 FILLER_80_585 ();
 sg13g2_fill_1 FILLER_80_643 ();
 sg13g2_fill_1 FILLER_80_677 ();
 sg13g2_fill_1 FILLER_80_734 ();
 sg13g2_fill_2 FILLER_80_761 ();
 sg13g2_fill_1 FILLER_80_856 ();
 sg13g2_fill_1 FILLER_80_929 ();
 sg13g2_fill_1 FILLER_80_969 ();
 sg13g2_fill_2 FILLER_80_987 ();
 sg13g2_fill_1 FILLER_80_989 ();
 sg13g2_fill_2 FILLER_80_1004 ();
 sg13g2_fill_1 FILLER_80_1006 ();
 sg13g2_fill_2 FILLER_80_1024 ();
 sg13g2_fill_1 FILLER_80_1026 ();
 sg13g2_decap_4 FILLER_80_1136 ();
 sg13g2_fill_1 FILLER_80_1174 ();
 sg13g2_fill_1 FILLER_80_1211 ();
 sg13g2_decap_8 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1252 ();
 sg13g2_decap_8 FILLER_80_1259 ();
 sg13g2_decap_8 FILLER_80_1274 ();
 sg13g2_decap_4 FILLER_80_1285 ();
 sg13g2_fill_2 FILLER_80_1297 ();
 sg13g2_fill_1 FILLER_80_1299 ();
 sg13g2_fill_2 FILLER_80_1313 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_decap_8 FILLER_80_1333 ();
 sg13g2_decap_4 FILLER_80_1340 ();
 sg13g2_fill_2 FILLER_80_1344 ();
 sg13g2_fill_2 FILLER_80_1354 ();
 sg13g2_fill_1 FILLER_80_1356 ();
 sg13g2_fill_2 FILLER_80_1362 ();
 sg13g2_fill_2 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1379 ();
 sg13g2_decap_8 FILLER_80_1386 ();
 sg13g2_decap_4 FILLER_80_1393 ();
 sg13g2_fill_1 FILLER_80_1397 ();
 sg13g2_fill_2 FILLER_80_1415 ();
 sg13g2_fill_1 FILLER_80_1417 ();
 sg13g2_fill_2 FILLER_80_1467 ();
 sg13g2_fill_1 FILLER_80_1469 ();
 sg13g2_fill_2 FILLER_80_1519 ();
 sg13g2_fill_2 FILLER_80_1570 ();
 sg13g2_fill_1 FILLER_80_1654 ();
 sg13g2_decap_8 FILLER_80_1728 ();
 sg13g2_decap_8 FILLER_80_1735 ();
 sg13g2_decap_8 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1749 ();
 sg13g2_fill_1 FILLER_80_1756 ();
 sg13g2_decap_8 FILLER_80_1767 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_4 FILLER_80_1788 ();
 sg13g2_fill_1 FILLER_80_1792 ();
 sg13g2_decap_4 FILLER_80_1797 ();
 sg13g2_fill_1 FILLER_80_1801 ();
 sg13g2_decap_8 FILLER_80_1806 ();
 sg13g2_fill_2 FILLER_80_1813 ();
 sg13g2_decap_4 FILLER_80_1819 ();
 sg13g2_fill_2 FILLER_80_1827 ();
 sg13g2_decap_4 FILLER_80_1855 ();
 sg13g2_fill_1 FILLER_80_1859 ();
 sg13g2_decap_4 FILLER_80_1864 ();
 sg13g2_fill_1 FILLER_80_1868 ();
 sg13g2_fill_2 FILLER_80_1895 ();
 sg13g2_fill_1 FILLER_80_1897 ();
 sg13g2_decap_4 FILLER_80_1903 ();
 sg13g2_fill_2 FILLER_80_1938 ();
 sg13g2_fill_1 FILLER_80_1940 ();
 sg13g2_fill_1 FILLER_80_1945 ();
 sg13g2_decap_8 FILLER_80_1980 ();
 sg13g2_fill_2 FILLER_80_1987 ();
 sg13g2_decap_8 FILLER_80_2015 ();
 sg13g2_fill_2 FILLER_80_2022 ();
 sg13g2_fill_1 FILLER_80_2024 ();
 sg13g2_decap_4 FILLER_80_2051 ();
 sg13g2_fill_2 FILLER_80_2055 ();
 sg13g2_fill_2 FILLER_80_2083 ();
 sg13g2_fill_2 FILLER_80_2147 ();
 sg13g2_fill_2 FILLER_80_2193 ();
 sg13g2_fill_1 FILLER_80_2195 ();
 sg13g2_fill_2 FILLER_80_2286 ();
 sg13g2_fill_2 FILLER_80_2314 ();
 sg13g2_fill_1 FILLER_80_2316 ();
 sg13g2_fill_2 FILLER_80_2377 ();
 sg13g2_fill_1 FILLER_80_2379 ();
 sg13g2_fill_2 FILLER_80_2390 ();
 sg13g2_fill_2 FILLER_80_2439 ();
 sg13g2_fill_2 FILLER_80_2519 ();
 sg13g2_fill_2 FILLER_80_2555 ();
 sg13g2_decap_8 FILLER_80_2596 ();
 sg13g2_decap_8 FILLER_80_2603 ();
 sg13g2_decap_8 FILLER_80_2610 ();
 sg13g2_decap_8 FILLER_80_2617 ();
 sg13g2_decap_8 FILLER_80_2624 ();
 sg13g2_decap_8 FILLER_80_2631 ();
 sg13g2_decap_8 FILLER_80_2638 ();
 sg13g2_decap_8 FILLER_80_2645 ();
 sg13g2_decap_8 FILLER_80_2652 ();
 sg13g2_decap_8 FILLER_80_2659 ();
 sg13g2_decap_8 FILLER_80_2666 ();
 sg13g2_fill_1 FILLER_80_2673 ();
 assign uio_oe[0] = net2923;
 assign uio_oe[3] = net2924;
 assign uio_oe[6] = net2925;
 assign uio_oe[7] = net2926;
 assign uio_out[6] = net2927;
endmodule
