module tt_um_rejunity_lgn_mnist (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire \calc_categories[0].sum_bits.popcount128.ad0.genblk1[105].add3.a ;
 wire \calc_categories[4].sum_bits.popcount128.add3.genblk1[12].add3.c ;
 wire \calc_categories[6].sum_bits.popcount128.ad0.genblk1[108].add3.a ;
 wire \net.in[0] ;
 wire \net.in[100] ;
 wire \net.in[101] ;
 wire \net.in[102] ;
 wire \net.in[103] ;
 wire \net.in[104] ;
 wire \net.in[105] ;
 wire \net.in[106] ;
 wire \net.in[107] ;
 wire \net.in[108] ;
 wire \net.in[109] ;
 wire \net.in[10] ;
 wire \net.in[110] ;
 wire \net.in[111] ;
 wire \net.in[112] ;
 wire \net.in[113] ;
 wire \net.in[114] ;
 wire \net.in[115] ;
 wire \net.in[116] ;
 wire \net.in[117] ;
 wire \net.in[118] ;
 wire \net.in[119] ;
 wire \net.in[11] ;
 wire \net.in[120] ;
 wire \net.in[121] ;
 wire \net.in[122] ;
 wire \net.in[123] ;
 wire \net.in[124] ;
 wire \net.in[125] ;
 wire \net.in[126] ;
 wire \net.in[127] ;
 wire \net.in[128] ;
 wire \net.in[129] ;
 wire \net.in[130] ;
 wire \net.in[131] ;
 wire \net.in[132] ;
 wire \net.in[133] ;
 wire \net.in[134] ;
 wire \net.in[135] ;
 wire \net.in[136] ;
 wire \net.in[137] ;
 wire \net.in[138] ;
 wire \net.in[139] ;
 wire \net.in[13] ;
 wire \net.in[140] ;
 wire \net.in[141] ;
 wire \net.in[143] ;
 wire \net.in[144] ;
 wire \net.in[145] ;
 wire \net.in[146] ;
 wire \net.in[147] ;
 wire \net.in[148] ;
 wire \net.in[149] ;
 wire \net.in[14] ;
 wire \net.in[150] ;
 wire \net.in[151] ;
 wire \net.in[152] ;
 wire \net.in[154] ;
 wire \net.in[155] ;
 wire \net.in[156] ;
 wire \net.in[157] ;
 wire \net.in[158] ;
 wire \net.in[159] ;
 wire \net.in[15] ;
 wire \net.in[160] ;
 wire \net.in[161] ;
 wire \net.in[162] ;
 wire \net.in[163] ;
 wire \net.in[164] ;
 wire \net.in[165] ;
 wire \net.in[166] ;
 wire \net.in[167] ;
 wire \net.in[168] ;
 wire \net.in[169] ;
 wire \net.in[16] ;
 wire \net.in[170] ;
 wire \net.in[171] ;
 wire \net.in[172] ;
 wire \net.in[173] ;
 wire \net.in[174] ;
 wire \net.in[175] ;
 wire \net.in[176] ;
 wire \net.in[177] ;
 wire \net.in[178] ;
 wire \net.in[179] ;
 wire \net.in[17] ;
 wire \net.in[180] ;
 wire \net.in[181] ;
 wire \net.in[182] ;
 wire \net.in[183] ;
 wire \net.in[184] ;
 wire \net.in[185] ;
 wire \net.in[186] ;
 wire \net.in[187] ;
 wire \net.in[188] ;
 wire \net.in[189] ;
 wire \net.in[18] ;
 wire \net.in[190] ;
 wire \net.in[191] ;
 wire \net.in[192] ;
 wire \net.in[193] ;
 wire \net.in[194] ;
 wire \net.in[195] ;
 wire \net.in[196] ;
 wire \net.in[197] ;
 wire \net.in[198] ;
 wire \net.in[199] ;
 wire \net.in[19] ;
 wire \net.in[1] ;
 wire \net.in[200] ;
 wire \net.in[201] ;
 wire \net.in[202] ;
 wire \net.in[203] ;
 wire \net.in[204] ;
 wire \net.in[205] ;
 wire \net.in[206] ;
 wire \net.in[207] ;
 wire \net.in[208] ;
 wire \net.in[209] ;
 wire \net.in[20] ;
 wire \net.in[210] ;
 wire \net.in[211] ;
 wire \net.in[212] ;
 wire \net.in[213] ;
 wire \net.in[214] ;
 wire \net.in[215] ;
 wire \net.in[216] ;
 wire \net.in[217] ;
 wire \net.in[218] ;
 wire \net.in[219] ;
 wire \net.in[21] ;
 wire \net.in[220] ;
 wire \net.in[221] ;
 wire \net.in[222] ;
 wire \net.in[223] ;
 wire \net.in[224] ;
 wire \net.in[225] ;
 wire \net.in[226] ;
 wire \net.in[227] ;
 wire \net.in[228] ;
 wire \net.in[229] ;
 wire \net.in[22] ;
 wire \net.in[230] ;
 wire \net.in[231] ;
 wire \net.in[232] ;
 wire \net.in[233] ;
 wire \net.in[234] ;
 wire \net.in[235] ;
 wire \net.in[236] ;
 wire \net.in[237] ;
 wire \net.in[238] ;
 wire \net.in[239] ;
 wire \net.in[23] ;
 wire \net.in[240] ;
 wire \net.in[241] ;
 wire \net.in[242] ;
 wire \net.in[243] ;
 wire \net.in[244] ;
 wire \net.in[245] ;
 wire \net.in[246] ;
 wire \net.in[247] ;
 wire \net.in[248] ;
 wire \net.in[249] ;
 wire \net.in[24] ;
 wire \net.in[250] ;
 wire \net.in[251] ;
 wire \net.in[252] ;
 wire \net.in[253] ;
 wire \net.in[25] ;
 wire \net.in[26] ;
 wire \net.in[27] ;
 wire \net.in[28] ;
 wire \net.in[29] ;
 wire \net.in[2] ;
 wire \net.in[30] ;
 wire \net.in[31] ;
 wire \net.in[32] ;
 wire \net.in[33] ;
 wire \net.in[34] ;
 wire \net.in[35] ;
 wire \net.in[36] ;
 wire \net.in[37] ;
 wire \net.in[38] ;
 wire \net.in[39] ;
 wire \net.in[3] ;
 wire \net.in[40] ;
 wire \net.in[41] ;
 wire \net.in[42] ;
 wire \net.in[43] ;
 wire \net.in[44] ;
 wire \net.in[45] ;
 wire \net.in[46] ;
 wire \net.in[47] ;
 wire \net.in[48] ;
 wire \net.in[49] ;
 wire \net.in[4] ;
 wire \net.in[50] ;
 wire \net.in[51] ;
 wire \net.in[52] ;
 wire \net.in[53] ;
 wire \net.in[54] ;
 wire \net.in[55] ;
 wire \net.in[56] ;
 wire \net.in[57] ;
 wire \net.in[58] ;
 wire \net.in[59] ;
 wire \net.in[5] ;
 wire \net.in[60] ;
 wire \net.in[61] ;
 wire \net.in[62] ;
 wire \net.in[63] ;
 wire \net.in[64] ;
 wire \net.in[65] ;
 wire \net.in[66] ;
 wire \net.in[67] ;
 wire \net.in[68] ;
 wire \net.in[69] ;
 wire \net.in[6] ;
 wire \net.in[70] ;
 wire \net.in[71] ;
 wire \net.in[72] ;
 wire \net.in[73] ;
 wire \net.in[74] ;
 wire \net.in[75] ;
 wire \net.in[76] ;
 wire \net.in[77] ;
 wire \net.in[78] ;
 wire \net.in[79] ;
 wire \net.in[7] ;
 wire \net.in[80] ;
 wire \net.in[81] ;
 wire \net.in[82] ;
 wire \net.in[83] ;
 wire \net.in[84] ;
 wire \net.in[85] ;
 wire \net.in[86] ;
 wire \net.in[87] ;
 wire \net.in[88] ;
 wire \net.in[89] ;
 wire \net.in[8] ;
 wire \net.in[90] ;
 wire \net.in[91] ;
 wire \net.in[92] ;
 wire \net.in[93] ;
 wire \net.in[94] ;
 wire \net.in[95] ;
 wire \net.in[96] ;
 wire \net.in[97] ;
 wire \net.in[98] ;
 wire \net.in[99] ;
 wire \net.in[9] ;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire clknet_leaf_0_clk;
 wire net11;
 wire net12;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;

 sg13g2_inv_2 _10349_ (.Y(_05000_),
    .A(\net.in[133] ));
 sg13g2_inv_2 _10350_ (.Y(_05011_),
    .A(net2699));
 sg13g2_inv_4 _10351_ (.A(net2430),
    .Y(_05022_));
 sg13g2_inv_1 _10352_ (.Y(_05033_),
    .A(net2522));
 sg13g2_inv_8 _10353_ (.Y(_05044_),
    .A(net2472));
 sg13g2_inv_2 _10354_ (.Y(_05055_),
    .A(net2259));
 sg13g2_inv_8 _10355_ (.Y(_05066_),
    .A(net2307));
 sg13g2_inv_4 _10356_ (.A(net2295),
    .Y(_05077_));
 sg13g2_inv_4 _10357_ (.A(net2499),
    .Y(_05088_));
 sg13g2_inv_8 _10358_ (.Y(_05099_),
    .A(net318));
 sg13g2_inv_1 _10359_ (.Y(_05110_),
    .A(net2241));
 sg13g2_inv_8 _10360_ (.Y(_05121_),
    .A(net2345));
 sg13g2_inv_2 _10361_ (.Y(_05132_),
    .A(net2219));
 sg13g2_inv_4 _10362_ (.A(net2765),
    .Y(_05143_));
 sg13g2_inv_8 _10363_ (.Y(_05154_),
    .A(net2806));
 sg13g2_inv_2 _10364_ (.Y(_05165_),
    .A(net2506));
 sg13g2_inv_8 _10365_ (.Y(_05176_),
    .A(net2554));
 sg13g2_inv_8 _10366_ (.Y(_05187_),
    .A(net2467));
 sg13g2_inv_1 _10367_ (.Y(_05198_),
    .A(net2519));
 sg13g2_inv_8 _10368_ (.Y(_05209_),
    .A(net2340));
 sg13g2_inv_4 _10369_ (.A(net2559),
    .Y(_05220_));
 sg13g2_inv_1 _10370_ (.Y(_05231_),
    .A(net2613));
 sg13g2_inv_2 _10371_ (.Y(_05242_),
    .A(net2528));
 sg13g2_inv_8 _10372_ (.Y(_05253_),
    .A(net2186));
 sg13g2_inv_4 _10373_ (.A(net2424),
    .Y(_05264_));
 sg13g2_inv_4 _10374_ (.A(net354),
    .Y(_05275_));
 sg13g2_inv_2 _10375_ (.Y(_05286_),
    .A(\net.in[149] ));
 sg13g2_inv_8 _10376_ (.Y(_05297_),
    .A(net2442));
 sg13g2_inv_4 _10377_ (.A(net2391),
    .Y(_05308_));
 sg13g2_inv_4 _10378_ (.A(net2312),
    .Y(_05319_));
 sg13g2_inv_8 _10379_ (.Y(_05330_),
    .A(net2557));
 sg13g2_inv_1 _10380_ (.Y(_05341_),
    .A(net2497));
 sg13g2_inv_8 _10381_ (.Y(_05352_),
    .A(net2414));
 sg13g2_inv_8 _10382_ (.Y(_05363_),
    .A(net2383));
 sg13g2_inv_4 _10383_ (.A(net2463),
    .Y(_05374_));
 sg13g2_inv_8 _10384_ (.Y(_05385_),
    .A(net2566));
 sg13g2_inv_2 _10385_ (.Y(_05396_),
    .A(net2192));
 sg13g2_inv_4 _10386_ (.A(net2447),
    .Y(_05407_));
 sg13g2_inv_8 _10387_ (.Y(_05418_),
    .A(net2439));
 sg13g2_inv_1 _10388_ (.Y(_05429_),
    .A(net2360));
 sg13g2_inv_2 _10389_ (.Y(_05440_),
    .A(\net.in[139] ));
 sg13g2_inv_8 _10390_ (.Y(_05451_),
    .A(net337));
 sg13g2_inv_8 _10391_ (.Y(_05462_),
    .A(net2379));
 sg13g2_inv_4 _10392_ (.A(net2356),
    .Y(_05473_));
 sg13g2_inv_8 _10393_ (.Y(_05484_),
    .A(net2293));
 sg13g2_inv_8 _10394_ (.Y(_05495_),
    .A(net2755));
 sg13g2_inv_8 _10395_ (.Y(_05506_),
    .A(\net.in[10] ));
 sg13g2_inv_1 _10396_ (.Y(_05517_),
    .A(net2224));
 sg13g2_inv_2 _10397_ (.Y(_05528_),
    .A(net2267));
 sg13g2_inv_4 _10398_ (.A(net2387),
    .Y(_05539_));
 sg13g2_inv_2 _10399_ (.Y(_05550_),
    .A(net2200));
 sg13g2_inv_8 _10400_ (.Y(_05561_),
    .A(net2710));
 sg13g2_inv_2 _10401_ (.Y(_05572_),
    .A(net2653));
 sg13g2_inv_1 _10402_ (.Y(_05583_),
    .A(net2189));
 sg13g2_inv_4 _10403_ (.A(net2631),
    .Y(_05594_));
 sg13g2_inv_1 _10404_ (.Y(_05605_),
    .A(net2196));
 sg13g2_inv_1 _10405_ (.Y(_05616_),
    .A(net2216));
 sg13g2_inv_2 _10406_ (.Y(_05627_),
    .A(net2770));
 sg13g2_inv_2 _10407_ (.Y(_05638_),
    .A(net2377));
 sg13g2_inv_1 _10408_ (.Y(_05649_),
    .A(net2759));
 sg13g2_inv_4 _10409_ (.A(net2795),
    .Y(_05660_));
 sg13g2_inv_1 _10410_ (.Y(_05671_),
    .A(net2489));
 sg13g2_inv_4 _10411_ (.A(net2589),
    .Y(_05682_));
 sg13g2_inv_8 _10412_ (.Y(_05693_),
    .A(net2581));
 sg13g2_inv_4 _10413_ (.A(net2223),
    .Y(_05704_));
 sg13g2_inv_4 _10414_ (.A(net2675),
    .Y(_05715_));
 sg13g2_inv_4 _10415_ (.A(net2636),
    .Y(_05726_));
 sg13g2_inv_4 _10416_ (.A(net2204),
    .Y(_05737_));
 sg13g2_inv_1 _10417_ (.Y(_05748_),
    .A(net2707));
 sg13g2_inv_1 _10418_ (.Y(_05759_),
    .A(net2230));
 sg13g2_inv_8 _10419_ (.Y(_05770_),
    .A(net2616));
 sg13g2_inv_1 _10420_ (.Y(_05781_),
    .A(net2369));
 sg13g2_inv_8 _10421_ (.Y(_05792_),
    .A(net2682));
 sg13g2_inv_2 _10422_ (.Y(_05803_),
    .A(net2328));
 sg13g2_inv_4 _10423_ (.A(net2563),
    .Y(_05814_));
 sg13g2_inv_1 _10424_ (.Y(_05825_),
    .A(net381));
 sg13g2_inv_4 _10425_ (.A(net2659),
    .Y(_05836_));
 sg13g2_inv_8 _10426_ (.Y(_05847_),
    .A(net2255));
 sg13g2_inv_4 _10427_ (.A(net2595),
    .Y(_05858_));
 sg13g2_inv_4 _10428_ (.A(net2784),
    .Y(_05869_));
 sg13g2_inv_1 _10429_ (.Y(_05880_),
    .A(net2648));
 sg13g2_inv_4 _10430_ (.A(net2746),
    .Y(_05891_));
 sg13g2_inv_1 _10431_ (.Y(_05902_),
    .A(\net.in[207] ));
 sg13g2_inv_8 _10432_ (.Y(_05913_),
    .A(net2791));
 sg13g2_inv_4 _10433_ (.A(\net.in[237] ),
    .Y(_05924_));
 sg13g2_inv_1 _10434_ (.Y(_05935_),
    .A(net2275));
 sg13g2_inv_8 _10435_ (.Y(_05946_),
    .A(net2739));
 sg13g2_inv_8 _10436_ (.Y(_05957_),
    .A(net2714));
 sg13g2_inv_4 _10437_ (.A(net2409),
    .Y(_05968_));
 sg13g2_inv_8 _10438_ (.Y(_05979_),
    .A(net2640));
 sg13g2_inv_1 _10439_ (.Y(_05990_),
    .A(net2287));
 sg13g2_inv_2 _10440_ (.Y(_06001_),
    .A(net2744));
 sg13g2_inv_4 _10441_ (.A(net2197),
    .Y(_06012_));
 sg13g2_inv_4 _10442_ (.A(net2761),
    .Y(_06023_));
 sg13g2_inv_2 _10443_ (.Y(_06034_),
    .A(net2210));
 sg13g2_inv_8 _10444_ (.Y(_06045_),
    .A(net2813));
 sg13g2_inv_2 _10445_ (.Y(_06056_),
    .A(net357));
 sg13g2_inv_1 _10446_ (.Y(_06067_),
    .A(\net.in[222] ));
 sg13g2_inv_4 _10447_ (.A(\net.in[31] ),
    .Y(_06078_));
 sg13g2_inv_1 _10448_ (.Y(_06089_),
    .A(_00013_));
 sg13g2_inv_1 _10449_ (.Y(_06100_),
    .A(_00015_));
 sg13g2_inv_1 _10450_ (.Y(_06111_),
    .A(_00017_));
 sg13g2_inv_1 _10451_ (.Y(_06122_),
    .A(_00020_));
 sg13g2_xnor2_1 _10452_ (.Y(_06133_),
    .A(net2463),
    .B(net2409));
 sg13g2_xor2_1 _10453_ (.B(\net.in[49] ),
    .A(net2550),
    .X(_06144_));
 sg13g2_nor2_2 _10454_ (.A(_06133_),
    .B(_06144_),
    .Y(_06155_));
 sg13g2_nor2_1 _10455_ (.A(net2531),
    .B(net2577),
    .Y(_06166_));
 sg13g2_xor2_1 _10456_ (.B(net2575),
    .A(net2530),
    .X(_06177_));
 sg13g2_xnor2_1 _10457_ (.Y(_06188_),
    .A(net2295),
    .B(net2231));
 sg13g2_nor2b_1 _10458_ (.A(net2732),
    .B_N(net2700),
    .Y(_06199_));
 sg13g2_xnor2_1 _10459_ (.Y(_06210_),
    .A(_06188_),
    .B(_06199_));
 sg13g2_nand2b_1 _10460_ (.Y(_06221_),
    .B(_06177_),
    .A_N(_06210_));
 sg13g2_nor2b_1 _10461_ (.A(_06177_),
    .B_N(_06210_),
    .Y(_06232_));
 sg13g2_xor2_1 _10462_ (.B(_06210_),
    .A(_06177_),
    .X(_06243_));
 sg13g2_xor2_1 _10463_ (.B(net2796),
    .A(net2769),
    .X(_06254_));
 sg13g2_xnor2_1 _10464_ (.Y(_06265_),
    .A(net2264),
    .B(net2704));
 sg13g2_xnor2_1 _10465_ (.Y(_06276_),
    .A(_06254_),
    .B(_06265_));
 sg13g2_xnor2_1 _10466_ (.Y(_06287_),
    .A(_06243_),
    .B(_06276_));
 sg13g2_xor2_1 _10467_ (.B(net2548),
    .A(net2760),
    .X(_06298_));
 sg13g2_xnor2_1 _10468_ (.Y(_06309_),
    .A(net2534),
    .B(net2496));
 sg13g2_nor2_1 _10469_ (.A(net2710),
    .B(net2757),
    .Y(_06320_));
 sg13g2_nor2_1 _10470_ (.A(net2752),
    .B(net2662),
    .Y(_06331_));
 sg13g2_xnor2_1 _10471_ (.Y(_06342_),
    .A(_06320_),
    .B(_06331_));
 sg13g2_nor2b_1 _10472_ (.A(_06309_),
    .B_N(_06342_),
    .Y(_06353_));
 sg13g2_nor2b_1 _10473_ (.A(_06342_),
    .B_N(_06309_),
    .Y(_06364_));
 sg13g2_xnor2_1 _10474_ (.Y(_06375_),
    .A(_06309_),
    .B(_06342_));
 sg13g2_xnor2_1 _10475_ (.Y(_06386_),
    .A(_06298_),
    .B(_06375_));
 sg13g2_nand2_1 _10476_ (.Y(_06397_),
    .A(_06287_),
    .B(_06386_));
 sg13g2_or2_1 _10477_ (.X(_06408_),
    .B(_06386_),
    .A(_06287_));
 sg13g2_xnor2_1 _10478_ (.Y(_06419_),
    .A(_06287_),
    .B(_06386_));
 sg13g2_xor2_1 _10479_ (.B(net2646),
    .A(net2699),
    .X(_06430_));
 sg13g2_nor2_1 _10480_ (.A(net2750),
    .B(net2787),
    .Y(_06441_));
 sg13g2_nor2_1 _10481_ (.A(net2301),
    .B(net2790),
    .Y(_06452_));
 sg13g2_xnor2_1 _10482_ (.Y(_06463_),
    .A(_06441_),
    .B(_06452_));
 sg13g2_nor2_1 _10483_ (.A(_06430_),
    .B(_06463_),
    .Y(_06474_));
 sg13g2_nand2_1 _10484_ (.Y(_06485_),
    .A(_06430_),
    .B(_06463_));
 sg13g2_nor2b_1 _10485_ (.A(_06474_),
    .B_N(_06485_),
    .Y(_06496_));
 sg13g2_xnor2_1 _10486_ (.Y(_06507_),
    .A(net2765),
    .B(net2690));
 sg13g2_or3_2 _10487_ (.A(net2256),
    .B(net2608),
    .C(_06507_),
    .X(_06518_));
 sg13g2_xnor2_1 _10488_ (.Y(_06529_),
    .A(_06496_),
    .B(_06518_));
 sg13g2_xnor2_1 _10489_ (.Y(_06540_),
    .A(_06419_),
    .B(_06529_));
 sg13g2_nor2_1 _10490_ (.A(net2583),
    .B(net2537),
    .Y(_06551_));
 sg13g2_xor2_1 _10491_ (.B(net2537),
    .A(net2583),
    .X(_06562_));
 sg13g2_xnor2_1 _10492_ (.Y(_06573_),
    .A(net2581),
    .B(net2534));
 sg13g2_xnor2_1 _10493_ (.Y(_06584_),
    .A(net2725),
    .B(net2790));
 sg13g2_xor2_1 _10494_ (.B(net2623),
    .A(net2447),
    .X(_06595_));
 sg13g2_xnor2_1 _10495_ (.Y(_06606_),
    .A(_06584_),
    .B(_06595_));
 sg13g2_nor2b_1 _10496_ (.A(net2796),
    .B_N(net2467),
    .Y(_06617_));
 sg13g2_xnor2_1 _10497_ (.Y(_06628_),
    .A(net2367),
    .B(net2502));
 sg13g2_xnor2_1 _10498_ (.Y(_06639_),
    .A(_06617_),
    .B(_06628_));
 sg13g2_nor2b_1 _10499_ (.A(_06606_),
    .B_N(_06639_),
    .Y(_06650_));
 sg13g2_nor2b_1 _10500_ (.A(_06639_),
    .B_N(_06606_),
    .Y(_06661_));
 sg13g2_xnor2_1 _10501_ (.Y(_06672_),
    .A(_06606_),
    .B(_06639_));
 sg13g2_xnor2_1 _10502_ (.Y(_06683_),
    .A(_06573_),
    .B(_06672_));
 sg13g2_nor2_1 _10503_ (.A(net2593),
    .B(net2545),
    .Y(_06694_));
 sg13g2_xor2_1 _10504_ (.B(net2547),
    .A(net2592),
    .X(_06705_));
 sg13g2_xnor2_1 _10505_ (.Y(_06716_),
    .A(net2729),
    .B(_06705_));
 sg13g2_xnor2_1 _10506_ (.Y(_06727_),
    .A(net2539),
    .B(net2496));
 sg13g2_xnor2_1 _10507_ (.Y(_06738_),
    .A(net2521),
    .B(net2437));
 sg13g2_nand2_1 _10508_ (.Y(_06749_),
    .A(_06727_),
    .B(_06738_));
 sg13g2_nor2_1 _10509_ (.A(_06727_),
    .B(_06738_),
    .Y(_06760_));
 sg13g2_xnor2_1 _10510_ (.Y(_06771_),
    .A(_06727_),
    .B(_06738_));
 sg13g2_xnor2_1 _10511_ (.Y(_06782_),
    .A(_06716_),
    .B(_06771_));
 sg13g2_nor2_1 _10512_ (.A(_06683_),
    .B(_06782_),
    .Y(_06793_));
 sg13g2_xor2_1 _10513_ (.B(_06782_),
    .A(_06683_),
    .X(_06804_));
 sg13g2_xor2_1 _10514_ (.B(net2642),
    .A(net2699),
    .X(_06815_));
 sg13g2_nor2_1 _10515_ (.A(_05022_),
    .B(net2787),
    .Y(_06826_));
 sg13g2_xor2_1 _10516_ (.B(net2447),
    .A(net2484),
    .X(_06837_));
 sg13g2_xor2_1 _10517_ (.B(net2255),
    .A(net2729),
    .X(_06848_));
 sg13g2_a21oi_2 _10518_ (.B1(_06848_),
    .Y(_06859_),
    .A2(_06837_),
    .A1(_06826_));
 sg13g2_inv_1 _10519_ (.Y(_06870_),
    .A(_06859_));
 sg13g2_and3_1 _10520_ (.X(_06881_),
    .A(_06826_),
    .B(_06837_),
    .C(_06848_));
 sg13g2_nor2_1 _10521_ (.A(_06859_),
    .B(_06881_),
    .Y(_06892_));
 sg13g2_xnor2_1 _10522_ (.Y(_06903_),
    .A(_06815_),
    .B(_06892_));
 sg13g2_xnor2_1 _10523_ (.Y(_06914_),
    .A(_06804_),
    .B(_06903_));
 sg13g2_nand2_1 _10524_ (.Y(_06925_),
    .A(_06540_),
    .B(_06914_));
 sg13g2_or2_1 _10525_ (.X(_06936_),
    .B(_06914_),
    .A(_06540_));
 sg13g2_nand2_1 _10526_ (.Y(_06947_),
    .A(_06925_),
    .B(_06936_));
 sg13g2_xnor2_1 _10527_ (.Y(_06958_),
    .A(_06155_),
    .B(_06947_));
 sg13g2_nor2_1 _10528_ (.A(net2221),
    .B(net2285),
    .Y(_06969_));
 sg13g2_xor2_1 _10529_ (.B(net2285),
    .A(net2220),
    .X(_06980_));
 sg13g2_xor2_1 _10530_ (.B(net2309),
    .A(net2357),
    .X(_06991_));
 sg13g2_nor2_1 _10531_ (.A(_06980_),
    .B(_06991_),
    .Y(_07002_));
 sg13g2_nor2_1 _10532_ (.A(net2602),
    .B(net2547),
    .Y(_07013_));
 sg13g2_nor2_1 _10533_ (.A(net2705),
    .B(net2320),
    .Y(_07024_));
 sg13g2_xor2_1 _10534_ (.B(net2460),
    .A(net2325),
    .X(_07035_));
 sg13g2_xnor2_1 _10535_ (.Y(_07046_),
    .A(_07024_),
    .B(_07035_));
 sg13g2_nor3_1 _10536_ (.A(net2214),
    .B(_07013_),
    .C(_07046_),
    .Y(_07057_));
 sg13g2_o21ai_1 _10537_ (.B1(_07046_),
    .Y(_07068_),
    .A1(net2214),
    .A2(_07013_));
 sg13g2_nand2b_1 _10538_ (.Y(_07079_),
    .B(_07068_),
    .A_N(_07057_));
 sg13g2_xnor2_1 _10539_ (.Y(_07090_),
    .A(_07002_),
    .B(_07079_));
 sg13g2_nor2_1 _10540_ (.A(net2502),
    .B(net2552),
    .Y(_07101_));
 sg13g2_a21oi_1 _10541_ (.A1(net2722),
    .A2(net2274),
    .Y(_07112_),
    .B1(_07101_));
 sg13g2_o21ai_1 _10542_ (.B1(_07112_),
    .Y(_07123_),
    .A1(net2722),
    .A2(net2274));
 sg13g2_nor3_2 _10543_ (.A(net2548),
    .B(\net.in[253] ),
    .C(_06111_),
    .Y(_07134_));
 sg13g2_xor2_1 _10544_ (.B(net2207),
    .A(net2259),
    .X(_07145_));
 sg13g2_xnor2_1 _10545_ (.Y(_07156_),
    .A(net2285),
    .B(_07145_));
 sg13g2_nor2b_1 _10546_ (.A(_07156_),
    .B_N(_07134_),
    .Y(_07167_));
 sg13g2_nand2b_1 _10547_ (.Y(_07178_),
    .B(_07156_),
    .A_N(_07134_));
 sg13g2_o21ai_1 _10548_ (.B1(_07178_),
    .Y(_07189_),
    .A1(_07123_),
    .A2(_07167_));
 sg13g2_xor2_1 _10549_ (.B(_07156_),
    .A(_07134_),
    .X(_07200_));
 sg13g2_xnor2_1 _10550_ (.Y(_07211_),
    .A(_07123_),
    .B(_07200_));
 sg13g2_nor2_1 _10551_ (.A(net2194),
    .B(_05957_),
    .Y(_07222_));
 sg13g2_nand2_1 _10552_ (.Y(_07233_),
    .A(net2694),
    .B(net2682));
 sg13g2_xnor2_1 _10553_ (.Y(_07244_),
    .A(_07222_),
    .B(_07233_));
 sg13g2_xnor2_1 _10554_ (.Y(_07255_),
    .A(net2513),
    .B(net2717));
 sg13g2_xnor2_1 _10555_ (.Y(_07266_),
    .A(net2218),
    .B(net2325));
 sg13g2_nand2_1 _10556_ (.Y(_07277_),
    .A(_07255_),
    .B(_07266_));
 sg13g2_nor2b_1 _10557_ (.A(net2764),
    .B_N(net2380),
    .Y(_07288_));
 sg13g2_nor2b_1 _10558_ (.A(net2602),
    .B_N(net2714),
    .Y(_07299_));
 sg13g2_xnor2_1 _10559_ (.Y(_07310_),
    .A(_07288_),
    .B(_07299_));
 sg13g2_nor2b_1 _10560_ (.A(_07277_),
    .B_N(_07310_),
    .Y(_07321_));
 sg13g2_a21o_1 _10561_ (.A2(_07266_),
    .A1(_07255_),
    .B1(_07310_),
    .X(_07332_));
 sg13g2_xor2_1 _10562_ (.B(_07310_),
    .A(_07277_),
    .X(_07343_));
 sg13g2_a21oi_2 _10563_ (.B1(_07321_),
    .Y(_07354_),
    .A2(_07332_),
    .A1(_07244_));
 sg13g2_xnor2_1 _10564_ (.Y(_07365_),
    .A(_07244_),
    .B(_07343_));
 sg13g2_inv_1 _10565_ (.Y(_07376_),
    .A(_07365_));
 sg13g2_nor2_1 _10566_ (.A(_07211_),
    .B(_07376_),
    .Y(_07387_));
 sg13g2_nand2_1 _10567_ (.Y(_07398_),
    .A(_07211_),
    .B(_07376_));
 sg13g2_xnor2_1 _10568_ (.Y(_07409_),
    .A(_07211_),
    .B(_07365_));
 sg13g2_xnor2_1 _10569_ (.Y(_07420_),
    .A(_07090_),
    .B(_07409_));
 sg13g2_xor2_1 _10570_ (.B(net2581),
    .A(net2530),
    .X(_07431_));
 sg13g2_nor3_2 _10571_ (.A(net2652),
    .B(net2548),
    .C(_07431_),
    .Y(_07442_));
 sg13g2_nor2_2 _10572_ (.A(\net.in[154] ),
    .B(net2369),
    .Y(_07453_));
 sg13g2_or2_1 _10573_ (.X(_07464_),
    .B(net2367),
    .A(net2416));
 sg13g2_xnor2_1 _10574_ (.Y(_07475_),
    .A(net2279),
    .B(net2362));
 sg13g2_xor2_1 _10575_ (.B(net2363),
    .A(net2280),
    .X(_07486_));
 sg13g2_xor2_1 _10576_ (.B(net2602),
    .A(net2517),
    .X(_07497_));
 sg13g2_nand3_1 _10577_ (.B(_07475_),
    .C(_07497_),
    .A(_07464_),
    .Y(_07508_));
 sg13g2_a21o_1 _10578_ (.A2(_07475_),
    .A1(_07464_),
    .B1(_07497_),
    .X(_07519_));
 sg13g2_nand2_1 _10579_ (.Y(_07530_),
    .A(_07508_),
    .B(_07519_));
 sg13g2_xnor2_1 _10580_ (.Y(_07541_),
    .A(_07442_),
    .B(_07530_));
 sg13g2_xnor2_1 _10581_ (.Y(_07552_),
    .A(net2216),
    .B(net2715));
 sg13g2_xor2_1 _10582_ (.B(net2349),
    .A(net2434),
    .X(_07563_));
 sg13g2_o21ai_1 _10583_ (.B1(_07563_),
    .Y(_07574_),
    .A1(net2734),
    .A2(net2682));
 sg13g2_nor2b_1 _10584_ (.A(net2287),
    .B_N(net2222),
    .Y(_07585_));
 sg13g2_xor2_1 _10585_ (.B(net2288),
    .A(net2222),
    .X(_07596_));
 sg13g2_nor2_1 _10586_ (.A(net2190),
    .B(net2743),
    .Y(_07607_));
 sg13g2_xnor2_1 _10587_ (.Y(_07618_),
    .A(_07596_),
    .B(_07607_));
 sg13g2_xnor2_1 _10588_ (.Y(_07629_),
    .A(_07574_),
    .B(_07618_));
 sg13g2_xnor2_1 _10589_ (.Y(_07640_),
    .A(_07552_),
    .B(_07629_));
 sg13g2_nand2_1 _10590_ (.Y(_07651_),
    .A(_07541_),
    .B(_07640_));
 sg13g2_nor2_1 _10591_ (.A(_07541_),
    .B(_07640_),
    .Y(_07662_));
 sg13g2_xor2_1 _10592_ (.B(_07640_),
    .A(_07541_),
    .X(_07673_));
 sg13g2_xnor2_1 _10593_ (.Y(_07684_),
    .A(net2694),
    .B(net2738));
 sg13g2_nand2b_1 _10594_ (.Y(_07695_),
    .B(net2757),
    .A_N(net2412));
 sg13g2_nor2_1 _10595_ (.A(net2596),
    .B(net2502),
    .Y(_07706_));
 sg13g2_xnor2_1 _10596_ (.Y(_07717_),
    .A(_07695_),
    .B(_07706_));
 sg13g2_nand2_1 _10597_ (.Y(_07728_),
    .A(_07684_),
    .B(_07717_));
 sg13g2_or2_1 _10598_ (.X(_07739_),
    .B(_07717_),
    .A(_07684_));
 sg13g2_nand2_1 _10599_ (.Y(_07750_),
    .A(_07728_),
    .B(_07739_));
 sg13g2_nor2_1 _10600_ (.A(net2786),
    .B(net2748),
    .Y(_07761_));
 sg13g2_xor2_1 _10601_ (.B(net2781),
    .A(net2707),
    .X(_07772_));
 sg13g2_xnor2_1 _10602_ (.Y(_07783_),
    .A(_07761_),
    .B(_07772_));
 sg13g2_xor2_1 _10603_ (.B(_07783_),
    .A(_07750_),
    .X(_07794_));
 sg13g2_xnor2_1 _10604_ (.Y(_07805_),
    .A(_07673_),
    .B(_07794_));
 sg13g2_nand2_1 _10605_ (.Y(_07816_),
    .A(_07420_),
    .B(_07805_));
 sg13g2_or2_1 _10606_ (.X(_07827_),
    .B(_07805_),
    .A(_07420_));
 sg13g2_nand2_1 _10607_ (.Y(_07838_),
    .A(_07816_),
    .B(_07827_));
 sg13g2_xnor2_1 _10608_ (.Y(_07849_),
    .A(net2430),
    .B(net2345));
 sg13g2_or3_2 _10609_ (.A(net2799),
    .B(net2309),
    .C(_07849_),
    .X(_07860_));
 sg13g2_xnor2_1 _10610_ (.Y(_07871_),
    .A(net2389),
    .B(net2220));
 sg13g2_nor2_1 _10611_ (.A(\net.in[253] ),
    .B(_07871_),
    .Y(_07882_));
 sg13g2_xor2_1 _10612_ (.B(net2638),
    .A(net2729),
    .X(_07893_));
 sg13g2_a21oi_2 _10613_ (.B1(_07893_),
    .Y(_07904_),
    .A2(_05418_),
    .A1(_05264_));
 sg13g2_nand2_1 _10614_ (.Y(_07915_),
    .A(_07882_),
    .B(_07904_));
 sg13g2_xnor2_1 _10615_ (.Y(_07926_),
    .A(_07882_),
    .B(_07904_));
 sg13g2_xnor2_1 _10616_ (.Y(_07937_),
    .A(_07860_),
    .B(_07926_));
 sg13g2_nor2_1 _10617_ (.A(net2722),
    .B(net2562),
    .Y(_07948_));
 sg13g2_xnor2_1 _10618_ (.Y(_07959_),
    .A(net2652),
    .B(_07948_));
 sg13g2_nor2_2 _10619_ (.A(net2686),
    .B(net2341),
    .Y(_07970_));
 sg13g2_xnor2_1 _10620_ (.Y(_07981_),
    .A(_07145_),
    .B(_07970_));
 sg13g2_a21o_1 _10621_ (.A2(net2370),
    .A1(net2460),
    .B1(_07981_),
    .X(_07992_));
 sg13g2_nand3_1 _10622_ (.B(net2370),
    .C(_07981_),
    .A(net2460),
    .Y(_08003_));
 sg13g2_nand2_1 _10623_ (.Y(_08014_),
    .A(_07992_),
    .B(_08003_));
 sg13g2_xnor2_1 _10624_ (.Y(_08025_),
    .A(_07959_),
    .B(_08014_));
 sg13g2_nand2_1 _10625_ (.Y(_08036_),
    .A(_07937_),
    .B(_08025_));
 sg13g2_or2_1 _10626_ (.X(_08047_),
    .B(_08025_),
    .A(_07937_));
 sg13g2_nand2_1 _10627_ (.Y(_08058_),
    .A(_08036_),
    .B(_08047_));
 sg13g2_xor2_1 _10628_ (.B(net2547),
    .A(net2757),
    .X(_08069_));
 sg13g2_xor2_1 _10629_ (.B(net2760),
    .A(net2393),
    .X(_08080_));
 sg13g2_nand2_1 _10630_ (.Y(_08091_),
    .A(_08069_),
    .B(_08080_));
 sg13g2_nor2b_1 _10631_ (.A(net2304),
    .B_N(net2249),
    .Y(_08102_));
 sg13g2_nor3_1 _10632_ (.A(net2357),
    .B(_05330_),
    .C(_08102_),
    .Y(_08113_));
 sg13g2_o21ai_1 _10633_ (.B1(_08113_),
    .Y(_08124_),
    .A1(_05066_),
    .A2(net2248));
 sg13g2_xor2_1 _10634_ (.B(_08124_),
    .A(_08091_),
    .X(_08135_));
 sg13g2_nor2_1 _10635_ (.A(net2264),
    .B(net2707),
    .Y(_08146_));
 sg13g2_nor2_1 _10636_ (.A(net2614),
    .B(net2725),
    .Y(_08157_));
 sg13g2_xnor2_1 _10637_ (.Y(_08168_),
    .A(_08146_),
    .B(_08157_));
 sg13g2_xnor2_1 _10638_ (.Y(_08179_),
    .A(_08135_),
    .B(_08168_));
 sg13g2_xor2_1 _10639_ (.B(_08179_),
    .A(_08058_),
    .X(_08190_));
 sg13g2_xor2_1 _10640_ (.B(_08190_),
    .A(_07838_),
    .X(_08201_));
 sg13g2_and2_1 _10641_ (.A(_06958_),
    .B(_08201_),
    .X(_08212_));
 sg13g2_xor2_1 _10642_ (.B(_08201_),
    .A(_06958_),
    .X(_08223_));
 sg13g2_nor2_1 _10643_ (.A(net2662),
    .B(net2642),
    .Y(_08234_));
 sg13g2_xnor2_1 _10644_ (.Y(_08245_),
    .A(net2732),
    .B(_08234_));
 sg13g2_xnor2_1 _10645_ (.Y(_08256_),
    .A(net2646),
    .B(net2320));
 sg13g2_nor2_2 _10646_ (.A(net2729),
    .B(net2762),
    .Y(_08267_));
 sg13g2_nor2_1 _10647_ (.A(net2699),
    .B(net2757),
    .Y(_08278_));
 sg13g2_xor2_1 _10648_ (.B(_08278_),
    .A(_08267_),
    .X(_08289_));
 sg13g2_nor2_1 _10649_ (.A(_08256_),
    .B(_08289_),
    .Y(_08300_));
 sg13g2_nand2_1 _10650_ (.Y(_08311_),
    .A(_08256_),
    .B(_08289_));
 sg13g2_nand2b_1 _10651_ (.Y(_08322_),
    .B(_08311_),
    .A_N(_08300_));
 sg13g2_xnor2_1 _10652_ (.Y(_08333_),
    .A(_08245_),
    .B(_08322_));
 sg13g2_xor2_1 _10653_ (.B(net2781),
    .A(net2311),
    .X(_08344_));
 sg13g2_nor2_2 _10654_ (.A(_06133_),
    .B(_08344_),
    .Y(_08355_));
 sg13g2_nor2b_1 _10655_ (.A(net2190),
    .B_N(net2252),
    .Y(_08366_));
 sg13g2_xor2_1 _10656_ (.B(net2251),
    .A(net2191),
    .X(_08377_));
 sg13g2_nor2_1 _10657_ (.A(net2729),
    .B(net2200),
    .Y(_08388_));
 sg13g2_nor2_1 _10658_ (.A(_08377_),
    .B(_08388_),
    .Y(_08399_));
 sg13g2_nor2_1 _10659_ (.A(net2342),
    .B(net2395),
    .Y(_08410_));
 sg13g2_xor2_1 _10660_ (.B(net2395),
    .A(net2343),
    .X(_08421_));
 sg13g2_nand2b_1 _10661_ (.Y(_08432_),
    .B(net2492),
    .A_N(net2704));
 sg13g2_xnor2_1 _10662_ (.Y(_08443_),
    .A(_08421_),
    .B(_08432_));
 sg13g2_nor3_1 _10663_ (.A(_08377_),
    .B(_08388_),
    .C(_08443_),
    .Y(_08454_));
 sg13g2_nand2b_1 _10664_ (.Y(_08465_),
    .B(_08443_),
    .A_N(_08399_));
 sg13g2_xnor2_1 _10665_ (.Y(_08476_),
    .A(_08399_),
    .B(_08443_));
 sg13g2_xnor2_1 _10666_ (.Y(_08487_),
    .A(_08355_),
    .B(_08476_));
 sg13g2_nor2_1 _10667_ (.A(net2448),
    .B(net2291),
    .Y(_08498_));
 sg13g2_xnor2_1 _10668_ (.Y(_08509_),
    .A(net2750),
    .B(net2311));
 sg13g2_xor2_1 _10669_ (.B(_08509_),
    .A(_08498_),
    .X(_08520_));
 sg13g2_xnor2_1 _10670_ (.Y(_08531_),
    .A(net2711),
    .B(net2732));
 sg13g2_nor2b_1 _10671_ (.A(net2707),
    .B_N(net2762),
    .Y(_08542_));
 sg13g2_xnor2_1 _10672_ (.Y(_08553_),
    .A(net2694),
    .B(net2320));
 sg13g2_xnor2_1 _10673_ (.Y(_08564_),
    .A(_08542_),
    .B(_08553_));
 sg13g2_nor2_1 _10674_ (.A(_08531_),
    .B(_08564_),
    .Y(_08575_));
 sg13g2_xnor2_1 _10675_ (.Y(_08586_),
    .A(_08531_),
    .B(_08564_));
 sg13g2_a21oi_1 _10676_ (.A1(_08531_),
    .A2(_08564_),
    .Y(_08597_),
    .B1(_08520_));
 sg13g2_nor2_2 _10677_ (.A(_08575_),
    .B(_08597_),
    .Y(_08608_));
 sg13g2_xnor2_1 _10678_ (.Y(_08619_),
    .A(_08520_),
    .B(_08586_));
 sg13g2_nor2_1 _10679_ (.A(_08487_),
    .B(_08619_),
    .Y(_08630_));
 sg13g2_nand2_1 _10680_ (.Y(_08641_),
    .A(_08487_),
    .B(_08619_));
 sg13g2_a21oi_1 _10681_ (.A1(_08333_),
    .A2(_08641_),
    .Y(_08652_),
    .B1(_08630_));
 sg13g2_nand2b_1 _10682_ (.Y(_08663_),
    .B(_08641_),
    .A_N(_08630_));
 sg13g2_xnor2_1 _10683_ (.Y(_08674_),
    .A(_08333_),
    .B(_08663_));
 sg13g2_xor2_1 _10684_ (.B(net2700),
    .A(net2389),
    .X(_08685_));
 sg13g2_xnor2_1 _10685_ (.Y(_08696_),
    .A(net2304),
    .B(net2405));
 sg13g2_nand2_2 _10686_ (.Y(_08707_),
    .A(_08685_),
    .B(_08696_));
 sg13g2_xnor2_1 _10687_ (.Y(_08718_),
    .A(net2471),
    .B(net2322));
 sg13g2_nor3_2 _10688_ (.A(net2354),
    .B(net2316),
    .C(_08718_),
    .Y(_08729_));
 sg13g2_nor2_1 _10689_ (.A(net2591),
    .B(net2548),
    .Y(_08740_));
 sg13g2_nand2_1 _10690_ (.Y(_08751_),
    .A(net2539),
    .B(net2729));
 sg13g2_xor2_1 _10691_ (.B(_08751_),
    .A(_08740_),
    .X(_08762_));
 sg13g2_nand2_1 _10692_ (.Y(_08773_),
    .A(_08729_),
    .B(_08762_));
 sg13g2_nor2_1 _10693_ (.A(_08729_),
    .B(_08762_),
    .Y(_08784_));
 sg13g2_xor2_1 _10694_ (.B(_08762_),
    .A(_08729_),
    .X(_08795_));
 sg13g2_xnor2_1 _10695_ (.Y(_08806_),
    .A(_08707_),
    .B(_08795_));
 sg13g2_nor2_1 _10696_ (.A(net2405),
    .B(net2707),
    .Y(_08817_));
 sg13g2_o21ai_1 _10697_ (.B1(_08817_),
    .Y(_08828_),
    .A1(net2506),
    .A2(net2575));
 sg13g2_xor2_1 _10698_ (.B(net2310),
    .A(net2222),
    .X(_08839_));
 sg13g2_or3_2 _10699_ (.A(net2357),
    .B(net2773),
    .C(_08839_),
    .X(_08850_));
 sg13g2_inv_1 _10700_ (.Y(_08861_),
    .A(_08850_));
 sg13g2_xnor2_1 _10701_ (.Y(_08872_),
    .A(net2764),
    .B(net2349));
 sg13g2_xnor2_1 _10702_ (.Y(_08883_),
    .A(_06969_),
    .B(_08872_));
 sg13g2_nand2_1 _10703_ (.Y(_08894_),
    .A(_08861_),
    .B(_08883_));
 sg13g2_xnor2_1 _10704_ (.Y(_08905_),
    .A(_08850_),
    .B(_08883_));
 sg13g2_xnor2_1 _10705_ (.Y(_08916_),
    .A(_08828_),
    .B(_08905_));
 sg13g2_nand2_1 _10706_ (.Y(_08927_),
    .A(_08806_),
    .B(_08916_));
 sg13g2_nor2_1 _10707_ (.A(_08806_),
    .B(_08916_),
    .Y(_08938_));
 sg13g2_xnor2_1 _10708_ (.Y(_08949_),
    .A(_08806_),
    .B(_08916_));
 sg13g2_nor2_1 _10709_ (.A(net2772),
    .B(net2361),
    .Y(_08960_));
 sg13g2_o21ai_1 _10710_ (.B1(_08960_),
    .Y(_08971_),
    .A1(net2453),
    .A2(net2442));
 sg13g2_a21oi_2 _10711_ (.B1(_08971_),
    .Y(_08982_),
    .A2(net2442),
    .A1(net2454));
 sg13g2_a22oi_1 _10712_ (.Y(_08993_),
    .B1(net2203),
    .B2(\net.in[252] ),
    .A2(net2722),
    .A1(_05077_));
 sg13g2_o21ai_1 _10713_ (.B1(_08993_),
    .Y(_09004_),
    .A1(net2203),
    .A2(\net.in[252] ));
 sg13g2_nor2_1 _10714_ (.A(net2179),
    .B(net2407),
    .Y(_09015_));
 sg13g2_o21ai_1 _10715_ (.B1(_09004_),
    .Y(_09026_),
    .A1(net2179),
    .A2(net2407));
 sg13g2_nor2b_1 _10716_ (.A(_09004_),
    .B_N(_09015_),
    .Y(_09037_));
 sg13g2_xnor2_1 _10717_ (.Y(_09048_),
    .A(_09004_),
    .B(_09015_));
 sg13g2_a21oi_2 _10718_ (.B1(_09037_),
    .Y(_09059_),
    .A2(_09026_),
    .A1(_08982_));
 sg13g2_xnor2_1 _10719_ (.Y(_09070_),
    .A(_08982_),
    .B(_09048_));
 sg13g2_or2_1 _10720_ (.X(_09081_),
    .B(_09070_),
    .A(_08938_));
 sg13g2_xnor2_1 _10721_ (.Y(_09092_),
    .A(_08949_),
    .B(_09070_));
 sg13g2_nor2_1 _10722_ (.A(net2448),
    .B(net2311),
    .Y(_09103_));
 sg13g2_o21ai_1 _10723_ (.B1(_09103_),
    .Y(_09114_),
    .A1(net2376),
    .A2(net2602));
 sg13g2_nor2b_1 _10724_ (.A(net2448),
    .B_N(net2463),
    .Y(_09125_));
 sg13g2_xnor2_1 _10725_ (.Y(_09136_),
    .A(net2752),
    .B(net2291));
 sg13g2_xnor2_1 _10726_ (.Y(_09147_),
    .A(_09125_),
    .B(_09136_));
 sg13g2_xnor2_1 _10727_ (.Y(_09158_),
    .A(net2716),
    .B(net2629));
 sg13g2_nor2_1 _10728_ (.A(net2312),
    .B(net2246),
    .Y(_09169_));
 sg13g2_xnor2_1 _10729_ (.Y(_09180_),
    .A(_09158_),
    .B(_09169_));
 sg13g2_inv_1 _10730_ (.Y(_09191_),
    .A(_09180_));
 sg13g2_nand2_1 _10731_ (.Y(_09202_),
    .A(_09147_),
    .B(_09191_));
 sg13g2_nor2_1 _10732_ (.A(_09147_),
    .B(_09191_),
    .Y(_09213_));
 sg13g2_xnor2_1 _10733_ (.Y(_09224_),
    .A(_09147_),
    .B(_09180_));
 sg13g2_xnor2_1 _10734_ (.Y(_09235_),
    .A(_09114_),
    .B(_09224_));
 sg13g2_nor2_2 _10735_ (.A(net2259),
    .B(_05803_),
    .Y(_09246_));
 sg13g2_xor2_1 _10736_ (.B(net2328),
    .A(net2259),
    .X(_09257_));
 sg13g2_and3_2 _10737_ (.X(_09268_),
    .A(_05275_),
    .B(net2722),
    .C(_09257_));
 sg13g2_nor2_1 _10738_ (.A(net2792),
    .B(net2710),
    .Y(_09279_));
 sg13g2_nor2_1 _10739_ (.A(net2614),
    .B(\net.in[238] ),
    .Y(_09290_));
 sg13g2_xor2_1 _10740_ (.B(_09290_),
    .A(_09279_),
    .X(_09301_));
 sg13g2_nand2_1 _10741_ (.Y(_09312_),
    .A(_09268_),
    .B(_09301_));
 sg13g2_xnor2_1 _10742_ (.Y(_09323_),
    .A(_09268_),
    .B(_09301_));
 sg13g2_xor2_1 _10743_ (.B(net2757),
    .A(net2492),
    .X(_09334_));
 sg13g2_xnor2_1 _10744_ (.Y(_09345_),
    .A(_09323_),
    .B(_09334_));
 sg13g2_nor2_1 _10745_ (.A(_09235_),
    .B(_09345_),
    .Y(_09356_));
 sg13g2_nand2_1 _10746_ (.Y(_09367_),
    .A(_09235_),
    .B(_09345_));
 sg13g2_xor2_1 _10747_ (.B(_09345_),
    .A(_09235_),
    .X(_09378_));
 sg13g2_xnor2_1 _10748_ (.Y(_09389_),
    .A(net2566),
    .B(net2501));
 sg13g2_nor2_1 _10749_ (.A(net2660),
    .B(_09389_),
    .Y(_09400_));
 sg13g2_nor2_1 _10750_ (.A(net2603),
    .B(net2596),
    .Y(_09411_));
 sg13g2_nor3_2 _10751_ (.A(net2332),
    .B(net2316),
    .C(_09411_),
    .Y(_09422_));
 sg13g2_nor2_2 _10752_ (.A(net2639),
    .B(net2700),
    .Y(_09433_));
 sg13g2_nor2_1 _10753_ (.A(net2311),
    .B(net2651),
    .Y(_09444_));
 sg13g2_xnor2_1 _10754_ (.Y(_09455_),
    .A(_09433_),
    .B(_09444_));
 sg13g2_nand2b_1 _10755_ (.Y(_09466_),
    .B(_09422_),
    .A_N(_09455_));
 sg13g2_nand2b_1 _10756_ (.Y(_09477_),
    .B(_09455_),
    .A_N(_09422_));
 sg13g2_nand2_1 _10757_ (.Y(_09488_),
    .A(_09466_),
    .B(_09477_));
 sg13g2_xor2_1 _10758_ (.B(_09488_),
    .A(_09400_),
    .X(_09499_));
 sg13g2_xnor2_1 _10759_ (.Y(_09510_),
    .A(_09378_),
    .B(_09499_));
 sg13g2_inv_1 _10760_ (.Y(_09521_),
    .A(_09510_));
 sg13g2_nor2_1 _10761_ (.A(_09092_),
    .B(_09521_),
    .Y(_09532_));
 sg13g2_nor2_1 _10762_ (.A(_08674_),
    .B(_09532_),
    .Y(_09543_));
 sg13g2_a21oi_2 _10763_ (.B1(_09543_),
    .Y(_09554_),
    .A2(_09521_),
    .A1(_09092_));
 sg13g2_xnor2_1 _10764_ (.Y(_09565_),
    .A(_09092_),
    .B(_09510_));
 sg13g2_xnor2_1 _10765_ (.Y(_09576_),
    .A(_08674_),
    .B(_09565_));
 sg13g2_xor2_1 _10766_ (.B(net2743),
    .A(net2606),
    .X(_09587_));
 sg13g2_xor2_1 _10767_ (.B(net2194),
    .A(net2231),
    .X(_09598_));
 sg13g2_xnor2_1 _10768_ (.Y(_09609_),
    .A(_09587_),
    .B(_09598_));
 sg13g2_or2_1 _10769_ (.X(_09620_),
    .B(_09609_),
    .A(_06705_));
 sg13g2_xor2_1 _10770_ (.B(_09609_),
    .A(_06705_),
    .X(_09631_));
 sg13g2_xor2_1 _10771_ (.B(net2364),
    .A(net2586),
    .X(_09642_));
 sg13g2_xnor2_1 _10772_ (.Y(_09653_),
    .A(_09631_),
    .B(_09642_));
 sg13g2_o21ai_1 _10773_ (.B1(_00000_),
    .Y(_09664_),
    .A1(net2567),
    .A2(net2458));
 sg13g2_a21oi_1 _10774_ (.A1(net2566),
    .A2(net2458),
    .Y(_09675_),
    .B1(_09664_));
 sg13g2_xnor2_1 _10775_ (.Y(_09686_),
    .A(net2510),
    .B(net2410));
 sg13g2_inv_4 _10776_ (.A(_09686_),
    .Y(_09697_));
 sg13g2_nor2_1 _10777_ (.A(net2305),
    .B(_05110_),
    .Y(_09708_));
 sg13g2_nor2_2 _10778_ (.A(_05066_),
    .B(net2241),
    .Y(_09719_));
 sg13g2_nor3_2 _10779_ (.A(_06254_),
    .B(_09708_),
    .C(_09719_),
    .Y(_09730_));
 sg13g2_nor2_1 _10780_ (.A(_09697_),
    .B(_09730_),
    .Y(_09741_));
 sg13g2_xnor2_1 _10781_ (.Y(_09752_),
    .A(_09686_),
    .B(_09730_));
 sg13g2_xnor2_1 _10782_ (.Y(_09763_),
    .A(_09675_),
    .B(_09752_));
 sg13g2_nand2_1 _10783_ (.Y(_09774_),
    .A(_09653_),
    .B(_09763_));
 sg13g2_nor2_1 _10784_ (.A(_09653_),
    .B(_09763_),
    .Y(_09785_));
 sg13g2_xor2_1 _10785_ (.B(_09763_),
    .A(_09653_),
    .X(_09796_));
 sg13g2_nor2_1 _10786_ (.A(_05022_),
    .B(net2534),
    .Y(_09807_));
 sg13g2_nor2b_1 _10787_ (.A(net2430),
    .B_N(net2534),
    .Y(_09818_));
 sg13g2_xor2_1 _10788_ (.B(net2605),
    .A(net2705),
    .X(_09829_));
 sg13g2_nor3_2 _10789_ (.A(_09807_),
    .B(_09818_),
    .C(_09829_),
    .Y(_09840_));
 sg13g2_nand2_1 _10790_ (.Y(_09850_),
    .A(_05209_),
    .B(net2592));
 sg13g2_nor2_1 _10791_ (.A(_05209_),
    .B(net2592),
    .Y(_09855_));
 sg13g2_nor3_1 _10792_ (.A(net2548),
    .B(\net.in[238] ),
    .C(_09855_),
    .Y(_00279_));
 sg13g2_xnor2_1 _10793_ (.Y(_00285_),
    .A(net2752),
    .B(net2675));
 sg13g2_a21oi_1 _10794_ (.A1(_09850_),
    .A2(_00279_),
    .Y(_00287_),
    .B1(_00285_));
 sg13g2_nand3_1 _10795_ (.B(_00279_),
    .C(_00285_),
    .A(_09850_),
    .Y(_00290_));
 sg13g2_nand2b_1 _10796_ (.Y(_00294_),
    .B(_00290_),
    .A_N(_00287_));
 sg13g2_xnor2_1 _10797_ (.Y(_00297_),
    .A(_09840_),
    .B(_00294_));
 sg13g2_xnor2_1 _10798_ (.Y(_00301_),
    .A(_09796_),
    .B(_00297_));
 sg13g2_xor2_1 _10799_ (.B(net2488),
    .A(net2530),
    .X(_00305_));
 sg13g2_nor2_1 _10800_ (.A(net2403),
    .B(net2393),
    .Y(_00310_));
 sg13g2_nor2_1 _10801_ (.A(net2521),
    .B(net2473),
    .Y(_00314_));
 sg13g2_xnor2_1 _10802_ (.Y(_00320_),
    .A(_00310_),
    .B(_00314_));
 sg13g2_nand2b_1 _10803_ (.Y(_00324_),
    .B(net2740),
    .A_N(net2729));
 sg13g2_xnor2_1 _10804_ (.Y(_00329_),
    .A(net2530),
    .B(net2458));
 sg13g2_xnor2_1 _10805_ (.Y(_00333_),
    .A(_00324_),
    .B(_00329_));
 sg13g2_nand2_1 _10806_ (.Y(_00338_),
    .A(_00320_),
    .B(_00333_));
 sg13g2_xor2_1 _10807_ (.B(_00333_),
    .A(_00320_),
    .X(_00344_));
 sg13g2_xnor2_1 _10808_ (.Y(_00348_),
    .A(_00305_),
    .B(_00344_));
 sg13g2_xnor2_1 _10809_ (.Y(_00353_),
    .A(net2646),
    .B(net2725));
 sg13g2_nand2_2 _10810_ (.Y(_00358_),
    .A(_07563_),
    .B(_00353_));
 sg13g2_nor2_1 _10811_ (.A(net2799),
    .B(net2279),
    .Y(_00364_));
 sg13g2_xnor2_1 _10812_ (.Y(_00369_),
    .A(net2416),
    .B(net2295));
 sg13g2_xnor2_1 _10813_ (.Y(_00374_),
    .A(_00364_),
    .B(_00369_));
 sg13g2_nor2_1 _10814_ (.A(_00358_),
    .B(_00374_),
    .Y(_00378_));
 sg13g2_nand2_1 _10815_ (.Y(_00384_),
    .A(_00358_),
    .B(_00374_));
 sg13g2_xor2_1 _10816_ (.B(_00374_),
    .A(_00358_),
    .X(_00389_));
 sg13g2_xnor2_1 _10817_ (.Y(_00395_),
    .A(net2307),
    .B(_00014_));
 sg13g2_xnor2_1 _10818_ (.Y(_00400_),
    .A(net2449),
    .B(_00395_));
 sg13g2_xnor2_1 _10819_ (.Y(_00405_),
    .A(_00389_),
    .B(_00400_));
 sg13g2_nand2_1 _10820_ (.Y(_00411_),
    .A(_00348_),
    .B(_00405_));
 sg13g2_xnor2_1 _10821_ (.Y(_00416_),
    .A(_00348_),
    .B(_00405_));
 sg13g2_nor2_2 _10822_ (.A(net2256),
    .B(net2230),
    .Y(_00421_));
 sg13g2_nor3_2 _10823_ (.A(net2256),
    .B(net2230),
    .C(_00015_),
    .Y(_00425_));
 sg13g2_nor2_1 _10824_ (.A(net2547),
    .B(net2548),
    .Y(_00430_));
 sg13g2_xnor2_1 _10825_ (.Y(_00435_),
    .A(net2388),
    .B(net2393));
 sg13g2_inv_2 _10826_ (.Y(_00439_),
    .A(_00435_));
 sg13g2_nor2_2 _10827_ (.A(net2381),
    .B(_00435_),
    .Y(_00443_));
 sg13g2_nor2_1 _10828_ (.A(_05363_),
    .B(net2393),
    .Y(_00447_));
 sg13g2_or3_1 _10829_ (.A(_00430_),
    .B(_00443_),
    .C(_00447_),
    .X(_00450_));
 sg13g2_o21ai_1 _10830_ (.B1(_00430_),
    .Y(_00454_),
    .A1(_00443_),
    .A2(_00447_));
 sg13g2_nand2_1 _10831_ (.Y(_00459_),
    .A(_00450_),
    .B(_00454_));
 sg13g2_xor2_1 _10832_ (.B(_00459_),
    .A(_00425_),
    .X(_00464_));
 sg13g2_xnor2_1 _10833_ (.Y(_00470_),
    .A(_00416_),
    .B(_00464_));
 sg13g2_nand2b_2 _10834_ (.Y(_00472_),
    .B(net2671),
    .A_N(net2560));
 sg13g2_xnor2_1 _10835_ (.Y(_00473_),
    .A(net2669),
    .B(net2606));
 sg13g2_nand2_1 _10836_ (.Y(_00474_),
    .A(net2559),
    .B(_00473_));
 sg13g2_nand2_2 _10837_ (.Y(_00475_),
    .A(_00472_),
    .B(_00474_));
 sg13g2_nand2_1 _10838_ (.Y(_00476_),
    .A(net2227),
    .B(net2363));
 sg13g2_nor2_2 _10839_ (.A(net2226),
    .B(net2362),
    .Y(_00477_));
 sg13g2_o21ai_1 _10840_ (.B1(_00476_),
    .Y(_00478_),
    .A1(_05143_),
    .A2(net2379));
 sg13g2_o21ai_1 _10841_ (.B1(_00430_),
    .Y(_00479_),
    .A1(net2177),
    .A2(net2407));
 sg13g2_o21ai_1 _10842_ (.B1(_00479_),
    .Y(_00480_),
    .A1(_00477_),
    .A2(_00478_));
 sg13g2_or3_1 _10843_ (.A(_00477_),
    .B(_00478_),
    .C(_00479_),
    .X(_00481_));
 sg13g2_nand2_1 _10844_ (.Y(_00482_),
    .A(_00480_),
    .B(_00481_));
 sg13g2_xor2_1 _10845_ (.B(_00482_),
    .A(_00475_),
    .X(_00483_));
 sg13g2_xor2_1 _10846_ (.B(net2547),
    .A(net2769),
    .X(_00484_));
 sg13g2_nand2b_1 _10847_ (.Y(_00485_),
    .B(net2788),
    .A_N(net2724));
 sg13g2_nor2_1 _10848_ (.A(net2789),
    .B(net2720),
    .Y(_00486_));
 sg13g2_xnor2_1 _10849_ (.Y(_00487_),
    .A(net2787),
    .B(net2722));
 sg13g2_xnor2_1 _10850_ (.Y(_00488_),
    .A(_00484_),
    .B(_00487_));
 sg13g2_nand2_1 _10851_ (.Y(_00489_),
    .A(net2216),
    .B(net2734));
 sg13g2_nor2_1 _10852_ (.A(net2368),
    .B(net2285),
    .Y(_00490_));
 sg13g2_xor2_1 _10853_ (.B(_00490_),
    .A(_00489_),
    .X(_00491_));
 sg13g2_inv_1 _10854_ (.Y(_00492_),
    .A(_00491_));
 sg13g2_nor2_1 _10855_ (.A(_00488_),
    .B(_00492_),
    .Y(_00493_));
 sg13g2_xnor2_1 _10856_ (.Y(_00494_),
    .A(_00488_),
    .B(_00491_));
 sg13g2_xor2_1 _10857_ (.B(net2790),
    .A(net2689),
    .X(_00495_));
 sg13g2_nor2_1 _10858_ (.A(net2553),
    .B(net2264),
    .Y(_00496_));
 sg13g2_xnor2_1 _10859_ (.Y(_00497_),
    .A(_00495_),
    .B(_00496_));
 sg13g2_xnor2_1 _10860_ (.Y(_00498_),
    .A(_00494_),
    .B(_00497_));
 sg13g2_nand2b_1 _10861_ (.Y(_00499_),
    .B(net2575),
    .A_N(net2481));
 sg13g2_xnor2_1 _10862_ (.Y(_00500_),
    .A(net2492),
    .B(net2535));
 sg13g2_xnor2_1 _10863_ (.Y(_00501_),
    .A(_00499_),
    .B(_00500_));
 sg13g2_nand2b_1 _10864_ (.Y(_00502_),
    .B(net2571),
    .A_N(net2453));
 sg13g2_xnor2_1 _10865_ (.Y(_00503_),
    .A(net2562),
    .B(net2606));
 sg13g2_xnor2_1 _10866_ (.Y(_00504_),
    .A(_00502_),
    .B(_00503_));
 sg13g2_inv_1 _10867_ (.Y(_00505_),
    .A(_00504_));
 sg13g2_nand2_1 _10868_ (.Y(_00506_),
    .A(_00501_),
    .B(_00505_));
 sg13g2_nor2_1 _10869_ (.A(_00501_),
    .B(_00505_),
    .Y(_00507_));
 sg13g2_xor2_1 _10870_ (.B(_00504_),
    .A(_00501_),
    .X(_00508_));
 sg13g2_nor2_2 _10871_ (.A(net2449),
    .B(net2745),
    .Y(_00509_));
 sg13g2_nor2_1 _10872_ (.A(net2509),
    .B(net2457),
    .Y(_00510_));
 sg13g2_xor2_1 _10873_ (.B(_00510_),
    .A(_00509_),
    .X(_00511_));
 sg13g2_a21oi_2 _10874_ (.B1(_00507_),
    .Y(_00512_),
    .A2(_00511_),
    .A1(_00506_));
 sg13g2_xnor2_1 _10875_ (.Y(_00513_),
    .A(_00508_),
    .B(_00511_));
 sg13g2_nand2b_1 _10876_ (.Y(_00514_),
    .B(_00513_),
    .A_N(_00498_));
 sg13g2_nor2b_1 _10877_ (.A(_00513_),
    .B_N(_00498_),
    .Y(_00515_));
 sg13g2_xnor2_1 _10878_ (.Y(_00516_),
    .A(_00498_),
    .B(_00513_));
 sg13g2_o21ai_1 _10879_ (.B1(_00514_),
    .Y(_00517_),
    .A1(_00483_),
    .A2(_00515_));
 sg13g2_xnor2_1 _10880_ (.Y(_00518_),
    .A(_00483_),
    .B(_00516_));
 sg13g2_nand2b_1 _10881_ (.Y(_00519_),
    .B(_00518_),
    .A_N(_00470_));
 sg13g2_nand2b_1 _10882_ (.Y(_00520_),
    .B(_00470_),
    .A_N(_00518_));
 sg13g2_xor2_1 _10883_ (.B(_00518_),
    .A(_00470_),
    .X(_00521_));
 sg13g2_xnor2_1 _10884_ (.Y(_00522_),
    .A(_00301_),
    .B(_00521_));
 sg13g2_nand2_1 _10885_ (.Y(_00523_),
    .A(_09576_),
    .B(_00522_));
 sg13g2_xor2_1 _10886_ (.B(_00522_),
    .A(_09576_),
    .X(_00524_));
 sg13g2_nor2_1 _10887_ (.A(net2237),
    .B(net2766),
    .Y(_00525_));
 sg13g2_xnor2_1 _10888_ (.Y(_00526_),
    .A(net2299),
    .B(net2740));
 sg13g2_xnor2_1 _10889_ (.Y(_00527_),
    .A(_00525_),
    .B(_00526_));
 sg13g2_and2_1 _10890_ (.A(net2603),
    .B(net2596),
    .X(_00528_));
 sg13g2_nor4_2 _10891_ (.A(net2235),
    .B(net2279),
    .C(_09411_),
    .Y(_00529_),
    .D(_00528_));
 sg13g2_o21ai_1 _10892_ (.B1(net2517),
    .Y(_00530_),
    .A1(net2677),
    .A2(net2652));
 sg13g2_inv_1 _10893_ (.Y(_00531_),
    .A(_00530_));
 sg13g2_xnor2_1 _10894_ (.Y(_00532_),
    .A(_00529_),
    .B(_00531_));
 sg13g2_a21o_1 _10895_ (.A2(_00531_),
    .A1(_00529_),
    .B1(_00527_),
    .X(_00533_));
 sg13g2_o21ai_1 _10896_ (.B1(_00533_),
    .Y(_00534_),
    .A1(_00529_),
    .A2(_00531_));
 sg13g2_xnor2_1 _10897_ (.Y(_00535_),
    .A(_00527_),
    .B(_00532_));
 sg13g2_xor2_1 _10898_ (.B(net2717),
    .A(net2218),
    .X(_00536_));
 sg13g2_xnor2_1 _10899_ (.Y(_00537_),
    .A(net2311),
    .B(net2248));
 sg13g2_nand2_1 _10900_ (.Y(_00538_),
    .A(_00536_),
    .B(_00537_));
 sg13g2_nor2b_1 _10901_ (.A(net2453),
    .B_N(net2418),
    .Y(_00539_));
 sg13g2_nor2_1 _10902_ (.A(net2364),
    .B(net2282),
    .Y(_00540_));
 sg13g2_xnor2_1 _10903_ (.Y(_00541_),
    .A(_00539_),
    .B(_00540_));
 sg13g2_nor2_1 _10904_ (.A(net2769),
    .B(net2364),
    .Y(_00542_));
 sg13g2_xor2_1 _10905_ (.B(net2416),
    .A(net2453),
    .X(_00543_));
 sg13g2_xnor2_1 _10906_ (.Y(_00544_),
    .A(_00542_),
    .B(_00543_));
 sg13g2_nand2_1 _10907_ (.Y(_00545_),
    .A(_00541_),
    .B(_00544_));
 sg13g2_nor2_1 _10908_ (.A(_00541_),
    .B(_00544_),
    .Y(_00546_));
 sg13g2_xor2_1 _10909_ (.B(_00544_),
    .A(_00541_),
    .X(_00547_));
 sg13g2_xnor2_1 _10910_ (.Y(_00548_),
    .A(_00538_),
    .B(_00547_));
 sg13g2_nand2_1 _10911_ (.Y(_00549_),
    .A(_00535_),
    .B(_00548_));
 sg13g2_or2_1 _10912_ (.X(_00550_),
    .B(_00548_),
    .A(_00535_));
 sg13g2_nand2_1 _10913_ (.Y(_00551_),
    .A(_00549_),
    .B(_00550_));
 sg13g2_nor2_1 _10914_ (.A(net2255),
    .B(net2199),
    .Y(_00552_));
 sg13g2_nor2_1 _10915_ (.A(net2517),
    .B(net2389),
    .Y(_00553_));
 sg13g2_xnor2_1 _10916_ (.Y(_00554_),
    .A(net2558),
    .B(_00553_));
 sg13g2_nor2_1 _10917_ (.A(net2786),
    .B(net2738),
    .Y(_00555_));
 sg13g2_nand2_1 _10918_ (.Y(_00556_),
    .A(net2716),
    .B(_05946_));
 sg13g2_xnor2_1 _10919_ (.Y(_00557_),
    .A(net2717),
    .B(_00555_));
 sg13g2_nor2b_1 _10920_ (.A(_00554_),
    .B_N(_00557_),
    .Y(_00558_));
 sg13g2_nand2b_1 _10921_ (.Y(_00559_),
    .B(_00554_),
    .A_N(_00557_));
 sg13g2_nor2b_1 _10922_ (.A(_00558_),
    .B_N(_00559_),
    .Y(_00560_));
 sg13g2_xnor2_1 _10923_ (.Y(_00561_),
    .A(_00552_),
    .B(_00560_));
 sg13g2_xor2_1 _10924_ (.B(_00561_),
    .A(_00551_),
    .X(_00562_));
 sg13g2_nand2b_2 _10925_ (.Y(_00563_),
    .B(net2556),
    .A_N(net2747));
 sg13g2_nor3_2 _10926_ (.A(net2405),
    .B(net2190),
    .C(_00563_),
    .Y(_00564_));
 sg13g2_xor2_1 _10927_ (.B(net2738),
    .A(net2786),
    .X(_00565_));
 sg13g2_nor2_1 _10928_ (.A(net2764),
    .B(net2787),
    .Y(_00566_));
 sg13g2_xnor2_1 _10929_ (.Y(_00567_),
    .A(_00565_),
    .B(_00566_));
 sg13g2_nor2b_1 _10930_ (.A(_00567_),
    .B_N(_00564_),
    .Y(_00568_));
 sg13g2_nand2b_1 _10931_ (.Y(_00569_),
    .B(_00567_),
    .A_N(_00564_));
 sg13g2_nor2b_1 _10932_ (.A(_00568_),
    .B_N(_00569_),
    .Y(_00570_));
 sg13g2_xnor2_1 _10933_ (.Y(_00571_),
    .A(net2442),
    .B(net2570));
 sg13g2_xnor2_1 _10934_ (.Y(_00572_),
    .A(_08267_),
    .B(_00571_));
 sg13g2_xor2_1 _10935_ (.B(_00572_),
    .A(_00570_),
    .X(_00573_));
 sg13g2_nor2_1 _10936_ (.A(net2684),
    .B(net2761),
    .Y(_00574_));
 sg13g2_xor2_1 _10937_ (.B(net2760),
    .A(net2682),
    .X(_00575_));
 sg13g2_o21ai_1 _10938_ (.B1(_00016_),
    .Y(_00576_),
    .A1(net2762),
    .A2(_05946_));
 sg13g2_nor2b_2 _10939_ (.A(net2755),
    .B_N(net2687),
    .Y(_00577_));
 sg13g2_xnor2_1 _10940_ (.Y(_00578_),
    .A(net2760),
    .B(_00577_));
 sg13g2_nand2_1 _10941_ (.Y(_00579_),
    .A(_00576_),
    .B(_00578_));
 sg13g2_nor2_1 _10942_ (.A(_00576_),
    .B(_00578_),
    .Y(_00580_));
 sg13g2_xnor2_1 _10943_ (.Y(_00581_),
    .A(_00576_),
    .B(_00578_));
 sg13g2_xnor2_1 _10944_ (.Y(_00582_),
    .A(_00575_),
    .B(_00581_));
 sg13g2_xnor2_1 _10945_ (.Y(_00583_),
    .A(net2642),
    .B(net2407));
 sg13g2_xnor2_1 _10946_ (.Y(_00584_),
    .A(net2662),
    .B(net2722));
 sg13g2_nor2_1 _10947_ (.A(_00583_),
    .B(_00584_),
    .Y(_00585_));
 sg13g2_nor2b_1 _10948_ (.A(net2207),
    .B_N(net2388),
    .Y(_00586_));
 sg13g2_or2_1 _10949_ (.X(_00587_),
    .B(net2499),
    .A(net2295));
 sg13g2_nand2b_1 _10950_ (.Y(_00588_),
    .B(net2513),
    .A_N(net2407));
 sg13g2_nand2b_1 _10951_ (.Y(_00589_),
    .B(net2501),
    .A_N(net2437));
 sg13g2_a22oi_1 _10952_ (.Y(_00590_),
    .B1(_00588_),
    .B2(_00589_),
    .A2(_00587_),
    .A1(_00586_));
 sg13g2_nand4_1 _10953_ (.B(_00587_),
    .C(_00588_),
    .A(_00586_),
    .Y(_00591_),
    .D(_00589_));
 sg13g2_nand2b_1 _10954_ (.Y(_00592_),
    .B(_00591_),
    .A_N(_00590_));
 sg13g2_xnor2_1 _10955_ (.Y(_00593_),
    .A(_00585_),
    .B(_00592_));
 sg13g2_nand2_1 _10956_ (.Y(_00594_),
    .A(_00582_),
    .B(_00593_));
 sg13g2_o21ai_1 _10957_ (.B1(_00573_),
    .Y(_00595_),
    .A1(_00582_),
    .A2(_00593_));
 sg13g2_nand2_1 _10958_ (.Y(_00596_),
    .A(_00594_),
    .B(_00595_));
 sg13g2_xor2_1 _10959_ (.B(_00593_),
    .A(_00582_),
    .X(_00597_));
 sg13g2_xnor2_1 _10960_ (.Y(_00598_),
    .A(_00573_),
    .B(_00597_));
 sg13g2_or2_1 _10961_ (.X(_00599_),
    .B(net2570),
    .A(net2460));
 sg13g2_o21ai_1 _10962_ (.B1(_00599_),
    .Y(_00600_),
    .A1(net2725),
    .A2(net2760));
 sg13g2_a21oi_1 _10963_ (.A1(net2460),
    .A2(net2570),
    .Y(_00601_),
    .B1(_00600_));
 sg13g2_xor2_1 _10964_ (.B(net2200),
    .A(net2389),
    .X(_00602_));
 sg13g2_nor2_1 _10965_ (.A(net2279),
    .B(net2309),
    .Y(_00603_));
 sg13g2_xnor2_1 _10966_ (.Y(_00604_),
    .A(net2711),
    .B(net2618));
 sg13g2_xnor2_1 _10967_ (.Y(_00605_),
    .A(_00603_),
    .B(_00604_));
 sg13g2_nor2b_1 _10968_ (.A(_00605_),
    .B_N(_00602_),
    .Y(_00606_));
 sg13g2_nand2b_1 _10969_ (.Y(_00607_),
    .B(_00605_),
    .A_N(_00602_));
 sg13g2_xnor2_1 _10970_ (.Y(_00608_),
    .A(_00602_),
    .B(_00605_));
 sg13g2_xnor2_1 _10971_ (.Y(_00609_),
    .A(_00601_),
    .B(_00608_));
 sg13g2_xor2_1 _10972_ (.B(net2668),
    .A(net2189),
    .X(_00610_));
 sg13g2_o21ai_1 _10973_ (.B1(_00610_),
    .Y(_00611_),
    .A1(net2570),
    .A2(net2502));
 sg13g2_xnor2_1 _10974_ (.Y(_00612_),
    .A(net2734),
    .B(net2711));
 sg13g2_xnor2_1 _10975_ (.Y(_00613_),
    .A(net2311),
    .B(_00612_));
 sg13g2_nor2b_1 _10976_ (.A(net2322),
    .B_N(net2467),
    .Y(_00614_));
 sg13g2_nor2_1 _10977_ (.A(net2457),
    .B(net2409),
    .Y(_00615_));
 sg13g2_xnor2_1 _10978_ (.Y(_00616_),
    .A(_00614_),
    .B(_00615_));
 sg13g2_nor2_1 _10979_ (.A(_00613_),
    .B(_00616_),
    .Y(_00617_));
 sg13g2_nand2_1 _10980_ (.Y(_00618_),
    .A(_00613_),
    .B(_00616_));
 sg13g2_xnor2_1 _10981_ (.Y(_00619_),
    .A(_00613_),
    .B(_00616_));
 sg13g2_o21ai_1 _10982_ (.B1(_00618_),
    .Y(_00620_),
    .A1(_00611_),
    .A2(_00617_));
 sg13g2_xnor2_1 _10983_ (.Y(_00621_),
    .A(_00611_),
    .B(_00619_));
 sg13g2_nand2_1 _10984_ (.Y(_00622_),
    .A(_00609_),
    .B(_00621_));
 sg13g2_or2_1 _10985_ (.X(_00623_),
    .B(_00621_),
    .A(_00609_));
 sg13g2_xor2_1 _10986_ (.B(_00621_),
    .A(_00609_),
    .X(_00624_));
 sg13g2_xor2_1 _10987_ (.B(net2598),
    .A(net2586),
    .X(_00625_));
 sg13g2_xnor2_1 _10988_ (.Y(_00626_),
    .A(net2453),
    .B(net2656));
 sg13g2_nand2_1 _10989_ (.Y(_00627_),
    .A(_00625_),
    .B(_00626_));
 sg13g2_xor2_1 _10990_ (.B(net2562),
    .A(net2453),
    .X(_00628_));
 sg13g2_nand2_1 _10991_ (.Y(_00629_),
    .A(_08509_),
    .B(_00628_));
 sg13g2_nor2_1 _10992_ (.A(net2304),
    .B(net2481),
    .Y(_00630_));
 sg13g2_xnor2_1 _10993_ (.Y(_00631_),
    .A(net2389),
    .B(_00630_));
 sg13g2_nand2b_1 _10994_ (.Y(_00632_),
    .B(_00631_),
    .A_N(_00629_));
 sg13g2_nor2b_1 _10995_ (.A(_00631_),
    .B_N(_00629_),
    .Y(_00633_));
 sg13g2_xnor2_1 _10996_ (.Y(_00634_),
    .A(_00629_),
    .B(_00631_));
 sg13g2_xnor2_1 _10997_ (.Y(_00635_),
    .A(_00627_),
    .B(_00634_));
 sg13g2_xnor2_1 _10998_ (.Y(_00636_),
    .A(_00624_),
    .B(_00635_));
 sg13g2_nor2_1 _10999_ (.A(_00598_),
    .B(_00636_),
    .Y(_00637_));
 sg13g2_and2_1 _11000_ (.A(_00598_),
    .B(_00636_),
    .X(_00638_));
 sg13g2_nor2_1 _11001_ (.A(_00637_),
    .B(_00638_),
    .Y(_00639_));
 sg13g2_xnor2_1 _11002_ (.Y(_00640_),
    .A(_00562_),
    .B(_00639_));
 sg13g2_o21ai_1 _11003_ (.B1(_00640_),
    .Y(_00641_),
    .A1(_09576_),
    .A2(_00522_));
 sg13g2_xnor2_1 _11004_ (.Y(_00642_),
    .A(_00524_),
    .B(_00640_));
 sg13g2_xnor2_1 _11005_ (.Y(_00643_),
    .A(_08223_),
    .B(_00642_));
 sg13g2_xnor2_1 _11006_ (.Y(_00644_),
    .A(net2418),
    .B(net2509));
 sg13g2_xnor2_1 _11007_ (.Y(_00645_),
    .A(net2390),
    .B(net2439));
 sg13g2_nand2b_1 _11008_ (.Y(_00646_),
    .B(net2209),
    .A_N(net2200));
 sg13g2_xnor2_1 _11009_ (.Y(_00647_),
    .A(\net.in[209] ),
    .B(net2409));
 sg13g2_xnor2_1 _11010_ (.Y(_00648_),
    .A(_00646_),
    .B(_00647_));
 sg13g2_nand2b_1 _11011_ (.Y(_00649_),
    .B(_00645_),
    .A_N(_00648_));
 sg13g2_nand2b_1 _11012_ (.Y(_00650_),
    .B(_00648_),
    .A_N(_00645_));
 sg13g2_xnor2_1 _11013_ (.Y(_00651_),
    .A(_00645_),
    .B(_00648_));
 sg13g2_nand2b_1 _11014_ (.Y(_00652_),
    .B(_00649_),
    .A_N(_00644_));
 sg13g2_xnor2_1 _11015_ (.Y(_00653_),
    .A(_00644_),
    .B(_00651_));
 sg13g2_nand2_1 _11016_ (.Y(_00654_),
    .A(net2299),
    .B(net2207));
 sg13g2_xnor2_1 _11017_ (.Y(_00655_),
    .A(net2367),
    .B(_00654_));
 sg13g2_nor2_1 _11018_ (.A(net2367),
    .B(net2320),
    .Y(_00656_));
 sg13g2_nor3_2 _11019_ (.A(net2570),
    .B(net2605),
    .C(_00656_),
    .Y(_00657_));
 sg13g2_xor2_1 _11020_ (.B(net2319),
    .A(net2409),
    .X(_00658_));
 sg13g2_nor2_1 _11021_ (.A(net2211),
    .B(_00658_),
    .Y(_00659_));
 sg13g2_nand2b_1 _11022_ (.Y(_00660_),
    .B(_00659_),
    .A_N(_00657_));
 sg13g2_nor2b_1 _11023_ (.A(_00659_),
    .B_N(_00657_),
    .Y(_00661_));
 sg13g2_xor2_1 _11024_ (.B(_00659_),
    .A(_00657_),
    .X(_00662_));
 sg13g2_xnor2_1 _11025_ (.Y(_00663_),
    .A(_00655_),
    .B(_00662_));
 sg13g2_nand2b_1 _11026_ (.Y(_00664_),
    .B(_00663_),
    .A_N(_00653_));
 sg13g2_nor2b_1 _11027_ (.A(_00663_),
    .B_N(_00653_),
    .Y(_00665_));
 sg13g2_nand2b_2 _11028_ (.Y(_00666_),
    .B(net2634),
    .A_N(net2711));
 sg13g2_nor2_2 _11029_ (.A(net2515),
    .B(_05869_),
    .Y(_00667_));
 sg13g2_xnor2_1 _11030_ (.Y(_00668_),
    .A(_00666_),
    .B(_00667_));
 sg13g2_nor2b_1 _11031_ (.A(net2534),
    .B_N(net2566),
    .Y(_00669_));
 sg13g2_nor3_2 _11032_ (.A(net2341),
    .B(net2656),
    .C(_00669_),
    .Y(_00670_));
 sg13g2_nor2_1 _11033_ (.A(net2481),
    .B(net2662),
    .Y(_00671_));
 sg13g2_nor2_1 _11034_ (.A(net2393),
    .B(net2281),
    .Y(_00672_));
 sg13g2_xnor2_1 _11035_ (.Y(_00673_),
    .A(_00671_),
    .B(_00672_));
 sg13g2_nor2b_1 _11036_ (.A(_00673_),
    .B_N(_00670_),
    .Y(_00674_));
 sg13g2_nand2b_1 _11037_ (.Y(_00675_),
    .B(_00673_),
    .A_N(_00670_));
 sg13g2_nand2b_1 _11038_ (.Y(_00676_),
    .B(_00675_),
    .A_N(_00674_));
 sg13g2_xor2_1 _11039_ (.B(_00676_),
    .A(_00668_),
    .X(_00677_));
 sg13g2_a21oi_2 _11040_ (.B1(_00665_),
    .Y(_00678_),
    .A2(_00677_),
    .A1(_00664_));
 sg13g2_nand2_1 _11041_ (.Y(_00679_),
    .A(_05077_),
    .B(net2252));
 sg13g2_xnor2_1 _11042_ (.Y(_00680_),
    .A(\net.in[10] ),
    .B(net2222));
 sg13g2_xnor2_1 _11043_ (.Y(_00681_),
    .A(_00679_),
    .B(_00680_));
 sg13g2_nor2_1 _11044_ (.A(net2796),
    .B(net2253),
    .Y(_00682_));
 sg13g2_xnor2_1 _11045_ (.Y(_00683_),
    .A(_00013_),
    .B(_00682_));
 sg13g2_nand2_1 _11046_ (.Y(_00684_),
    .A(_00435_),
    .B(_00683_));
 sg13g2_xnor2_1 _11047_ (.Y(_00685_),
    .A(_00439_),
    .B(_00683_));
 sg13g2_o21ai_1 _11048_ (.B1(_00681_),
    .Y(_00686_),
    .A1(_00435_),
    .A2(_00683_));
 sg13g2_xor2_1 _11049_ (.B(_00685_),
    .A(_00681_),
    .X(_00687_));
 sg13g2_nor2_1 _11050_ (.A(net2525),
    .B(net2575),
    .Y(_00688_));
 sg13g2_nor2b_1 _11051_ (.A(net2282),
    .B_N(net2418),
    .Y(_00689_));
 sg13g2_xnor2_1 _11052_ (.Y(_00690_),
    .A(net2332),
    .B(_00689_));
 sg13g2_nor2_1 _11053_ (.A(net2295),
    .B(net2381),
    .Y(_00691_));
 sg13g2_nor2_1 _11054_ (.A(net2606),
    .B(net2596),
    .Y(_00692_));
 sg13g2_xor2_1 _11055_ (.B(_00692_),
    .A(_00691_),
    .X(_00693_));
 sg13g2_nand2_1 _11056_ (.Y(_00694_),
    .A(_00690_),
    .B(_00693_));
 sg13g2_xnor2_1 _11057_ (.Y(_00695_),
    .A(_00690_),
    .B(_00693_));
 sg13g2_xnor2_1 _11058_ (.Y(_00696_),
    .A(_00688_),
    .B(_00695_));
 sg13g2_nand2_1 _11059_ (.Y(_00697_),
    .A(_00687_),
    .B(_00696_));
 sg13g2_xor2_1 _11060_ (.B(net2502),
    .A(net2558),
    .X(_00698_));
 sg13g2_nand2_2 _11061_ (.Y(_00699_),
    .A(_05693_),
    .B(_05979_));
 sg13g2_a21oi_1 _11062_ (.A1(net2581),
    .A2(net2638),
    .Y(_00700_),
    .B1(net2492));
 sg13g2_xnor2_1 _11063_ (.Y(_00701_),
    .A(net2336),
    .B(net2222));
 sg13g2_a21oi_1 _11064_ (.A1(_00699_),
    .A2(_00700_),
    .Y(_00702_),
    .B1(_00701_));
 sg13g2_inv_1 _11065_ (.Y(_00703_),
    .A(_00702_));
 sg13g2_and3_1 _11066_ (.X(_00704_),
    .A(_00699_),
    .B(_00700_),
    .C(_00701_));
 sg13g2_nor2_1 _11067_ (.A(_00702_),
    .B(_00704_),
    .Y(_00705_));
 sg13g2_xor2_1 _11068_ (.B(_00705_),
    .A(_00698_),
    .X(_00706_));
 sg13g2_or2_1 _11069_ (.X(_00707_),
    .B(_00696_),
    .A(_00687_));
 sg13g2_nand2_1 _11070_ (.Y(_00708_),
    .A(_00697_),
    .B(_00706_));
 sg13g2_nor2_1 _11071_ (.A(net2211),
    .B(net2362),
    .Y(_00709_));
 sg13g2_nor2_1 _11072_ (.A(net2187),
    .B(net2796),
    .Y(_00710_));
 sg13g2_xnor2_1 _11073_ (.Y(_00711_),
    .A(_00709_),
    .B(_00710_));
 sg13g2_o21ai_1 _11074_ (.B1(net2581),
    .Y(_00712_),
    .A1(net2694),
    .A2(net2740));
 sg13g2_or3_1 _11075_ (.A(net2694),
    .B(net2740),
    .C(net2581),
    .X(_00713_));
 sg13g2_xor2_1 _11076_ (.B(net2623),
    .A(net2807),
    .X(_00714_));
 sg13g2_a21oi_1 _11077_ (.A1(_00712_),
    .A2(_00713_),
    .Y(_00715_),
    .B1(_00714_));
 sg13g2_nand3_1 _11078_ (.B(_00713_),
    .C(_00714_),
    .A(_00712_),
    .Y(_00716_));
 sg13g2_nand2b_1 _11079_ (.Y(_00717_),
    .B(_00716_),
    .A_N(_00715_));
 sg13g2_xor2_1 _11080_ (.B(_00717_),
    .A(_00711_),
    .X(_00718_));
 sg13g2_nor2_1 _11081_ (.A(net2409),
    .B(net2211),
    .Y(_00719_));
 sg13g2_xor2_1 _11082_ (.B(net2743),
    .A(net2800),
    .X(_00720_));
 sg13g2_xnor2_1 _11083_ (.Y(_00721_),
    .A(_00719_),
    .B(_00720_));
 sg13g2_xnor2_1 _11084_ (.Y(_00722_),
    .A(net2364),
    .B(net2702));
 sg13g2_nand2_1 _11085_ (.Y(_00723_),
    .A(net2269),
    .B(net2220));
 sg13g2_or2_1 _11086_ (.X(_00724_),
    .B(net2220),
    .A(net2269));
 sg13g2_nand3_1 _11087_ (.B(_00723_),
    .C(_00724_),
    .A(_00722_),
    .Y(_00725_));
 sg13g2_nor2_1 _11088_ (.A(net2189),
    .B(net2252),
    .Y(_00726_));
 sg13g2_xor2_1 _11089_ (.B(_00726_),
    .A(_00724_),
    .X(_00727_));
 sg13g2_xnor2_1 _11090_ (.Y(_00728_),
    .A(_00725_),
    .B(_00727_));
 sg13g2_a21o_1 _11091_ (.A2(_00727_),
    .A1(_00725_),
    .B1(_00721_),
    .X(_00729_));
 sg13g2_o21ai_1 _11092_ (.B1(_00729_),
    .Y(_00730_),
    .A1(_00725_),
    .A2(_00727_));
 sg13g2_xnor2_1 _11093_ (.Y(_00731_),
    .A(_00721_),
    .B(_00728_));
 sg13g2_nand2_1 _11094_ (.Y(_00732_),
    .A(_00718_),
    .B(_00731_));
 sg13g2_xnor2_1 _11095_ (.Y(_00733_),
    .A(net2289),
    .B(net2224));
 sg13g2_xor2_1 _11096_ (.B(net2623),
    .A(net2525),
    .X(_00734_));
 sg13g2_xnor2_1 _11097_ (.Y(_00735_),
    .A(net2558),
    .B(net2656));
 sg13g2_nor2b_1 _11098_ (.A(net2299),
    .B_N(net2291),
    .Y(_00736_));
 sg13g2_nor2b_1 _11099_ (.A(net2248),
    .B_N(net2226),
    .Y(_00737_));
 sg13g2_xnor2_1 _11100_ (.Y(_00738_),
    .A(_00736_),
    .B(_00737_));
 sg13g2_a21oi_1 _11101_ (.A1(_00734_),
    .A2(_00735_),
    .Y(_00739_),
    .B1(_00738_));
 sg13g2_nand3_1 _11102_ (.B(_00735_),
    .C(_00738_),
    .A(_00734_),
    .Y(_00740_));
 sg13g2_nor2b_1 _11103_ (.A(_00739_),
    .B_N(_00740_),
    .Y(_00741_));
 sg13g2_xnor2_1 _11104_ (.Y(_00742_),
    .A(_00733_),
    .B(_00741_));
 sg13g2_or2_1 _11105_ (.X(_00743_),
    .B(_00731_),
    .A(_00718_));
 sg13g2_nand2_1 _11106_ (.Y(_00744_),
    .A(_00732_),
    .B(_00742_));
 sg13g2_a22oi_1 _11107_ (.Y(_00745_),
    .B1(_00743_),
    .B2(_00744_),
    .A2(_00708_),
    .A1(_00707_));
 sg13g2_inv_1 _11108_ (.Y(_00746_),
    .A(_00745_));
 sg13g2_and4_1 _11109_ (.A(_00707_),
    .B(_00708_),
    .C(_00743_),
    .D(_00744_),
    .X(_00747_));
 sg13g2_a21oi_1 _11110_ (.A1(_00678_),
    .A2(_00746_),
    .Y(_00748_),
    .B1(_00747_));
 sg13g2_a21o_1 _11111_ (.A2(_00747_),
    .A1(_00678_),
    .B1(_00748_),
    .X(_00749_));
 sg13g2_o21ai_1 _11112_ (.B1(_00749_),
    .Y(_00750_),
    .A1(_00678_),
    .A2(_00746_));
 sg13g2_nor2_2 _11113_ (.A(net2816),
    .B(\net.in[208] ),
    .Y(_00751_));
 sg13g2_and2_1 _11114_ (.A(net2816),
    .B(\net.in[208] ),
    .X(_00752_));
 sg13g2_xnor2_1 _11115_ (.Y(_00753_),
    .A(net2806),
    .B(net2211));
 sg13g2_o21ai_1 _11116_ (.B1(_00753_),
    .Y(_00754_),
    .A1(_00751_),
    .A2(_00752_));
 sg13g2_nand2_1 _11117_ (.Y(_00755_),
    .A(net2259),
    .B(net2270));
 sg13g2_nor2_1 _11118_ (.A(net2457),
    .B(net2408),
    .Y(_00756_));
 sg13g2_xor2_1 _11119_ (.B(_00756_),
    .A(_00755_),
    .X(_00757_));
 sg13g2_nand2b_1 _11120_ (.Y(_00758_),
    .B(_00757_),
    .A_N(_07431_));
 sg13g2_nand2b_1 _11121_ (.Y(_00759_),
    .B(_07431_),
    .A_N(_00757_));
 sg13g2_xor2_1 _11122_ (.B(_00757_),
    .A(_07431_),
    .X(_00760_));
 sg13g2_xnor2_1 _11123_ (.Y(_00761_),
    .A(_00754_),
    .B(_00760_));
 sg13g2_nor2_2 _11124_ (.A(net2183),
    .B(net2727),
    .Y(_00762_));
 sg13g2_nor2_1 _11125_ (.A(net2555),
    .B(net2609),
    .Y(_00763_));
 sg13g2_xnor2_1 _11126_ (.Y(_00764_),
    .A(_00762_),
    .B(_00763_));
 sg13g2_xor2_1 _11127_ (.B(net2809),
    .A(net2359),
    .X(_00765_));
 sg13g2_xnor2_1 _11128_ (.Y(_00766_),
    .A(net2359),
    .B(net2809));
 sg13g2_nor2b_1 _11129_ (.A(net2606),
    .B_N(net2666),
    .Y(_00767_));
 sg13g2_nor2b_1 _11130_ (.A(net2666),
    .B_N(net2606),
    .Y(_00768_));
 sg13g2_nor2b_1 _11131_ (.A(net2674),
    .B_N(net2426),
    .Y(_00769_));
 sg13g2_nor3_2 _11132_ (.A(_00767_),
    .B(_00768_),
    .C(_00769_),
    .Y(_00770_));
 sg13g2_nand2_1 _11133_ (.Y(_00771_),
    .A(_00765_),
    .B(_00770_));
 sg13g2_nor2_1 _11134_ (.A(_00765_),
    .B(_00770_),
    .Y(_00772_));
 sg13g2_xnor2_1 _11135_ (.Y(_00773_),
    .A(_00766_),
    .B(_00770_));
 sg13g2_xnor2_1 _11136_ (.Y(_00774_),
    .A(_00764_),
    .B(_00773_));
 sg13g2_nand2_1 _11137_ (.Y(_00775_),
    .A(_00761_),
    .B(_00774_));
 sg13g2_nor2_1 _11138_ (.A(net2482),
    .B(net2525),
    .Y(_00776_));
 sg13g2_nor2_1 _11139_ (.A(net2592),
    .B(net2646),
    .Y(_00777_));
 sg13g2_xnor2_1 _11140_ (.Y(_00778_),
    .A(_00776_),
    .B(_00777_));
 sg13g2_nor2_1 _11141_ (.A(net2398),
    .B(net2221),
    .Y(_00779_));
 sg13g2_xnor2_1 _11142_ (.Y(_00780_),
    .A(net2517),
    .B(_00779_));
 sg13g2_xor2_1 _11143_ (.B(net2513),
    .A(net2336),
    .X(_00781_));
 sg13g2_nand3b_1 _11144_ (.B(_06078_),
    .C(_00781_),
    .Y(_00782_),
    .A_N(net2493));
 sg13g2_nand2_1 _11145_ (.Y(_00783_),
    .A(_00780_),
    .B(_00782_));
 sg13g2_or2_1 _11146_ (.X(_00784_),
    .B(_00782_),
    .A(_00780_));
 sg13g2_nand2_1 _11147_ (.Y(_00785_),
    .A(_00783_),
    .B(_00784_));
 sg13g2_xnor2_1 _11148_ (.Y(_00786_),
    .A(_00778_),
    .B(_00785_));
 sg13g2_or2_1 _11149_ (.X(_00787_),
    .B(_00774_),
    .A(_00761_));
 sg13g2_nand2_1 _11150_ (.Y(_00788_),
    .A(_00775_),
    .B(_00786_));
 sg13g2_xnor2_1 _11151_ (.Y(_00789_),
    .A(net2539),
    .B(net2592));
 sg13g2_xor2_1 _11152_ (.B(net2237),
    .A(net2492),
    .X(_00790_));
 sg13g2_nor2_1 _11153_ (.A(_00789_),
    .B(_00790_),
    .Y(_00791_));
 sg13g2_nor2_1 _11154_ (.A(net2311),
    .B(net2189),
    .Y(_00792_));
 sg13g2_xor2_1 _11155_ (.B(net2218),
    .A(net2304),
    .X(_00793_));
 sg13g2_xnor2_1 _11156_ (.Y(_00794_),
    .A(_00792_),
    .B(_00793_));
 sg13g2_nand2_1 _11157_ (.Y(_00795_),
    .A(_00791_),
    .B(_00794_));
 sg13g2_nor2_1 _11158_ (.A(_00791_),
    .B(_00794_),
    .Y(_00796_));
 sg13g2_xnor2_1 _11159_ (.Y(_00797_),
    .A(_00791_),
    .B(_00794_));
 sg13g2_nand2_1 _11160_ (.Y(_00798_),
    .A(net2575),
    .B(net2635));
 sg13g2_o21ai_1 _11161_ (.B1(_00798_),
    .Y(_00799_),
    .A1(net2635),
    .A2(_06177_));
 sg13g2_xnor2_1 _11162_ (.Y(_00800_),
    .A(_00797_),
    .B(_00799_));
 sg13g2_nand2_1 _11163_ (.Y(_00801_),
    .A(net2674),
    .B(net2364));
 sg13g2_or2_1 _11164_ (.X(_00802_),
    .B(net2364),
    .A(net2674));
 sg13g2_nand2b_1 _11165_ (.Y(_00803_),
    .B(net2606),
    .A_N(net2407));
 sg13g2_and2_1 _11166_ (.A(_00801_),
    .B(_00803_),
    .X(_00804_));
 sg13g2_nand3_1 _11167_ (.B(_00802_),
    .C(_00803_),
    .A(_00801_),
    .Y(_00805_));
 sg13g2_nor2_1 _11168_ (.A(net2448),
    .B(net2677),
    .Y(_00806_));
 sg13g2_xor2_1 _11169_ (.B(net2237),
    .A(net2488),
    .X(_00807_));
 sg13g2_xnor2_1 _11170_ (.Y(_00808_),
    .A(_00806_),
    .B(_00807_));
 sg13g2_a21oi_1 _11171_ (.A1(_00802_),
    .A2(_00804_),
    .Y(_00809_),
    .B1(_00808_));
 sg13g2_nand2b_1 _11172_ (.Y(_00810_),
    .B(_00808_),
    .A_N(_00805_));
 sg13g2_xnor2_1 _11173_ (.Y(_00811_),
    .A(_00805_),
    .B(_00808_));
 sg13g2_xor2_1 _11174_ (.B(net2339),
    .A(net2346),
    .X(_00812_));
 sg13g2_nor2_1 _11175_ (.A(net2406),
    .B(net2210),
    .Y(_00813_));
 sg13g2_xnor2_1 _11176_ (.Y(_00814_),
    .A(_00812_),
    .B(_00813_));
 sg13g2_xnor2_1 _11177_ (.Y(_00815_),
    .A(_00811_),
    .B(_00814_));
 sg13g2_nand2_1 _11178_ (.Y(_00816_),
    .A(_00800_),
    .B(_00815_));
 sg13g2_xor2_1 _11179_ (.B(net2571),
    .A(net2483),
    .X(_00817_));
 sg13g2_xnor2_1 _11180_ (.Y(_00818_),
    .A(net2521),
    .B(_00817_));
 sg13g2_xnor2_1 _11181_ (.Y(_00819_),
    .A(net2743),
    .B(\net.in[208] ));
 sg13g2_nand2b_1 _11182_ (.Y(_00820_),
    .B(_00819_),
    .A_N(_06254_));
 sg13g2_xnor2_1 _11183_ (.Y(_00821_),
    .A(net2478),
    .B(net2579));
 sg13g2_xnor2_1 _11184_ (.Y(_00822_),
    .A(net2659),
    .B(net2239));
 sg13g2_nand2_2 _11185_ (.Y(_00823_),
    .A(_00821_),
    .B(_00822_));
 sg13g2_nand2b_1 _11186_ (.Y(_00824_),
    .B(_00823_),
    .A_N(_00820_));
 sg13g2_nand2b_1 _11187_ (.Y(_00825_),
    .B(_00820_),
    .A_N(_00823_));
 sg13g2_and2_1 _11188_ (.A(_00824_),
    .B(_00825_),
    .X(_00826_));
 sg13g2_xnor2_1 _11189_ (.Y(_00827_),
    .A(_00818_),
    .B(_00826_));
 sg13g2_or2_1 _11190_ (.X(_00828_),
    .B(_00815_),
    .A(_00800_));
 sg13g2_nand2_1 _11191_ (.Y(_00829_),
    .A(_00816_),
    .B(_00827_));
 sg13g2_a22oi_1 _11192_ (.Y(_00830_),
    .B1(_00828_),
    .B2(_00829_),
    .A2(_00788_),
    .A1(_00787_));
 sg13g2_and4_1 _11193_ (.A(_00787_),
    .B(_00788_),
    .C(_00828_),
    .D(_00829_),
    .X(_00831_));
 sg13g2_inv_1 _11194_ (.Y(_00832_),
    .A(_00831_));
 sg13g2_nor2_1 _11195_ (.A(_00830_),
    .B(_00831_),
    .Y(_00833_));
 sg13g2_nor2_1 _11196_ (.A(_05055_),
    .B(net2235),
    .Y(_00834_));
 sg13g2_xnor2_1 _11197_ (.Y(_00835_),
    .A(net2291),
    .B(_00834_));
 sg13g2_xor2_1 _11198_ (.B(net2638),
    .A(net2354),
    .X(_00836_));
 sg13g2_nor2_1 _11199_ (.A(net2471),
    .B(net2467),
    .Y(_00837_));
 sg13g2_xnor2_1 _11200_ (.Y(_00838_),
    .A(net2457),
    .B(net2209));
 sg13g2_xnor2_1 _11201_ (.Y(_00839_),
    .A(_00837_),
    .B(_00838_));
 sg13g2_nor2_1 _11202_ (.A(_00836_),
    .B(_00839_),
    .Y(_00840_));
 sg13g2_xor2_1 _11203_ (.B(_00839_),
    .A(_00836_),
    .X(_00841_));
 sg13g2_xnor2_1 _11204_ (.Y(_00842_),
    .A(_00835_),
    .B(_00841_));
 sg13g2_nor2_2 _11205_ (.A(net2224),
    .B(net2197),
    .Y(_00843_));
 sg13g2_xnor2_1 _11206_ (.Y(_00844_),
    .A(net2550),
    .B(net2212));
 sg13g2_xnor2_1 _11207_ (.Y(_00845_),
    .A(_00843_),
    .B(_00844_));
 sg13g2_nand2_1 _11208_ (.Y(_00846_),
    .A(net2677),
    .B(net2245));
 sg13g2_xor2_1 _11209_ (.B(net2246),
    .A(net2681),
    .X(_00847_));
 sg13g2_a21o_1 _11210_ (.A2(net2398),
    .A1(_05319_),
    .B1(_00847_),
    .X(_00848_));
 sg13g2_nand2_1 _11211_ (.Y(_00849_),
    .A(net2218),
    .B(net2291));
 sg13g2_xor2_1 _11212_ (.B(net2310),
    .A(net2299),
    .X(_00850_));
 sg13g2_xnor2_1 _11213_ (.Y(_00851_),
    .A(_00849_),
    .B(_00850_));
 sg13g2_nand2b_1 _11214_ (.Y(_00852_),
    .B(_00848_),
    .A_N(_00851_));
 sg13g2_nand2b_1 _11215_ (.Y(_00853_),
    .B(_00851_),
    .A_N(_00848_));
 sg13g2_xnor2_1 _11216_ (.Y(_00854_),
    .A(_00848_),
    .B(_00851_));
 sg13g2_xnor2_1 _11217_ (.Y(_00855_),
    .A(_00845_),
    .B(_00854_));
 sg13g2_nor2_1 _11218_ (.A(_00842_),
    .B(_00855_),
    .Y(_00856_));
 sg13g2_nor2_1 _11219_ (.A(net2772),
    .B(net2320),
    .Y(_00857_));
 sg13g2_xnor2_1 _11220_ (.Y(_00858_),
    .A(net2367),
    .B(_00857_));
 sg13g2_xnor2_1 _11221_ (.Y(_00859_),
    .A(net2190),
    .B(net2220));
 sg13g2_nor2_1 _11222_ (.A(net2455),
    .B(\net.in[225] ),
    .Y(_00860_));
 sg13g2_nor2_1 _11223_ (.A(net2791),
    .B(\net.in[192] ),
    .Y(_00861_));
 sg13g2_xor2_1 _11224_ (.B(_00861_),
    .A(_00860_),
    .X(_00862_));
 sg13g2_nand2_2 _11225_ (.Y(_00863_),
    .A(_00859_),
    .B(_00862_));
 sg13g2_or2_1 _11226_ (.X(_00864_),
    .B(_00862_),
    .A(_00859_));
 sg13g2_nand2_1 _11227_ (.Y(_00865_),
    .A(_00863_),
    .B(_00864_));
 sg13g2_xnor2_1 _11228_ (.Y(_00866_),
    .A(_00858_),
    .B(_00865_));
 sg13g2_nand2_1 _11229_ (.Y(_00867_),
    .A(_00842_),
    .B(_00855_));
 sg13g2_o21ai_1 _11230_ (.B1(_00867_),
    .Y(_00868_),
    .A1(_00856_),
    .A2(_00866_));
 sg13g2_xor2_1 _11231_ (.B(_00868_),
    .A(_00833_),
    .X(_00869_));
 sg13g2_nor2_1 _11232_ (.A(_00750_),
    .B(_00869_),
    .Y(_00870_));
 sg13g2_nand2_1 _11233_ (.Y(_00871_),
    .A(_00750_),
    .B(_00869_));
 sg13g2_nand2_1 _11234_ (.Y(_00872_),
    .A(net2325),
    .B(net2412));
 sg13g2_o21ai_1 _11235_ (.B1(_00872_),
    .Y(_00873_),
    .A1(net2388),
    .A2(net2393));
 sg13g2_xnor2_1 _11236_ (.Y(_00874_),
    .A(net2668),
    .B(net2682));
 sg13g2_nand2_1 _11237_ (.Y(_00875_),
    .A(net2243),
    .B(net2534));
 sg13g2_xnor2_1 _11238_ (.Y(_00876_),
    .A(_00874_),
    .B(_00875_));
 sg13g2_nor2b_1 _11239_ (.A(net2484),
    .B_N(net2481),
    .Y(_00877_));
 sg13g2_nor2_1 _11240_ (.A(net2311),
    .B(net2586),
    .Y(_00878_));
 sg13g2_xnor2_1 _11241_ (.Y(_00879_),
    .A(_00877_),
    .B(_00878_));
 sg13g2_nor2b_1 _11242_ (.A(_00876_),
    .B_N(_00879_),
    .Y(_00880_));
 sg13g2_nand2b_1 _11243_ (.Y(_00881_),
    .B(_00876_),
    .A_N(_00879_));
 sg13g2_xnor2_1 _11244_ (.Y(_00882_),
    .A(_00876_),
    .B(_00879_));
 sg13g2_xnor2_1 _11245_ (.Y(_00883_),
    .A(_00873_),
    .B(_00882_));
 sg13g2_xnor2_1 _11246_ (.Y(_00884_),
    .A(net2481),
    .B(net2434));
 sg13g2_xnor2_1 _11247_ (.Y(_00885_),
    .A(net2521),
    .B(_00884_));
 sg13g2_xnor2_1 _11248_ (.Y(_00886_),
    .A(net2652),
    .B(net2570));
 sg13g2_xnor2_1 _11249_ (.Y(_00887_),
    .A(net2656),
    .B(net2605));
 sg13g2_nor4_2 _11250_ (.A(net2482),
    .B(net2484),
    .C(net2525),
    .Y(_00888_),
    .D(net2570));
 sg13g2_nand3_1 _11251_ (.B(_00887_),
    .C(_00888_),
    .A(_00886_),
    .Y(_00889_));
 sg13g2_a21oi_1 _11252_ (.A1(_00886_),
    .A2(_00887_),
    .Y(_00890_),
    .B1(_00888_));
 sg13g2_a21o_1 _11253_ (.A2(_00887_),
    .A1(_00886_),
    .B1(_00888_),
    .X(_00891_));
 sg13g2_nand2_1 _11254_ (.Y(_00892_),
    .A(_00889_),
    .B(_00891_));
 sg13g2_xnor2_1 _11255_ (.Y(_00893_),
    .A(_00885_),
    .B(_00892_));
 sg13g2_or2_1 _11256_ (.X(_00894_),
    .B(_00893_),
    .A(_00883_));
 sg13g2_xnor2_1 _11257_ (.Y(_00895_),
    .A(net2417),
    .B(net2512));
 sg13g2_or2_1 _11258_ (.X(_00896_),
    .B(net2600),
    .A(net2350));
 sg13g2_nor2b_1 _11259_ (.A(net2488),
    .B_N(net2480),
    .Y(_00897_));
 sg13g2_xnor2_1 _11260_ (.Y(_00898_),
    .A(net2201),
    .B(net2257));
 sg13g2_nor2_1 _11261_ (.A(net2390),
    .B(net2692),
    .Y(_00899_));
 sg13g2_xnor2_1 _11262_ (.Y(_00900_),
    .A(_00898_),
    .B(_00899_));
 sg13g2_a21oi_1 _11263_ (.A1(_00896_),
    .A2(_00897_),
    .Y(_00901_),
    .B1(_00900_));
 sg13g2_nand3_1 _11264_ (.B(_00897_),
    .C(_00900_),
    .A(_00896_),
    .Y(_00902_));
 sg13g2_nand2b_1 _11265_ (.Y(_00903_),
    .B(_00902_),
    .A_N(_00901_));
 sg13g2_xnor2_1 _11266_ (.Y(_00904_),
    .A(_00895_),
    .B(_00903_));
 sg13g2_nand2_1 _11267_ (.Y(_00905_),
    .A(_00883_),
    .B(_00893_));
 sg13g2_nand2_1 _11268_ (.Y(_00906_),
    .A(_00904_),
    .B(_00905_));
 sg13g2_nand2_1 _11269_ (.Y(_00907_),
    .A(_05286_),
    .B(net2356));
 sg13g2_nor2_1 _11270_ (.A(net2361),
    .B(net2208),
    .Y(_00908_));
 sg13g2_xnor2_1 _11271_ (.Y(_00909_),
    .A(_00907_),
    .B(_00908_));
 sg13g2_xnor2_1 _11272_ (.Y(_00910_),
    .A(net2346),
    .B(net2395));
 sg13g2_xor2_1 _11273_ (.B(net2369),
    .A(net2515),
    .X(_00911_));
 sg13g2_nor2_1 _11274_ (.A(_00910_),
    .B(_00911_),
    .Y(_00912_));
 sg13g2_nand2_1 _11275_ (.Y(_00913_),
    .A(_00910_),
    .B(_00911_));
 sg13g2_nor2b_1 _11276_ (.A(_00912_),
    .B_N(_00913_),
    .Y(_00914_));
 sg13g2_xnor2_1 _11277_ (.Y(_00915_),
    .A(_00909_),
    .B(_00914_));
 sg13g2_xor2_1 _11278_ (.B(net2501),
    .A(net2416),
    .X(_00916_));
 sg13g2_nand2_1 _11279_ (.Y(_00917_),
    .A(_05187_),
    .B(net2322));
 sg13g2_nand2b_1 _11280_ (.Y(_00918_),
    .B(net2426),
    .A_N(net2248));
 sg13g2_xnor2_1 _11281_ (.Y(_00919_),
    .A(net2345),
    .B(net2187));
 sg13g2_xnor2_1 _11282_ (.Y(_00920_),
    .A(_00918_),
    .B(_00919_));
 sg13g2_a21oi_1 _11283_ (.A1(_00751_),
    .A2(_00917_),
    .Y(_00921_),
    .B1(_00920_));
 sg13g2_nand3_1 _11284_ (.B(_00917_),
    .C(_00920_),
    .A(_00751_),
    .Y(_00922_));
 sg13g2_nand2b_1 _11285_ (.Y(_00923_),
    .B(_00922_),
    .A_N(_00921_));
 sg13g2_xnor2_1 _11286_ (.Y(_00924_),
    .A(_00916_),
    .B(_00923_));
 sg13g2_nand2_1 _11287_ (.Y(_00925_),
    .A(_00915_),
    .B(_00924_));
 sg13g2_xor2_1 _11288_ (.B(net2442),
    .A(net2481),
    .X(_00926_));
 sg13g2_nor2_1 _11289_ (.A(net2694),
    .B(net2700),
    .Y(_00927_));
 sg13g2_nor2_1 _11290_ (.A(net2380),
    .B(net2575),
    .Y(_00928_));
 sg13g2_xnor2_1 _11291_ (.Y(_00929_),
    .A(net2259),
    .B(net2231));
 sg13g2_nor3_1 _11292_ (.A(_00927_),
    .B(_00928_),
    .C(_00929_),
    .Y(_00930_));
 sg13g2_o21ai_1 _11293_ (.B1(_00929_),
    .Y(_00931_),
    .A1(_00927_),
    .A2(_00928_));
 sg13g2_nand2b_1 _11294_ (.Y(_00932_),
    .B(_00931_),
    .A_N(_00930_));
 sg13g2_xnor2_1 _11295_ (.Y(_00933_),
    .A(_00926_),
    .B(_00932_));
 sg13g2_or2_1 _11296_ (.X(_00934_),
    .B(_00924_),
    .A(_00915_));
 sg13g2_nand2b_1 _11297_ (.Y(_00935_),
    .B(_00934_),
    .A_N(_00933_));
 sg13g2_a22oi_1 _11298_ (.Y(_00936_),
    .B1(_00925_),
    .B2(_00935_),
    .A2(_00906_),
    .A1(_00894_));
 sg13g2_and4_1 _11299_ (.A(_00894_),
    .B(_00906_),
    .C(_00925_),
    .D(_00935_),
    .X(_00937_));
 sg13g2_nor2_1 _11300_ (.A(_00936_),
    .B(_00937_),
    .Y(_00938_));
 sg13g2_nor2_1 _11301_ (.A(net2289),
    .B(net2623),
    .Y(_00939_));
 sg13g2_a21oi_1 _11302_ (.A1(net2792),
    .A2(net2717),
    .Y(_00940_),
    .B1(_00939_));
 sg13g2_o21ai_1 _11303_ (.B1(_00940_),
    .Y(_00941_),
    .A1(net2792),
    .A2(net2717));
 sg13g2_xor2_1 _11304_ (.B(net2282),
    .A(net2370),
    .X(_00942_));
 sg13g2_nor3_2 _11305_ (.A(net2743),
    .B(net2496),
    .C(_00942_),
    .Y(_00943_));
 sg13g2_nor2_1 _11306_ (.A(net2448),
    .B(net2816),
    .Y(_00944_));
 sg13g2_nor2_1 _11307_ (.A(net2430),
    .B(net2422),
    .Y(_00945_));
 sg13g2_xor2_1 _11308_ (.B(_00945_),
    .A(_00944_),
    .X(_00946_));
 sg13g2_xnor2_1 _11309_ (.Y(_00947_),
    .A(_00943_),
    .B(_00946_));
 sg13g2_xnor2_1 _11310_ (.Y(_00948_),
    .A(_00941_),
    .B(_00947_));
 sg13g2_xor2_1 _11311_ (.B(net2328),
    .A(net2729),
    .X(_00949_));
 sg13g2_nand2b_1 _11312_ (.Y(_00950_),
    .B(net2315),
    .A_N(net2769));
 sg13g2_nand2b_1 _11313_ (.Y(_00951_),
    .B(net2769),
    .A_N(net2315));
 sg13g2_nand2b_1 _11314_ (.Y(_00952_),
    .B(net2623),
    .A_N(net2220));
 sg13g2_nand3_1 _11315_ (.B(_00951_),
    .C(_00952_),
    .A(_00950_),
    .Y(_00953_));
 sg13g2_xor2_1 _11316_ (.B(net2571),
    .A(net2525),
    .X(_00954_));
 sg13g2_inv_1 _11317_ (.Y(_00955_),
    .A(_00954_));
 sg13g2_nand2_1 _11318_ (.Y(_00956_),
    .A(_00953_),
    .B(_00955_));
 sg13g2_xnor2_1 _11319_ (.Y(_00957_),
    .A(_00953_),
    .B(_00954_));
 sg13g2_xnor2_1 _11320_ (.Y(_00958_),
    .A(_00949_),
    .B(_00957_));
 sg13g2_nor2_1 _11321_ (.A(_00948_),
    .B(_00958_),
    .Y(_00959_));
 sg13g2_nor2_1 _11322_ (.A(net2482),
    .B(net2403),
    .Y(_00960_));
 sg13g2_nor2_1 _11323_ (.A(net2473),
    .B(net2438),
    .Y(_00961_));
 sg13g2_xnor2_1 _11324_ (.Y(_00962_),
    .A(_00960_),
    .B(_00961_));
 sg13g2_xnor2_1 _11325_ (.Y(_00963_),
    .A(net2434),
    .B(net2388));
 sg13g2_nor2_1 _11326_ (.A(net2460),
    .B(net2329),
    .Y(_00964_));
 sg13g2_xnor2_1 _11327_ (.Y(_00965_),
    .A(_07453_),
    .B(_00964_));
 sg13g2_nor2_1 _11328_ (.A(_00963_),
    .B(_00965_),
    .Y(_00966_));
 sg13g2_xor2_1 _11329_ (.B(_00965_),
    .A(_00963_),
    .X(_00967_));
 sg13g2_xnor2_1 _11330_ (.Y(_00968_),
    .A(_00962_),
    .B(_00967_));
 sg13g2_a21oi_1 _11331_ (.A1(_00948_),
    .A2(_00958_),
    .Y(_00969_),
    .B1(_00968_));
 sg13g2_nor2_2 _11332_ (.A(_00959_),
    .B(_00969_),
    .Y(_00970_));
 sg13g2_xnor2_1 _11333_ (.Y(_00971_),
    .A(_00938_),
    .B(_00970_));
 sg13g2_o21ai_1 _11334_ (.B1(_00871_),
    .Y(_00972_),
    .A1(_00870_),
    .A2(_00971_));
 sg13g2_a21oi_1 _11335_ (.A1(_00836_),
    .A2(_00839_),
    .Y(_00973_),
    .B1(_00835_));
 sg13g2_nor2_1 _11336_ (.A(_00840_),
    .B(_00973_),
    .Y(_00974_));
 sg13g2_nand2_1 _11337_ (.Y(_00975_),
    .A(_00845_),
    .B(_00853_));
 sg13g2_nand2b_1 _11338_ (.Y(_00976_),
    .B(_00784_),
    .A_N(_00778_));
 sg13g2_a22oi_1 _11339_ (.Y(_00977_),
    .B1(_00976_),
    .B2(_00783_),
    .A2(_00975_),
    .A1(_00852_));
 sg13g2_nand4_1 _11340_ (.B(_00852_),
    .C(_00975_),
    .A(_00783_),
    .Y(_00978_),
    .D(_00976_));
 sg13g2_nor2b_1 _11341_ (.A(_00977_),
    .B_N(_00978_),
    .Y(_00979_));
 sg13g2_xnor2_1 _11342_ (.Y(_00980_),
    .A(_00974_),
    .B(_00979_));
 sg13g2_o21ai_1 _11343_ (.B1(_00771_),
    .Y(_00981_),
    .A1(_00764_),
    .A2(_00772_));
 sg13g2_nand2_1 _11344_ (.Y(_00982_),
    .A(_00754_),
    .B(_00759_));
 sg13g2_nand2b_1 _11345_ (.Y(_00983_),
    .B(_00825_),
    .A_N(_00818_));
 sg13g2_nand2_1 _11346_ (.Y(_00984_),
    .A(_00824_),
    .B(_00983_));
 sg13g2_a21oi_1 _11347_ (.A1(_00758_),
    .A2(_00982_),
    .Y(_00985_),
    .B1(_00984_));
 sg13g2_and3_1 _11348_ (.X(_00986_),
    .A(_00758_),
    .B(_00982_),
    .C(_00984_));
 sg13g2_nor2_1 _11349_ (.A(_00985_),
    .B(_00986_),
    .Y(_00987_));
 sg13g2_nor2_1 _11350_ (.A(_00981_),
    .B(_00985_),
    .Y(_00988_));
 sg13g2_nor2_2 _11351_ (.A(_00986_),
    .B(_00988_),
    .Y(_00989_));
 sg13g2_xor2_1 _11352_ (.B(_00987_),
    .A(_00981_),
    .X(_00990_));
 sg13g2_inv_1 _11353_ (.Y(_00991_),
    .A(_00990_));
 sg13g2_nand2b_1 _11354_ (.Y(_00992_),
    .B(_00990_),
    .A_N(_00980_));
 sg13g2_nand2_1 _11355_ (.Y(_00993_),
    .A(_00980_),
    .B(_00991_));
 sg13g2_nand2_1 _11356_ (.Y(_00994_),
    .A(_00992_),
    .B(_00993_));
 sg13g2_a21oi_1 _11357_ (.A1(_00711_),
    .A2(_00716_),
    .Y(_00995_),
    .B1(_00715_));
 sg13g2_nand2_1 _11358_ (.Y(_00996_),
    .A(_00858_),
    .B(_00864_));
 sg13g2_nand3_1 _11359_ (.B(_00863_),
    .C(_00996_),
    .A(_00730_),
    .Y(_00997_));
 sg13g2_a21oi_1 _11360_ (.A1(_00863_),
    .A2(_00996_),
    .Y(_00998_),
    .B1(_00730_));
 sg13g2_o21ai_1 _11361_ (.B1(_00997_),
    .Y(_00999_),
    .A1(_00995_),
    .A2(_00998_));
 sg13g2_a21o_1 _11362_ (.A2(_00998_),
    .A1(_00995_),
    .B1(_00999_),
    .X(_01000_));
 sg13g2_o21ai_1 _11363_ (.B1(_01000_),
    .Y(_01001_),
    .A1(_00995_),
    .A2(_00997_));
 sg13g2_xnor2_1 _11364_ (.Y(_01002_),
    .A(_00994_),
    .B(_01001_));
 sg13g2_nand2b_1 _11365_ (.Y(_01003_),
    .B(_00733_),
    .A_N(_00739_));
 sg13g2_nand2_2 _11366_ (.Y(_01004_),
    .A(_00740_),
    .B(_01003_));
 sg13g2_o21ai_1 _11367_ (.B1(_00688_),
    .Y(_01005_),
    .A1(_00690_),
    .A2(_00693_));
 sg13g2_nand2_1 _11368_ (.Y(_01006_),
    .A(_00694_),
    .B(_01005_));
 sg13g2_or2_1 _11369_ (.X(_01007_),
    .B(_01006_),
    .A(_01004_));
 sg13g2_and2_1 _11370_ (.A(_01004_),
    .B(_01006_),
    .X(_01008_));
 sg13g2_xor2_1 _11371_ (.B(_01006_),
    .A(_01004_),
    .X(_01009_));
 sg13g2_nand2_2 _11372_ (.Y(_01010_),
    .A(_00684_),
    .B(_00686_));
 sg13g2_xnor2_1 _11373_ (.Y(_01011_),
    .A(_01009_),
    .B(_01010_));
 sg13g2_o21ai_1 _11374_ (.B1(_00703_),
    .Y(_01012_),
    .A1(_00698_),
    .A2(_00704_));
 sg13g2_a21oi_1 _11375_ (.A1(_00650_),
    .A2(_00652_),
    .Y(_01013_),
    .B1(_01012_));
 sg13g2_nand3_1 _11376_ (.B(_00652_),
    .C(_01012_),
    .A(_00650_),
    .Y(_01014_));
 sg13g2_nand2b_1 _11377_ (.Y(_01015_),
    .B(_01014_),
    .A_N(_01013_));
 sg13g2_o21ai_1 _11378_ (.B1(_00660_),
    .Y(_01016_),
    .A1(_00655_),
    .A2(_00661_));
 sg13g2_xnor2_1 _11379_ (.Y(_01017_),
    .A(_01015_),
    .B(_01016_));
 sg13g2_nand2_1 _11380_ (.Y(_01018_),
    .A(_01011_),
    .B(_01017_));
 sg13g2_or2_1 _11381_ (.X(_01019_),
    .B(_01017_),
    .A(_01011_));
 sg13g2_inv_1 _11382_ (.Y(_01020_),
    .A(_01019_));
 sg13g2_nand2_1 _11383_ (.Y(_01021_),
    .A(_01018_),
    .B(_01019_));
 sg13g2_and2_1 _11384_ (.A(_00668_),
    .B(_00675_),
    .X(_01022_));
 sg13g2_o21ai_1 _11385_ (.B1(_00889_),
    .Y(_01023_),
    .A1(_00885_),
    .A2(_00890_));
 sg13g2_o21ai_1 _11386_ (.B1(_01023_),
    .Y(_01024_),
    .A1(_00674_),
    .A2(_01022_));
 sg13g2_or3_1 _11387_ (.A(_00674_),
    .B(_01022_),
    .C(_01023_),
    .X(_01025_));
 sg13g2_nand2_1 _11388_ (.Y(_01026_),
    .A(_01024_),
    .B(_01025_));
 sg13g2_a21oi_2 _11389_ (.B1(_00880_),
    .Y(_01027_),
    .A2(_00881_),
    .A1(_00873_));
 sg13g2_xor2_1 _11390_ (.B(_01027_),
    .A(_01026_),
    .X(_01028_));
 sg13g2_xor2_1 _11391_ (.B(_01028_),
    .A(_01021_),
    .X(_01029_));
 sg13g2_or2_1 _11392_ (.X(_01030_),
    .B(_01029_),
    .A(_01002_));
 sg13g2_nand2_1 _11393_ (.Y(_01031_),
    .A(_01002_),
    .B(_01029_));
 sg13g2_a21oi_2 _11394_ (.B1(_00930_),
    .Y(_01032_),
    .A2(_00931_),
    .A1(_00926_));
 sg13g2_a21o_1 _11395_ (.A2(_00946_),
    .A1(_00943_),
    .B1(_00941_),
    .X(_01033_));
 sg13g2_o21ai_1 _11396_ (.B1(_01033_),
    .Y(_01034_),
    .A1(_00943_),
    .A2(_00946_));
 sg13g2_nor2_1 _11397_ (.A(_01032_),
    .B(_01034_),
    .Y(_01035_));
 sg13g2_and2_1 _11398_ (.A(_01032_),
    .B(_01034_),
    .X(_01036_));
 sg13g2_nor2_1 _11399_ (.A(_01035_),
    .B(_01036_),
    .Y(_01037_));
 sg13g2_o21ai_1 _11400_ (.B1(_00949_),
    .Y(_01038_),
    .A1(_00953_),
    .A2(_00955_));
 sg13g2_nand2_2 _11401_ (.Y(_01039_),
    .A(_00956_),
    .B(_01038_));
 sg13g2_xnor2_1 _11402_ (.Y(_01040_),
    .A(_01037_),
    .B(_01039_));
 sg13g2_a21oi_2 _11403_ (.B1(_00901_),
    .Y(_01041_),
    .A2(_00902_),
    .A1(_00895_));
 sg13g2_a21oi_2 _11404_ (.B1(_00912_),
    .Y(_01042_),
    .A2(_00913_),
    .A1(_00909_));
 sg13g2_nor2b_1 _11405_ (.A(_01042_),
    .B_N(_01041_),
    .Y(_01043_));
 sg13g2_nand2b_1 _11406_ (.Y(_01044_),
    .B(_01042_),
    .A_N(_01041_));
 sg13g2_nand2b_1 _11407_ (.Y(_01045_),
    .B(_01044_),
    .A_N(_01043_));
 sg13g2_a21oi_1 _11408_ (.A1(_00916_),
    .A2(_00922_),
    .Y(_01046_),
    .B1(_00921_));
 sg13g2_xnor2_1 _11409_ (.Y(_01047_),
    .A(_01045_),
    .B(_01046_));
 sg13g2_nand2_1 _11410_ (.Y(_01048_),
    .A(_01040_),
    .B(_01047_));
 sg13g2_nor2_1 _11411_ (.A(_01040_),
    .B(_01047_),
    .Y(_01049_));
 sg13g2_xor2_1 _11412_ (.B(_01047_),
    .A(_01040_),
    .X(_01050_));
 sg13g2_nor2b_1 _11413_ (.A(net2253),
    .B_N(net2618),
    .Y(_01051_));
 sg13g2_nor2_1 _11414_ (.A(net2381),
    .B(net2388),
    .Y(_01052_));
 sg13g2_xor2_1 _11415_ (.B(net2194),
    .A(net2295),
    .X(_01053_));
 sg13g2_nor3_1 _11416_ (.A(_01051_),
    .B(_01052_),
    .C(_01053_),
    .Y(_01054_));
 sg13g2_o21ai_1 _11417_ (.B1(_01053_),
    .Y(_01055_),
    .A1(_01051_),
    .A2(_01052_));
 sg13g2_xnor2_1 _11418_ (.Y(_01056_),
    .A(net2207),
    .B(\net.in[223] ));
 sg13g2_o21ai_1 _11419_ (.B1(_01055_),
    .Y(_01057_),
    .A1(_01054_),
    .A2(_01056_));
 sg13g2_a21oi_1 _11420_ (.A1(_00963_),
    .A2(_00965_),
    .Y(_01058_),
    .B1(_00962_));
 sg13g2_nor2_2 _11421_ (.A(_00966_),
    .B(_01058_),
    .Y(_01059_));
 sg13g2_nor2_1 _11422_ (.A(_01057_),
    .B(_01059_),
    .Y(_01060_));
 sg13g2_xnor2_1 _11423_ (.Y(_01061_),
    .A(_01057_),
    .B(_01059_));
 sg13g2_xnor2_1 _11424_ (.Y(_01062_),
    .A(net2487),
    .B(net2481));
 sg13g2_nand2b_1 _11425_ (.Y(_01063_),
    .B(net2603),
    .A_N(net2517));
 sg13g2_xnor2_1 _11426_ (.Y(_01064_),
    .A(net2513),
    .B(net2463));
 sg13g2_and3_1 _11427_ (.X(_01065_),
    .A(_01062_),
    .B(_01063_),
    .C(_01064_));
 sg13g2_inv_1 _11428_ (.Y(_01066_),
    .A(_01065_));
 sg13g2_a21oi_1 _11429_ (.A1(_01062_),
    .A2(_01063_),
    .Y(_01067_),
    .B1(_01064_));
 sg13g2_xor2_1 _11430_ (.B(net2341),
    .A(net2226),
    .X(_01068_));
 sg13g2_xor2_1 _11431_ (.B(net2442),
    .A(\net.in[145] ),
    .X(_01069_));
 sg13g2_nor2_2 _11432_ (.A(_01068_),
    .B(_01069_),
    .Y(_01070_));
 sg13g2_a21oi_2 _11433_ (.B1(_01067_),
    .Y(_01071_),
    .A2(_01070_),
    .A1(_01066_));
 sg13g2_a21oi_1 _11434_ (.A1(_01057_),
    .A2(_01059_),
    .Y(_01072_),
    .B1(_01071_));
 sg13g2_xnor2_1 _11435_ (.Y(_01073_),
    .A(_01061_),
    .B(_01071_));
 sg13g2_xnor2_1 _11436_ (.Y(_01074_),
    .A(_01050_),
    .B(_01073_));
 sg13g2_nand2_1 _11437_ (.Y(_01075_),
    .A(_01030_),
    .B(_01074_));
 sg13g2_xnor2_1 _11438_ (.Y(_01076_),
    .A(_00948_),
    .B(_00958_));
 sg13g2_xnor2_1 _11439_ (.Y(_01077_),
    .A(_00968_),
    .B(_01076_));
 sg13g2_nor2b_1 _11440_ (.A(_01054_),
    .B_N(_01055_),
    .Y(_01078_));
 sg13g2_xor2_1 _11441_ (.B(_01078_),
    .A(_01056_),
    .X(_01079_));
 sg13g2_nor2_1 _11442_ (.A(_01065_),
    .B(_01067_),
    .Y(_01080_));
 sg13g2_xnor2_1 _11443_ (.Y(_01081_),
    .A(_01070_),
    .B(_01080_));
 sg13g2_inv_1 _11444_ (.Y(_01082_),
    .A(_01081_));
 sg13g2_nand2_1 _11445_ (.Y(_01083_),
    .A(_01079_),
    .B(_01082_));
 sg13g2_xor2_1 _11446_ (.B(_01081_),
    .A(_01079_),
    .X(_01084_));
 sg13g2_nor2_1 _11447_ (.A(net2332),
    .B(net2776),
    .Y(_01085_));
 sg13g2_xnor2_1 _11448_ (.Y(_01086_),
    .A(net2214),
    .B(_01085_));
 sg13g2_xor2_1 _11449_ (.B(net2656),
    .A(net2530),
    .X(_01087_));
 sg13g2_nand2_1 _11450_ (.Y(_01088_),
    .A(net2422),
    .B(_06045_));
 sg13g2_nor2_1 _11451_ (.A(net2359),
    .B(net2634),
    .Y(_01089_));
 sg13g2_xnor2_1 _11452_ (.Y(_01090_),
    .A(_01088_),
    .B(_01089_));
 sg13g2_nand2_1 _11453_ (.Y(_01091_),
    .A(_01087_),
    .B(_01090_));
 sg13g2_xor2_1 _11454_ (.B(_01090_),
    .A(_01087_),
    .X(_01092_));
 sg13g2_xnor2_1 _11455_ (.Y(_01093_),
    .A(_01086_),
    .B(_01092_));
 sg13g2_xnor2_1 _11456_ (.Y(_01094_),
    .A(_01084_),
    .B(_01093_));
 sg13g2_nor2_1 _11457_ (.A(_01077_),
    .B(_01094_),
    .Y(_01095_));
 sg13g2_and2_1 _11458_ (.A(_01077_),
    .B(_01094_),
    .X(_01096_));
 sg13g2_nor2_1 _11459_ (.A(_01095_),
    .B(_01096_),
    .Y(_01097_));
 sg13g2_xor2_1 _11460_ (.B(net2403),
    .A(net2482),
    .X(_01098_));
 sg13g2_a21oi_2 _11461_ (.B1(_00776_),
    .Y(_01099_),
    .A2(_01098_),
    .A1(net2525));
 sg13g2_xnor2_1 _11462_ (.Y(_01100_),
    .A(net2614),
    .B(net2362));
 sg13g2_xnor2_1 _11463_ (.Y(_01101_),
    .A(net2629),
    .B(_01100_));
 sg13g2_nor2_1 _11464_ (.A(net2407),
    .B(net2209),
    .Y(_01102_));
 sg13g2_xor2_1 _11465_ (.B(\net.in[209] ),
    .A(net2359),
    .X(_01103_));
 sg13g2_xnor2_1 _11466_ (.Y(_01104_),
    .A(_01102_),
    .B(_01103_));
 sg13g2_nor2_1 _11467_ (.A(_01101_),
    .B(_01104_),
    .Y(_01105_));
 sg13g2_nand2_1 _11468_ (.Y(_01106_),
    .A(_01101_),
    .B(_01104_));
 sg13g2_nor2b_1 _11469_ (.A(_01105_),
    .B_N(_01106_),
    .Y(_01107_));
 sg13g2_xnor2_1 _11470_ (.Y(_01108_),
    .A(_01099_),
    .B(_01107_));
 sg13g2_a21oi_1 _11471_ (.A1(net2555),
    .A2(_05572_),
    .Y(_01109_),
    .B1(net2550));
 sg13g2_a21oi_1 _11472_ (.A1(_05176_),
    .A2(net2654),
    .Y(_01110_),
    .B1(net2518));
 sg13g2_nand2_2 _11473_ (.Y(_01111_),
    .A(_01109_),
    .B(_01110_));
 sg13g2_nand2_1 _11474_ (.Y(_01112_),
    .A(net2389),
    .B(net2397));
 sg13g2_xnor2_1 _11475_ (.Y(_01113_),
    .A(net2398),
    .B(net2341));
 sg13g2_nand2_2 _11476_ (.Y(_01114_),
    .A(net2180),
    .B(_01113_));
 sg13g2_nand3_1 _11477_ (.B(_01112_),
    .C(_01114_),
    .A(_01111_),
    .Y(_01115_));
 sg13g2_a21o_1 _11478_ (.A2(_01114_),
    .A1(_01112_),
    .B1(_01111_),
    .X(_01116_));
 sg13g2_nand2_1 _11479_ (.Y(_01117_),
    .A(_01115_),
    .B(_01116_));
 sg13g2_xnor2_1 _11480_ (.Y(_01118_),
    .A(net2304),
    .B(net2214));
 sg13g2_xnor2_1 _11481_ (.Y(_01119_),
    .A(_01117_),
    .B(_01118_));
 sg13g2_or2_1 _11482_ (.X(_01120_),
    .B(_01119_),
    .A(_01108_));
 sg13g2_xnor2_1 _11483_ (.Y(_01121_),
    .A(_01108_),
    .B(_01119_));
 sg13g2_nor2_1 _11484_ (.A(net2389),
    .B(net2381),
    .Y(_01122_));
 sg13g2_nor2b_1 _11485_ (.A(net2354),
    .B_N(net2426),
    .Y(_01123_));
 sg13g2_xnor2_1 _11486_ (.Y(_01124_),
    .A(net2434),
    .B(_01123_));
 sg13g2_nor3_1 _11487_ (.A(_00421_),
    .B(_01122_),
    .C(_01124_),
    .Y(_01125_));
 sg13g2_o21ai_1 _11488_ (.B1(_01124_),
    .Y(_01126_),
    .A1(_00421_),
    .A2(_01122_));
 sg13g2_nor2b_1 _11489_ (.A(_01125_),
    .B_N(_01126_),
    .Y(_01127_));
 sg13g2_xnor2_1 _11490_ (.Y(_01128_),
    .A(net2539),
    .B(net2553));
 sg13g2_xor2_1 _11491_ (.B(_01128_),
    .A(_01127_),
    .X(_01129_));
 sg13g2_xnor2_1 _11492_ (.Y(_01130_),
    .A(_01121_),
    .B(_01129_));
 sg13g2_nor2_1 _11493_ (.A(_01095_),
    .B(_01130_),
    .Y(_01131_));
 sg13g2_nor2_2 _11494_ (.A(_01096_),
    .B(_01131_),
    .Y(_01132_));
 sg13g2_xor2_1 _11495_ (.B(_01130_),
    .A(_01097_),
    .X(_01133_));
 sg13g2_xor2_1 _11496_ (.B(\net.in[223] ),
    .A(net2211),
    .X(_01134_));
 sg13g2_xor2_1 _11497_ (.B(net2686),
    .A(net2259),
    .X(_01135_));
 sg13g2_nor2_2 _11498_ (.A(_01134_),
    .B(_01135_),
    .Y(_01136_));
 sg13g2_nor2_1 _11499_ (.A(net2799),
    .B(net2237),
    .Y(_01137_));
 sg13g2_xnor2_1 _11500_ (.Y(_01138_),
    .A(_00843_),
    .B(_01137_));
 sg13g2_nor2b_1 _11501_ (.A(net2370),
    .B_N(net2762),
    .Y(_01139_));
 sg13g2_xnor2_1 _11502_ (.Y(_01140_),
    .A(net2460),
    .B(net2816));
 sg13g2_xnor2_1 _11503_ (.Y(_01141_),
    .A(_01139_),
    .B(_01140_));
 sg13g2_nor2_1 _11504_ (.A(_01138_),
    .B(_01141_),
    .Y(_01142_));
 sg13g2_nand2_1 _11505_ (.Y(_01143_),
    .A(_01138_),
    .B(_01141_));
 sg13g2_nor2b_1 _11506_ (.A(_01142_),
    .B_N(_01143_),
    .Y(_01144_));
 sg13g2_nor2_2 _11507_ (.A(net2298),
    .B(net2302),
    .Y(_01145_));
 sg13g2_nor2_1 _11508_ (.A(net2191),
    .B(\net.in[247] ),
    .Y(_01146_));
 sg13g2_xnor2_1 _11509_ (.Y(_01147_),
    .A(_01145_),
    .B(_01146_));
 sg13g2_xnor2_1 _11510_ (.Y(_01148_),
    .A(_01144_),
    .B(_01147_));
 sg13g2_xor2_1 _11511_ (.B(net2634),
    .A(net2581),
    .X(_01149_));
 sg13g2_nor2_1 _11512_ (.A(net2345),
    .B(net2212),
    .Y(_01150_));
 sg13g2_xnor2_1 _11513_ (.Y(_01151_),
    .A(net2291),
    .B(net2248));
 sg13g2_xnor2_1 _11514_ (.Y(_01152_),
    .A(_01150_),
    .B(_01151_));
 sg13g2_nand2_1 _11515_ (.Y(_01153_),
    .A(_01149_),
    .B(_01152_));
 sg13g2_xnor2_1 _11516_ (.Y(_01154_),
    .A(_01149_),
    .B(_01152_));
 sg13g2_xnor2_1 _11517_ (.Y(_01155_),
    .A(\net.in[229] ),
    .B(net2395));
 sg13g2_nand2_1 _11518_ (.Y(_01156_),
    .A(net2230),
    .B(net2803));
 sg13g2_o21ai_1 _11519_ (.B1(_01156_),
    .Y(_01157_),
    .A1(net2803),
    .A2(_01155_));
 sg13g2_nand2_1 _11520_ (.Y(_01158_),
    .A(_01153_),
    .B(_01157_));
 sg13g2_o21ai_1 _11521_ (.B1(_01158_),
    .Y(_01159_),
    .A1(_01149_),
    .A2(_01152_));
 sg13g2_xnor2_1 _11522_ (.Y(_01160_),
    .A(_01154_),
    .B(_01157_));
 sg13g2_nand2b_1 _11523_ (.Y(_01161_),
    .B(net2517),
    .A_N(net2281));
 sg13g2_xnor2_1 _11524_ (.Y(_01162_),
    .A(net2623),
    .B(net2287));
 sg13g2_xnor2_1 _11525_ (.Y(_01163_),
    .A(_01161_),
    .B(_01162_));
 sg13g2_nor2_1 _11526_ (.A(net2752),
    .B(net2354),
    .Y(_01164_));
 sg13g2_nor2_1 _11527_ (.A(net2686),
    .B(net2407),
    .Y(_01165_));
 sg13g2_xnor2_1 _11528_ (.Y(_01166_),
    .A(_01164_),
    .B(_01165_));
 sg13g2_inv_1 _11529_ (.Y(_01167_),
    .A(_01166_));
 sg13g2_nor2_1 _11530_ (.A(_01163_),
    .B(_01167_),
    .Y(_01168_));
 sg13g2_xnor2_1 _11531_ (.Y(_01169_),
    .A(_01163_),
    .B(_01166_));
 sg13g2_xor2_1 _11532_ (.B(net2255),
    .A(net2226),
    .X(_01170_));
 sg13g2_xnor2_1 _11533_ (.Y(_01171_),
    .A(_01169_),
    .B(_01170_));
 sg13g2_or2_1 _11534_ (.X(_01172_),
    .B(_01171_),
    .A(_01160_));
 sg13g2_xnor2_1 _11535_ (.Y(_01173_),
    .A(_01160_),
    .B(_01171_));
 sg13g2_xnor2_1 _11536_ (.Y(_01174_),
    .A(_01148_),
    .B(_01173_));
 sg13g2_a21oi_1 _11537_ (.A1(net2430),
    .A2(_05418_),
    .Y(_01175_),
    .B1(net2357));
 sg13g2_a21oi_1 _11538_ (.A1(_05022_),
    .A2(net2437),
    .Y(_01176_),
    .B1(net2381));
 sg13g2_nand2_2 _11539_ (.Y(_01177_),
    .A(_01175_),
    .B(_01176_));
 sg13g2_and2_1 _11540_ (.A(net2367),
    .B(net2209),
    .X(_01178_));
 sg13g2_nor2_1 _11541_ (.A(net2367),
    .B(net2209),
    .Y(_01179_));
 sg13g2_nor2_1 _11542_ (.A(net2325),
    .B(net2586),
    .Y(_01180_));
 sg13g2_nor3_2 _11543_ (.A(_01178_),
    .B(_01179_),
    .C(_01180_),
    .Y(_01181_));
 sg13g2_nor2_1 _11544_ (.A(net2448),
    .B(net2488),
    .Y(_01182_));
 sg13g2_xnor2_1 _11545_ (.Y(_01183_),
    .A(net2276),
    .B(_01182_));
 sg13g2_nand2_1 _11546_ (.Y(_01184_),
    .A(_01181_),
    .B(_01183_));
 sg13g2_nor2_1 _11547_ (.A(_01181_),
    .B(_01183_),
    .Y(_01185_));
 sg13g2_a21oi_2 _11548_ (.B1(_01185_),
    .Y(_01186_),
    .A2(_01184_),
    .A1(_01177_));
 sg13g2_xor2_1 _11549_ (.B(_01183_),
    .A(_01181_),
    .X(_01187_));
 sg13g2_xnor2_1 _11550_ (.Y(_01188_),
    .A(_01177_),
    .B(_01187_));
 sg13g2_xnor2_1 _11551_ (.Y(_01189_),
    .A(net2792),
    .B(net2562));
 sg13g2_nor2_1 _11552_ (.A(net2525),
    .B(net2586),
    .Y(_01190_));
 sg13g2_xnor2_1 _11553_ (.Y(_01191_),
    .A(_07585_),
    .B(_01190_));
 sg13g2_inv_1 _11554_ (.Y(_01192_),
    .A(_01191_));
 sg13g2_nand2b_1 _11555_ (.Y(_01193_),
    .B(_01191_),
    .A_N(_01189_));
 sg13g2_xnor2_1 _11556_ (.Y(_01194_),
    .A(_01189_),
    .B(_01191_));
 sg13g2_xor2_1 _11557_ (.B(net2602),
    .A(net2652),
    .X(_01195_));
 sg13g2_xnor2_1 _11558_ (.Y(_01196_),
    .A(_01194_),
    .B(_01195_));
 sg13g2_nand2_1 _11559_ (.Y(_01197_),
    .A(_01188_),
    .B(_01196_));
 sg13g2_nor2_1 _11560_ (.A(_01188_),
    .B(_01196_),
    .Y(_01198_));
 sg13g2_xor2_1 _11561_ (.B(_01196_),
    .A(_01188_),
    .X(_01199_));
 sg13g2_nor2_2 _11562_ (.A(\net.in[145] ),
    .B(net2404),
    .Y(_01200_));
 sg13g2_o21ai_1 _11563_ (.B1(_01200_),
    .Y(_01201_),
    .A1(net2353),
    .A2(_05737_));
 sg13g2_xor2_1 _11564_ (.B(net2264),
    .A(net2295),
    .X(_01202_));
 sg13g2_xnor2_1 _11565_ (.Y(_01203_),
    .A(net2296),
    .B(net2264));
 sg13g2_nor2_1 _11566_ (.A(net2324),
    .B(_05484_),
    .Y(_01204_));
 sg13g2_xnor2_1 _11567_ (.Y(_01205_),
    .A(net2325),
    .B(net2291));
 sg13g2_nor2_1 _11568_ (.A(_01202_),
    .B(_01205_),
    .Y(_01206_));
 sg13g2_xnor2_1 _11569_ (.Y(_01207_),
    .A(_01203_),
    .B(_01205_));
 sg13g2_xnor2_1 _11570_ (.Y(_01208_),
    .A(_01201_),
    .B(_01207_));
 sg13g2_xnor2_1 _11571_ (.Y(_01209_),
    .A(_01199_),
    .B(_01208_));
 sg13g2_nor2_1 _11572_ (.A(_01174_),
    .B(_01209_),
    .Y(_01210_));
 sg13g2_and2_1 _11573_ (.A(_01174_),
    .B(_01209_),
    .X(_01211_));
 sg13g2_inv_1 _11574_ (.Y(_01212_),
    .A(_01211_));
 sg13g2_nor2_1 _11575_ (.A(_01210_),
    .B(_01211_),
    .Y(_01213_));
 sg13g2_a21oi_2 _11576_ (.B1(_01210_),
    .Y(_01214_),
    .A2(_01212_),
    .A1(_01136_));
 sg13g2_xnor2_1 _11577_ (.Y(_01215_),
    .A(_01136_),
    .B(_01213_));
 sg13g2_nor2_1 _11578_ (.A(_01133_),
    .B(_01215_),
    .Y(_01216_));
 sg13g2_xor2_1 _11579_ (.B(_01215_),
    .A(_01133_),
    .X(_01217_));
 sg13g2_xor2_1 _11580_ (.B(_00731_),
    .A(_00718_),
    .X(_01218_));
 sg13g2_xnor2_1 _11581_ (.Y(_01219_),
    .A(_00742_),
    .B(_01218_));
 sg13g2_xor2_1 _11582_ (.B(_00855_),
    .A(_00842_),
    .X(_01220_));
 sg13g2_xnor2_1 _11583_ (.Y(_01221_),
    .A(_00866_),
    .B(_01220_));
 sg13g2_inv_1 _11584_ (.Y(_01222_),
    .A(_01221_));
 sg13g2_nand2b_1 _11585_ (.Y(_01223_),
    .B(_01221_),
    .A_N(_01219_));
 sg13g2_nand2_1 _11586_ (.Y(_01224_),
    .A(_00697_),
    .B(_00707_));
 sg13g2_xnor2_1 _11587_ (.Y(_01225_),
    .A(_00706_),
    .B(_01224_));
 sg13g2_nand2_1 _11588_ (.Y(_01226_),
    .A(_01219_),
    .B(_01222_));
 sg13g2_nand2_1 _11589_ (.Y(_01227_),
    .A(_01225_),
    .B(_01226_));
 sg13g2_xnor2_1 _11590_ (.Y(_01228_),
    .A(_01219_),
    .B(_01221_));
 sg13g2_xnor2_1 _11591_ (.Y(_01229_),
    .A(_01225_),
    .B(_01228_));
 sg13g2_xor2_1 _11592_ (.B(net2330),
    .A(net2343),
    .X(_01230_));
 sg13g2_nor2_2 _11593_ (.A(net2374),
    .B(_01230_),
    .Y(_01231_));
 sg13g2_a21oi_2 _11594_ (.B1(_01231_),
    .Y(_01232_),
    .A2(_05803_),
    .A1(net2371));
 sg13g2_nor2_1 _11595_ (.A(net2352),
    .B(net2343),
    .Y(_01233_));
 sg13g2_xor2_1 _11596_ (.B(net2344),
    .A(net2352),
    .X(_01234_));
 sg13g2_xnor2_1 _11597_ (.Y(_01235_),
    .A(net2349),
    .B(net2341));
 sg13g2_nand2_1 _11598_ (.Y(_01236_),
    .A(_05066_),
    .B(net2312));
 sg13g2_nor2_1 _11599_ (.A(net2304),
    .B(net2299),
    .Y(_01237_));
 sg13g2_nor2b_1 _11600_ (.A(net2359),
    .B_N(net2430),
    .Y(_01238_));
 sg13g2_xnor2_1 _11601_ (.Y(_01239_),
    .A(_01237_),
    .B(_01238_));
 sg13g2_nand3_1 _11602_ (.B(_01236_),
    .C(_01239_),
    .A(_01235_),
    .Y(_01240_));
 sg13g2_a21o_1 _11603_ (.A2(_01236_),
    .A1(_01235_),
    .B1(_01239_),
    .X(_01241_));
 sg13g2_nand2_1 _11604_ (.Y(_01242_),
    .A(_01240_),
    .B(_01241_));
 sg13g2_xnor2_1 _11605_ (.Y(_01243_),
    .A(_01232_),
    .B(_01242_));
 sg13g2_nand2b_1 _11606_ (.Y(_01244_),
    .B(net2800),
    .A_N(net2345));
 sg13g2_nor2_1 _11607_ (.A(net2448),
    .B(net2814),
    .Y(_01245_));
 sg13g2_xnor2_1 _11608_ (.Y(_01246_),
    .A(_01244_),
    .B(_01245_));
 sg13g2_nor2_1 _11609_ (.A(net2662),
    .B(net2426),
    .Y(_01247_));
 sg13g2_nor2_1 _11610_ (.A(net2814),
    .B(net2315),
    .Y(_01248_));
 sg13g2_xnor2_1 _11611_ (.Y(_01249_),
    .A(_01247_),
    .B(_01248_));
 sg13g2_inv_1 _11612_ (.Y(_01250_),
    .A(_01249_));
 sg13g2_nand2_1 _11613_ (.Y(_01251_),
    .A(_01246_),
    .B(_01250_));
 sg13g2_nor2_1 _11614_ (.A(_01246_),
    .B(_01250_),
    .Y(_01252_));
 sg13g2_xnor2_1 _11615_ (.Y(_01253_),
    .A(_01246_),
    .B(_01249_));
 sg13g2_xor2_1 _11616_ (.B(net2812),
    .A(net2800),
    .X(_01254_));
 sg13g2_xnor2_1 _11617_ (.Y(_01255_),
    .A(_01253_),
    .B(_01254_));
 sg13g2_nor2_2 _11618_ (.A(net2404),
    .B(net2809),
    .Y(_01256_));
 sg13g2_nor2_1 _11619_ (.A(net2187),
    .B(net2700),
    .Y(_01257_));
 sg13g2_nand2b_1 _11620_ (.Y(_01258_),
    .B(net2471),
    .A_N(net2766));
 sg13g2_xnor2_1 _11621_ (.Y(_01259_),
    .A(_01257_),
    .B(_01258_));
 sg13g2_nor2b_1 _11622_ (.A(_01259_),
    .B_N(_01256_),
    .Y(_01260_));
 sg13g2_nand2b_1 _11623_ (.Y(_01261_),
    .B(_01259_),
    .A_N(_01256_));
 sg13g2_xnor2_1 _11624_ (.Y(_01262_),
    .A(_01256_),
    .B(_01259_));
 sg13g2_xnor2_1 _11625_ (.Y(_01263_),
    .A(net2336),
    .B(net2370));
 sg13g2_xnor2_1 _11626_ (.Y(_01264_),
    .A(_01262_),
    .B(_01263_));
 sg13g2_nor2b_1 _11627_ (.A(_01255_),
    .B_N(_01264_),
    .Y(_01265_));
 sg13g2_nand2b_1 _11628_ (.Y(_01266_),
    .B(_01255_),
    .A_N(_01264_));
 sg13g2_xnor2_1 _11629_ (.Y(_01267_),
    .A(_01255_),
    .B(_01264_));
 sg13g2_o21ai_1 _11630_ (.B1(_01266_),
    .Y(_01268_),
    .A1(_01243_),
    .A2(_01265_));
 sg13g2_xnor2_1 _11631_ (.Y(_01269_),
    .A(_01243_),
    .B(_01267_));
 sg13g2_xnor2_1 _11632_ (.Y(_01270_),
    .A(_00800_),
    .B(_00815_));
 sg13g2_xnor2_1 _11633_ (.Y(_01271_),
    .A(_00827_),
    .B(_01270_));
 sg13g2_xor2_1 _11634_ (.B(_01271_),
    .A(_01269_),
    .X(_01272_));
 sg13g2_nand2_1 _11635_ (.Y(_01273_),
    .A(_00775_),
    .B(_00787_));
 sg13g2_xnor2_1 _11636_ (.Y(_01274_),
    .A(_00786_),
    .B(_01273_));
 sg13g2_xnor2_1 _11637_ (.Y(_01275_),
    .A(_01272_),
    .B(_01274_));
 sg13g2_xor2_1 _11638_ (.B(_01275_),
    .A(_01229_),
    .X(_01276_));
 sg13g2_xor2_1 _11639_ (.B(_00663_),
    .A(_00653_),
    .X(_01277_));
 sg13g2_xnor2_1 _11640_ (.Y(_01278_),
    .A(_00677_),
    .B(_01277_));
 sg13g2_xor2_1 _11641_ (.B(_00893_),
    .A(_00883_),
    .X(_01279_));
 sg13g2_xnor2_1 _11642_ (.Y(_01280_),
    .A(_00904_),
    .B(_01279_));
 sg13g2_nor2_1 _11643_ (.A(_01278_),
    .B(_01280_),
    .Y(_01281_));
 sg13g2_nand2_1 _11644_ (.Y(_01282_),
    .A(_01278_),
    .B(_01280_));
 sg13g2_nand2b_1 _11645_ (.Y(_01283_),
    .B(_01282_),
    .A_N(_01281_));
 sg13g2_nand2_1 _11646_ (.Y(_01284_),
    .A(_00925_),
    .B(_00934_));
 sg13g2_xor2_1 _11647_ (.B(_01284_),
    .A(_00933_),
    .X(_01285_));
 sg13g2_xnor2_1 _11648_ (.Y(_01286_),
    .A(_01283_),
    .B(_01285_));
 sg13g2_xnor2_1 _11649_ (.Y(_01287_),
    .A(_01276_),
    .B(_01286_));
 sg13g2_a21oi_2 _11650_ (.B1(_01216_),
    .Y(_01288_),
    .A2(_01287_),
    .A1(_01217_));
 sg13g2_a21o_1 _11651_ (.A2(_01275_),
    .A1(_01229_),
    .B1(_01286_),
    .X(_01289_));
 sg13g2_o21ai_1 _11652_ (.B1(_01289_),
    .Y(_01290_),
    .A1(_01229_),
    .A2(_01275_));
 sg13g2_nor2b_1 _11653_ (.A(_01288_),
    .B_N(_01290_),
    .Y(_01291_));
 sg13g2_xor2_1 _11654_ (.B(_01290_),
    .A(_01288_),
    .X(_01292_));
 sg13g2_a21o_1 _11655_ (.A2(_01271_),
    .A1(_01269_),
    .B1(_01274_),
    .X(_01293_));
 sg13g2_o21ai_1 _11656_ (.B1(_01293_),
    .Y(_01294_),
    .A1(_01269_),
    .A2(_01271_));
 sg13g2_a21oi_1 _11657_ (.A1(_01223_),
    .A2(_01227_),
    .Y(_01295_),
    .B1(_01294_));
 sg13g2_and3_1 _11658_ (.X(_01296_),
    .A(_01223_),
    .B(_01227_),
    .C(_01294_));
 sg13g2_nor2_1 _11659_ (.A(_01295_),
    .B(_01296_),
    .Y(_01297_));
 sg13g2_o21ai_1 _11660_ (.B1(_01282_),
    .Y(_01298_),
    .A1(_01281_),
    .A2(_01285_));
 sg13g2_xnor2_1 _11661_ (.Y(_01299_),
    .A(_01297_),
    .B(_01298_));
 sg13g2_nand2_1 _11662_ (.Y(_01300_),
    .A(_01292_),
    .B(_01299_));
 sg13g2_nor2_1 _11663_ (.A(_01292_),
    .B(_01299_),
    .Y(_01301_));
 sg13g2_nand2_1 _11664_ (.Y(_01302_),
    .A(_01132_),
    .B(_01214_));
 sg13g2_nor2_1 _11665_ (.A(_01132_),
    .B(_01214_),
    .Y(_01303_));
 sg13g2_a21oi_1 _11666_ (.A1(_01268_),
    .A2(_01302_),
    .Y(_01304_),
    .B1(_01303_));
 sg13g2_xnor2_1 _11667_ (.Y(_01305_),
    .A(_01132_),
    .B(_01214_));
 sg13g2_xnor2_1 _11668_ (.Y(_01306_),
    .A(_01268_),
    .B(_01305_));
 sg13g2_a21oi_1 _11669_ (.A1(_01300_),
    .A2(_01306_),
    .Y(_01307_),
    .B1(_01301_));
 sg13g2_a21oi_1 _11670_ (.A1(_01031_),
    .A2(_01075_),
    .Y(_01308_),
    .B1(_01307_));
 sg13g2_nand3_1 _11671_ (.B(_01075_),
    .C(_01307_),
    .A(_01031_),
    .Y(_01309_));
 sg13g2_nand2b_1 _11672_ (.Y(_01310_),
    .B(_01309_),
    .A_N(_01308_));
 sg13g2_a21oi_1 _11673_ (.A1(_00972_),
    .A2(_01309_),
    .Y(_01311_),
    .B1(_01308_));
 sg13g2_xnor2_1 _11674_ (.Y(_01312_),
    .A(_00972_),
    .B(_01310_));
 sg13g2_inv_1 _11675_ (.Y(_01313_),
    .A(_01312_));
 sg13g2_nand2_1 _11676_ (.Y(_01314_),
    .A(_01030_),
    .B(_01031_));
 sg13g2_xor2_1 _11677_ (.B(_01314_),
    .A(_01074_),
    .X(_01315_));
 sg13g2_inv_1 _11678_ (.Y(_01316_),
    .A(_01315_));
 sg13g2_xor2_1 _11679_ (.B(_01299_),
    .A(_01292_),
    .X(_01317_));
 sg13g2_xnor2_1 _11680_ (.Y(_01318_),
    .A(_01306_),
    .B(_01317_));
 sg13g2_nand2b_1 _11681_ (.Y(_01319_),
    .B(_00871_),
    .A_N(_00870_));
 sg13g2_xnor2_1 _11682_ (.Y(_01320_),
    .A(_00971_),
    .B(_01319_));
 sg13g2_nand2_1 _11683_ (.Y(_01321_),
    .A(_01318_),
    .B(_01320_));
 sg13g2_nor2_1 _11684_ (.A(_01318_),
    .B(_01320_),
    .Y(_01322_));
 sg13g2_xnor2_1 _11685_ (.Y(_01323_),
    .A(_01318_),
    .B(_01320_));
 sg13g2_a21o_1 _11686_ (.A2(_01119_),
    .A1(_01108_),
    .B1(_01129_),
    .X(_01324_));
 sg13g2_o21ai_1 _11687_ (.B1(_01093_),
    .Y(_01325_),
    .A1(_01079_),
    .A2(_01082_));
 sg13g2_a22oi_1 _11688_ (.Y(_01326_),
    .B1(_01325_),
    .B2(_01083_),
    .A2(_01324_),
    .A1(_01120_));
 sg13g2_nand4_1 _11689_ (.B(_01120_),
    .C(_01324_),
    .A(_01083_),
    .Y(_01327_),
    .D(_01325_));
 sg13g2_nor2b_1 _11690_ (.A(_01326_),
    .B_N(_01327_),
    .Y(_01328_));
 sg13g2_a21oi_1 _11691_ (.A1(_01197_),
    .A2(_01208_),
    .Y(_01329_),
    .B1(_01198_));
 sg13g2_inv_1 _11692_ (.Y(_01330_),
    .A(_01329_));
 sg13g2_xnor2_1 _11693_ (.Y(_01331_),
    .A(_01328_),
    .B(_01330_));
 sg13g2_or2_1 _11694_ (.X(_01332_),
    .B(_01254_),
    .A(_01252_));
 sg13g2_a21o_1 _11695_ (.A2(_01171_),
    .A1(_01160_),
    .B1(_01148_),
    .X(_01333_));
 sg13g2_a22oi_1 _11696_ (.Y(_01334_),
    .B1(_01333_),
    .B2(_01172_),
    .A2(_01332_),
    .A1(_01251_));
 sg13g2_nand4_1 _11697_ (.B(_01251_),
    .C(_01332_),
    .A(_01172_),
    .Y(_01335_),
    .D(_01333_));
 sg13g2_nand2b_1 _11698_ (.Y(_01336_),
    .B(_01335_),
    .A_N(_01334_));
 sg13g2_a21o_1 _11699_ (.A2(_01263_),
    .A1(_01261_),
    .B1(_01260_),
    .X(_01337_));
 sg13g2_xor2_1 _11700_ (.B(_01337_),
    .A(_01336_),
    .X(_01338_));
 sg13g2_nand2_1 _11701_ (.Y(_01339_),
    .A(_01331_),
    .B(_01338_));
 sg13g2_or2_1 _11702_ (.X(_01340_),
    .B(_01338_),
    .A(_01331_));
 sg13g2_nand2_1 _11703_ (.Y(_01341_),
    .A(_01339_),
    .B(_01340_));
 sg13g2_o21ai_1 _11704_ (.B1(_00810_),
    .Y(_01342_),
    .A1(_00809_),
    .A2(_00814_));
 sg13g2_nand2b_1 _11705_ (.Y(_01343_),
    .B(_01240_),
    .A_N(_01232_));
 sg13g2_or2_1 _11706_ (.X(_01344_),
    .B(_00799_),
    .A(_00796_));
 sg13g2_a22oi_1 _11707_ (.Y(_01345_),
    .B1(_01344_),
    .B2(_00795_),
    .A2(_01343_),
    .A1(_01241_));
 sg13g2_and4_1 _11708_ (.A(_00795_),
    .B(_01241_),
    .C(_01343_),
    .D(_01344_),
    .X(_01346_));
 sg13g2_nor2_1 _11709_ (.A(_01345_),
    .B(_01346_),
    .Y(_01347_));
 sg13g2_xnor2_1 _11710_ (.Y(_01348_),
    .A(_01342_),
    .B(_01347_));
 sg13g2_xnor2_1 _11711_ (.Y(_01349_),
    .A(_01341_),
    .B(_01348_));
 sg13g2_xnor2_1 _11712_ (.Y(_01350_),
    .A(_01323_),
    .B(_01349_));
 sg13g2_nand2_1 _11713_ (.Y(_01351_),
    .A(_01316_),
    .B(_01350_));
 sg13g2_xnor2_1 _11714_ (.Y(_01352_),
    .A(_01316_),
    .B(_01350_));
 sg13g2_nand2b_1 _11715_ (.Y(_01353_),
    .B(_01128_),
    .A_N(_01125_));
 sg13g2_a21o_1 _11716_ (.A2(_01192_),
    .A1(_01189_),
    .B1(_01195_),
    .X(_01354_));
 sg13g2_a22oi_1 _11717_ (.Y(_01355_),
    .B1(_01354_),
    .B2(_01193_),
    .A2(_01353_),
    .A1(_01126_));
 sg13g2_nand4_1 _11718_ (.B(_01193_),
    .C(_01353_),
    .A(_01126_),
    .Y(_01356_),
    .D(_01354_));
 sg13g2_a21oi_2 _11719_ (.B1(_01355_),
    .Y(_01357_),
    .A2(_01356_),
    .A1(_01186_));
 sg13g2_or2_1 _11720_ (.X(_01358_),
    .B(_01356_),
    .A(_01186_));
 sg13g2_a22oi_1 _11721_ (.Y(_01359_),
    .B1(_01357_),
    .B2(_01358_),
    .A2(_01355_),
    .A1(_01186_));
 sg13g2_a21oi_1 _11722_ (.A1(_01099_),
    .A2(_01106_),
    .Y(_01360_),
    .B1(_01105_));
 sg13g2_o21ai_1 _11723_ (.B1(_01086_),
    .Y(_01361_),
    .A1(_01087_),
    .A2(_01090_));
 sg13g2_nand2_1 _11724_ (.Y(_01362_),
    .A(_01115_),
    .B(_01118_));
 sg13g2_a22oi_1 _11725_ (.Y(_01363_),
    .B1(_01362_),
    .B2(_01116_),
    .A2(_01361_),
    .A1(_01091_));
 sg13g2_nand4_1 _11726_ (.B(_01116_),
    .C(_01361_),
    .A(_01091_),
    .Y(_01364_),
    .D(_01362_));
 sg13g2_o21ai_1 _11727_ (.B1(_01364_),
    .Y(_01365_),
    .A1(_01360_),
    .A2(_01363_));
 sg13g2_or2_1 _11728_ (.X(_01366_),
    .B(_01364_),
    .A(_01360_));
 sg13g2_a22oi_1 _11729_ (.Y(_01367_),
    .B1(_01365_),
    .B2(_01366_),
    .A2(_01363_),
    .A1(_01360_));
 sg13g2_nand2_1 _11730_ (.Y(_01368_),
    .A(_01359_),
    .B(_01367_));
 sg13g2_or2_1 _11731_ (.X(_01369_),
    .B(_01367_),
    .A(_01359_));
 sg13g2_nand2_1 _11732_ (.Y(_01370_),
    .A(_01368_),
    .B(_01369_));
 sg13g2_nor2_1 _11733_ (.A(_01201_),
    .B(_01206_),
    .Y(_01371_));
 sg13g2_a21oi_2 _11734_ (.B1(_01371_),
    .Y(_01372_),
    .A2(_01205_),
    .A1(_01202_));
 sg13g2_nor2_1 _11735_ (.A(_01159_),
    .B(_01372_),
    .Y(_01373_));
 sg13g2_nand2_1 _11736_ (.Y(_01374_),
    .A(_01159_),
    .B(_01372_));
 sg13g2_nor2b_1 _11737_ (.A(_01373_),
    .B_N(_01374_),
    .Y(_01375_));
 sg13g2_nor2_1 _11738_ (.A(_01168_),
    .B(_01170_),
    .Y(_01376_));
 sg13g2_a21oi_2 _11739_ (.B1(_01376_),
    .Y(_01377_),
    .A2(_01167_),
    .A1(_01163_));
 sg13g2_xnor2_1 _11740_ (.Y(_01378_),
    .A(_01375_),
    .B(_01377_));
 sg13g2_xor2_1 _11741_ (.B(_01378_),
    .A(_01370_),
    .X(_01379_));
 sg13g2_xnor2_1 _11742_ (.Y(_01380_),
    .A(_01352_),
    .B(_01379_));
 sg13g2_o21ai_1 _11743_ (.B1(_01143_),
    .Y(_01381_),
    .A1(_01142_),
    .A2(_01147_));
 sg13g2_inv_1 _11744_ (.Y(_01382_),
    .A(_01381_));
 sg13g2_o21ai_1 _11745_ (.B1(_01379_),
    .Y(_01383_),
    .A1(_01316_),
    .A2(_01350_));
 sg13g2_nand2_1 _11746_ (.Y(_01384_),
    .A(_01351_),
    .B(_01383_));
 sg13g2_nand3_1 _11747_ (.B(_01382_),
    .C(_01384_),
    .A(_01380_),
    .Y(_01385_));
 sg13g2_a21o_1 _11748_ (.A2(_01382_),
    .A1(_01380_),
    .B1(_01384_),
    .X(_01386_));
 sg13g2_a21oi_1 _11749_ (.A1(_01321_),
    .A2(_01349_),
    .Y(_01387_),
    .B1(_01322_));
 sg13g2_a21o_1 _11750_ (.A2(_01386_),
    .A1(_01385_),
    .B1(_01387_),
    .X(_01388_));
 sg13g2_nand3_1 _11751_ (.B(_01386_),
    .C(_01387_),
    .A(_01385_),
    .Y(_01389_));
 sg13g2_and3_1 _11752_ (.X(_01390_),
    .A(_01313_),
    .B(_01388_),
    .C(_01389_));
 sg13g2_a21oi_1 _11753_ (.A1(_01388_),
    .A2(_01389_),
    .Y(_01391_),
    .B1(_01313_));
 sg13g2_nand2_1 _11754_ (.Y(_01392_),
    .A(_00992_),
    .B(_01001_));
 sg13g2_nand2_1 _11755_ (.Y(_01393_),
    .A(_01339_),
    .B(_01348_));
 sg13g2_a22oi_1 _11756_ (.Y(_01394_),
    .B1(_01393_),
    .B2(_01340_),
    .A2(_01392_),
    .A1(_00993_));
 sg13g2_nand4_1 _11757_ (.B(_01340_),
    .C(_01392_),
    .A(_00993_),
    .Y(_01395_),
    .D(_01393_));
 sg13g2_nor2b_1 _11758_ (.A(_01394_),
    .B_N(_01395_),
    .Y(_01396_));
 sg13g2_a21oi_2 _11759_ (.B1(_01020_),
    .Y(_01397_),
    .A2(_01028_),
    .A1(_01018_));
 sg13g2_xnor2_1 _11760_ (.Y(_01398_),
    .A(_01396_),
    .B(_01397_));
 sg13g2_or3_1 _11761_ (.A(_01390_),
    .B(_01391_),
    .C(_01398_),
    .X(_01399_));
 sg13g2_o21ai_1 _11762_ (.B1(_01398_),
    .Y(_01400_),
    .A1(_01390_),
    .A2(_01391_));
 sg13g2_nor2_1 _11763_ (.A(_01295_),
    .B(_01298_),
    .Y(_01401_));
 sg13g2_o21ai_1 _11764_ (.B1(_01304_),
    .Y(_01402_),
    .A1(_01296_),
    .A2(_01401_));
 sg13g2_nor3_1 _11765_ (.A(_01296_),
    .B(_01304_),
    .C(_01401_),
    .Y(_01403_));
 sg13g2_inv_1 _11766_ (.Y(_01404_),
    .A(_01403_));
 sg13g2_nand2_1 _11767_ (.Y(_01405_),
    .A(_01402_),
    .B(_01404_));
 sg13g2_o21ai_1 _11768_ (.B1(_00832_),
    .Y(_01406_),
    .A1(_00830_),
    .A2(_00868_));
 sg13g2_inv_1 _11769_ (.Y(_01407_),
    .A(_01406_));
 sg13g2_xnor2_1 _11770_ (.Y(_01408_),
    .A(_01405_),
    .B(_01406_));
 sg13g2_nand2_1 _11771_ (.Y(_01409_),
    .A(_01368_),
    .B(_01378_));
 sg13g2_a21oi_1 _11772_ (.A1(_01048_),
    .A2(_01073_),
    .Y(_01410_),
    .B1(_01049_));
 sg13g2_a21oi_2 _11773_ (.B1(_01410_),
    .Y(_01411_),
    .A2(_01409_),
    .A1(_01369_));
 sg13g2_and3_1 _11774_ (.X(_01412_),
    .A(_01369_),
    .B(_01409_),
    .C(_01410_));
 sg13g2_nor2_1 _11775_ (.A(_01411_),
    .B(_01412_),
    .Y(_01413_));
 sg13g2_xnor2_1 _11776_ (.Y(_01414_),
    .A(_01291_),
    .B(_01413_));
 sg13g2_nand2_1 _11777_ (.Y(_01415_),
    .A(_01408_),
    .B(_01414_));
 sg13g2_nor2_1 _11778_ (.A(_01408_),
    .B(_01414_),
    .Y(_01416_));
 sg13g2_xnor2_1 _11779_ (.Y(_01417_),
    .A(_01408_),
    .B(_01414_));
 sg13g2_nor2_1 _11780_ (.A(_00937_),
    .B(_00970_),
    .Y(_01418_));
 sg13g2_nor2_2 _11781_ (.A(_00936_),
    .B(_01418_),
    .Y(_01419_));
 sg13g2_nor2_1 _11782_ (.A(_00748_),
    .B(_01419_),
    .Y(_01420_));
 sg13g2_nand2_1 _11783_ (.Y(_01421_),
    .A(_00748_),
    .B(_01419_));
 sg13g2_nor2b_1 _11784_ (.A(_01420_),
    .B_N(_01421_),
    .Y(_01422_));
 sg13g2_o21ai_1 _11785_ (.B1(_01327_),
    .Y(_01423_),
    .A1(_01326_),
    .A2(_01330_));
 sg13g2_xnor2_1 _11786_ (.Y(_01424_),
    .A(_01422_),
    .B(_01423_));
 sg13g2_xnor2_1 _11787_ (.Y(_01425_),
    .A(_01417_),
    .B(_01424_));
 sg13g2_a21o_1 _11788_ (.A2(_01400_),
    .A1(_01399_),
    .B1(_01425_),
    .X(_01426_));
 sg13g2_nand3_1 _11789_ (.B(_01400_),
    .C(_01425_),
    .A(_01399_),
    .Y(_01427_));
 sg13g2_a21oi_2 _11790_ (.B1(_00977_),
    .Y(_01428_),
    .A2(_00978_),
    .A1(_00974_));
 sg13g2_nand2_1 _11791_ (.Y(_01429_),
    .A(_00999_),
    .B(_01428_));
 sg13g2_or2_1 _11792_ (.X(_01430_),
    .B(_01428_),
    .A(_00999_));
 sg13g2_nand2_1 _11793_ (.Y(_01431_),
    .A(_01429_),
    .B(_01430_));
 sg13g2_o21ai_1 _11794_ (.B1(_01007_),
    .Y(_01432_),
    .A1(_01008_),
    .A2(_01010_));
 sg13g2_xnor2_1 _11795_ (.Y(_01433_),
    .A(_01431_),
    .B(_01432_));
 sg13g2_nor2_1 _11796_ (.A(_01342_),
    .B(_01346_),
    .Y(_01434_));
 sg13g2_nor2_2 _11797_ (.A(_01345_),
    .B(_01434_),
    .Y(_01435_));
 sg13g2_a21oi_2 _11798_ (.B1(_01334_),
    .Y(_01436_),
    .A2(_01337_),
    .A1(_01335_));
 sg13g2_or2_1 _11799_ (.X(_01437_),
    .B(_01436_),
    .A(_01435_));
 sg13g2_nand2_1 _11800_ (.Y(_01438_),
    .A(_01435_),
    .B(_01436_));
 sg13g2_nand2_1 _11801_ (.Y(_01439_),
    .A(_01437_),
    .B(_01438_));
 sg13g2_xor2_1 _11802_ (.B(_01439_),
    .A(_00989_),
    .X(_01440_));
 sg13g2_nand2_1 _11803_ (.Y(_01441_),
    .A(_01433_),
    .B(_01440_));
 sg13g2_or2_1 _11804_ (.X(_01442_),
    .B(_01440_),
    .A(_01433_));
 sg13g2_nand2_1 _11805_ (.Y(_01443_),
    .A(_01441_),
    .B(_01442_));
 sg13g2_nand2_1 _11806_ (.Y(_01444_),
    .A(_01024_),
    .B(_01027_));
 sg13g2_and2_1 _11807_ (.A(_01025_),
    .B(_01444_),
    .X(_01445_));
 sg13g2_a21oi_1 _11808_ (.A1(_01014_),
    .A2(_01016_),
    .Y(_01446_),
    .B1(_01013_));
 sg13g2_nor2_1 _11809_ (.A(_01445_),
    .B(_01446_),
    .Y(_01447_));
 sg13g2_nand2_1 _11810_ (.Y(_01448_),
    .A(_01445_),
    .B(_01446_));
 sg13g2_nor2b_1 _11811_ (.A(_01447_),
    .B_N(_01448_),
    .Y(_01449_));
 sg13g2_a21o_2 _11812_ (.A2(_01046_),
    .A1(_01044_),
    .B1(_01043_),
    .X(_01450_));
 sg13g2_xnor2_1 _11813_ (.Y(_01451_),
    .A(_01449_),
    .B(_01450_));
 sg13g2_xnor2_1 _11814_ (.Y(_01452_),
    .A(_01443_),
    .B(_01451_));
 sg13g2_inv_1 _11815_ (.Y(_01453_),
    .A(_01452_));
 sg13g2_a21oi_1 _11816_ (.A1(_01426_),
    .A2(_01427_),
    .Y(_01454_),
    .B1(_01453_));
 sg13g2_nand3_1 _11817_ (.B(_01427_),
    .C(_01453_),
    .A(_01426_),
    .Y(_01455_));
 sg13g2_nand2b_1 _11818_ (.Y(_01456_),
    .B(_01455_),
    .A_N(_01454_));
 sg13g2_nor2_2 _11819_ (.A(_01060_),
    .B(_01072_),
    .Y(_01457_));
 sg13g2_nor2_1 _11820_ (.A(_01036_),
    .B(_01039_),
    .Y(_01458_));
 sg13g2_nor2_1 _11821_ (.A(_01035_),
    .B(_01458_),
    .Y(_01459_));
 sg13g2_and2_1 _11822_ (.A(_01457_),
    .B(_01459_),
    .X(_01460_));
 sg13g2_nor2_1 _11823_ (.A(_01457_),
    .B(_01459_),
    .Y(_01461_));
 sg13g2_nor2_1 _11824_ (.A(_01460_),
    .B(_01461_),
    .Y(_01462_));
 sg13g2_xnor2_1 _11825_ (.Y(_01463_),
    .A(_01365_),
    .B(_01462_));
 sg13g2_nand2b_1 _11826_ (.Y(_01464_),
    .B(_01463_),
    .A_N(_01357_));
 sg13g2_inv_1 _11827_ (.Y(_01465_),
    .A(_01464_));
 sg13g2_nand2b_1 _11828_ (.Y(_01466_),
    .B(_01357_),
    .A_N(_01463_));
 sg13g2_nand2_1 _11829_ (.Y(_01467_),
    .A(_01464_),
    .B(_01466_));
 sg13g2_a21oi_2 _11830_ (.B1(_01373_),
    .Y(_01468_),
    .A2(_01377_),
    .A1(_01374_));
 sg13g2_xor2_1 _11831_ (.B(_01468_),
    .A(_01467_),
    .X(_01469_));
 sg13g2_nand3b_1 _11832_ (.B(_01455_),
    .C(_01469_),
    .Y(_01470_),
    .A_N(_01454_));
 sg13g2_nand2_1 _11833_ (.Y(_01471_),
    .A(_01427_),
    .B(_01452_));
 sg13g2_nand2_1 _11834_ (.Y(_01472_),
    .A(_01426_),
    .B(_01471_));
 sg13g2_nand2_1 _11835_ (.Y(_01473_),
    .A(_01470_),
    .B(_01472_));
 sg13g2_nor2_1 _11836_ (.A(_01470_),
    .B(_01472_),
    .Y(_01474_));
 sg13g2_nor2b_1 _11837_ (.A(_01391_),
    .B_N(_01398_),
    .Y(_01475_));
 sg13g2_nor2_1 _11838_ (.A(_01390_),
    .B(_01475_),
    .Y(_01476_));
 sg13g2_a21oi_1 _11839_ (.A1(_01473_),
    .A2(_01476_),
    .Y(_01477_),
    .B1(_01474_));
 sg13g2_nand2_1 _11840_ (.Y(_01478_),
    .A(_01441_),
    .B(_01451_));
 sg13g2_or2_1 _11841_ (.X(_01479_),
    .B(_01424_),
    .A(_01416_));
 sg13g2_a22oi_1 _11842_ (.Y(_01480_),
    .B1(_01479_),
    .B2(_01415_),
    .A2(_01478_),
    .A1(_01442_));
 sg13g2_nand4_1 _11843_ (.B(_01442_),
    .C(_01478_),
    .A(_01415_),
    .Y(_01481_),
    .D(_01479_));
 sg13g2_o21ai_1 _11844_ (.B1(_01466_),
    .Y(_01482_),
    .A1(_01465_),
    .A2(_01468_));
 sg13g2_nand2b_1 _11845_ (.Y(_01483_),
    .B(_01482_),
    .A_N(_01480_));
 sg13g2_and3_1 _11846_ (.X(_01484_),
    .A(_01477_),
    .B(_01481_),
    .C(_01483_));
 sg13g2_a21o_1 _11847_ (.A2(_01483_),
    .A1(_01481_),
    .B1(_01477_),
    .X(_01485_));
 sg13g2_nand2b_1 _11848_ (.Y(_01486_),
    .B(_01386_),
    .A_N(_01387_));
 sg13g2_a21oi_1 _11849_ (.A1(_01385_),
    .A2(_01486_),
    .Y(_01487_),
    .B1(_01311_));
 sg13g2_nand3_1 _11850_ (.B(_01385_),
    .C(_01486_),
    .A(_01311_),
    .Y(_01488_));
 sg13g2_a21oi_1 _11851_ (.A1(_01395_),
    .A2(_01397_),
    .Y(_01489_),
    .B1(_01394_));
 sg13g2_inv_1 _11852_ (.Y(_01490_),
    .A(_01489_));
 sg13g2_o21ai_1 _11853_ (.B1(_01488_),
    .Y(_01491_),
    .A1(_01487_),
    .A2(_01490_));
 sg13g2_o21ai_1 _11854_ (.B1(_01485_),
    .Y(_01492_),
    .A1(_01484_),
    .A2(_01491_));
 sg13g2_nor2b_1 _11855_ (.A(_01484_),
    .B_N(_01485_),
    .Y(_01493_));
 sg13g2_xnor2_1 _11856_ (.Y(_01494_),
    .A(_01491_),
    .B(_01493_));
 sg13g2_o21ai_1 _11857_ (.B1(_01421_),
    .Y(_01495_),
    .A1(_01420_),
    .A2(_01423_));
 sg13g2_nor2_1 _11858_ (.A(_01291_),
    .B(_01412_),
    .Y(_01496_));
 sg13g2_a21oi_1 _11859_ (.A1(_01402_),
    .A2(_01407_),
    .Y(_01497_),
    .B1(_01403_));
 sg13g2_nor3_2 _11860_ (.A(_01411_),
    .B(_01496_),
    .C(_01497_),
    .Y(_01498_));
 sg13g2_o21ai_1 _11861_ (.B1(_01497_),
    .Y(_01499_),
    .A1(_01411_),
    .A2(_01496_));
 sg13g2_a21oi_2 _11862_ (.B1(_01498_),
    .Y(_01500_),
    .A2(_01499_),
    .A1(_01495_));
 sg13g2_or2_1 _11863_ (.X(_01501_),
    .B(_01499_),
    .A(_01495_));
 sg13g2_a22oi_1 _11864_ (.Y(_01502_),
    .B1(_01500_),
    .B2(_01501_),
    .A2(_01498_),
    .A1(_01495_));
 sg13g2_a21oi_1 _11865_ (.A1(_01448_),
    .A2(_01450_),
    .Y(_01503_),
    .B1(_01447_));
 sg13g2_nand2b_1 _11866_ (.Y(_01504_),
    .B(_01438_),
    .A_N(_00989_));
 sg13g2_nand2_1 _11867_ (.Y(_01505_),
    .A(_01430_),
    .B(_01432_));
 sg13g2_and4_1 _11868_ (.A(_01429_),
    .B(_01437_),
    .C(_01504_),
    .D(_01505_),
    .X(_01506_));
 sg13g2_a22oi_1 _11869_ (.Y(_01507_),
    .B1(_01505_),
    .B2(_01429_),
    .A2(_01504_),
    .A1(_01437_));
 sg13g2_inv_1 _11870_ (.Y(_01508_),
    .A(_01507_));
 sg13g2_o21ai_1 _11871_ (.B1(_01508_),
    .Y(_01509_),
    .A1(_01503_),
    .A2(_01506_));
 sg13g2_a21o_1 _11872_ (.A2(_01506_),
    .A1(_01503_),
    .B1(_01509_),
    .X(_01510_));
 sg13g2_o21ai_1 _11873_ (.B1(_01510_),
    .Y(_01511_),
    .A1(_01503_),
    .A2(_01508_));
 sg13g2_nand2b_1 _11874_ (.Y(_01512_),
    .B(_01511_),
    .A_N(_01502_));
 sg13g2_nor2b_1 _11875_ (.A(_01511_),
    .B_N(_01502_),
    .Y(_01513_));
 sg13g2_nor2_1 _11876_ (.A(_01365_),
    .B(_01461_),
    .Y(_01514_));
 sg13g2_nor2_2 _11877_ (.A(_01460_),
    .B(_01514_),
    .Y(_01515_));
 sg13g2_inv_1 _11878_ (.Y(_01516_),
    .A(_01515_));
 sg13g2_a21oi_1 _11879_ (.A1(_01512_),
    .A2(_01516_),
    .Y(_01517_),
    .B1(_01513_));
 sg13g2_xor2_1 _11880_ (.B(_01472_),
    .A(_01470_),
    .X(_01518_));
 sg13g2_xnor2_1 _11881_ (.Y(_01519_),
    .A(_01476_),
    .B(_01518_));
 sg13g2_nor2b_1 _11882_ (.A(_01480_),
    .B_N(_01481_),
    .Y(_01520_));
 sg13g2_xnor2_1 _11883_ (.Y(_01521_),
    .A(_01482_),
    .B(_01520_));
 sg13g2_nor2_1 _11884_ (.A(_01519_),
    .B(_01521_),
    .Y(_01522_));
 sg13g2_nand2_1 _11885_ (.Y(_01523_),
    .A(_01519_),
    .B(_01521_));
 sg13g2_nand2b_1 _11886_ (.Y(_01524_),
    .B(_01523_),
    .A_N(_01522_));
 sg13g2_nor2b_1 _11887_ (.A(_01487_),
    .B_N(_01488_),
    .Y(_01525_));
 sg13g2_xnor2_1 _11888_ (.Y(_01526_),
    .A(_01489_),
    .B(_01525_));
 sg13g2_xor2_1 _11889_ (.B(_01526_),
    .A(_01524_),
    .X(_01527_));
 sg13g2_xnor2_1 _11890_ (.Y(_01528_),
    .A(_01502_),
    .B(_01511_));
 sg13g2_xnor2_1 _11891_ (.Y(_01529_),
    .A(_01515_),
    .B(_01528_));
 sg13g2_o21ai_1 _11892_ (.B1(_01523_),
    .Y(_01530_),
    .A1(_01522_),
    .A2(_01526_));
 sg13g2_o21ai_1 _11893_ (.B1(_01530_),
    .Y(_01531_),
    .A1(_01527_),
    .A2(_01529_));
 sg13g2_or3_1 _11894_ (.A(_01527_),
    .B(_01529_),
    .C(_01530_),
    .X(_01532_));
 sg13g2_nand2_1 _11895_ (.Y(_01533_),
    .A(_01531_),
    .B(_01532_));
 sg13g2_xnor2_1 _11896_ (.Y(_01534_),
    .A(_01517_),
    .B(_01533_));
 sg13g2_nor2_1 _11897_ (.A(_01494_),
    .B(_01534_),
    .Y(_01535_));
 sg13g2_nand2_1 _11898_ (.Y(_01536_),
    .A(_01494_),
    .B(_01534_));
 sg13g2_o21ai_1 _11899_ (.B1(_01536_),
    .Y(_01537_),
    .A1(_01500_),
    .A2(_01535_));
 sg13g2_nor2b_1 _11900_ (.A(_01535_),
    .B_N(_01536_),
    .Y(_01538_));
 sg13g2_xnor2_1 _11901_ (.Y(_01539_),
    .A(_01500_),
    .B(_01538_));
 sg13g2_a21o_1 _11902_ (.A2(_01539_),
    .A1(_01509_),
    .B1(_01537_),
    .X(_01540_));
 sg13g2_nand3_1 _11903_ (.B(_01537_),
    .C(_01539_),
    .A(_01509_),
    .Y(_01541_));
 sg13g2_nand2_1 _11904_ (.Y(_01542_),
    .A(_01540_),
    .B(_01541_));
 sg13g2_nand2b_1 _11905_ (.Y(_01543_),
    .B(_01532_),
    .A_N(_01517_));
 sg13g2_nand2_1 _11906_ (.Y(_01544_),
    .A(_01531_),
    .B(_01543_));
 sg13g2_xor2_1 _11907_ (.B(_01544_),
    .A(_01542_),
    .X(_01545_));
 sg13g2_nand2_1 _11908_ (.Y(_01546_),
    .A(_01541_),
    .B(_01544_));
 sg13g2_a22oi_1 _11909_ (.Y(_01547_),
    .B1(_01546_),
    .B2(_01540_),
    .A2(_01545_),
    .A1(_01492_));
 sg13g2_inv_1 _11910_ (.Y(_01548_),
    .A(_01547_));
 sg13g2_a21o_1 _11911_ (.A2(_08124_),
    .A1(_08091_),
    .B1(_08168_),
    .X(_01549_));
 sg13g2_o21ai_1 _11912_ (.B1(_01549_),
    .Y(_01550_),
    .A1(_08091_),
    .A2(_08124_));
 sg13g2_nor2_1 _11913_ (.A(_06573_),
    .B(_06661_),
    .Y(_01551_));
 sg13g2_o21ai_1 _11914_ (.B1(_01550_),
    .Y(_01552_),
    .A1(_06650_),
    .A2(_01551_));
 sg13g2_or3_1 _11915_ (.A(_06650_),
    .B(_01550_),
    .C(_01551_),
    .X(_01553_));
 sg13g2_a21oi_1 _11916_ (.A1(_06716_),
    .A2(_06749_),
    .Y(_01554_),
    .B1(_06760_));
 sg13g2_nand2_1 _11917_ (.Y(_01555_),
    .A(_01552_),
    .B(_01554_));
 sg13g2_and2_1 _11918_ (.A(_01553_),
    .B(_01555_),
    .X(_01556_));
 sg13g2_or2_1 _11919_ (.X(_01557_),
    .B(_07057_),
    .A(_07002_));
 sg13g2_nand2_1 _11920_ (.Y(_01558_),
    .A(_07442_),
    .B(_07508_));
 sg13g2_a22oi_1 _11921_ (.Y(_01559_),
    .B1(_01558_),
    .B2(_07519_),
    .A2(_01557_),
    .A1(_07068_));
 sg13g2_nand4_1 _11922_ (.B(_07519_),
    .C(_01557_),
    .A(_07068_),
    .Y(_01560_),
    .D(_01558_));
 sg13g2_a21o_1 _11923_ (.A2(_07618_),
    .A1(_07574_),
    .B1(_07552_),
    .X(_01561_));
 sg13g2_o21ai_1 _11924_ (.B1(_01561_),
    .Y(_01562_),
    .A1(_07574_),
    .A2(_07618_));
 sg13g2_nand2b_1 _11925_ (.Y(_01563_),
    .B(_01562_),
    .A_N(_01559_));
 sg13g2_a21oi_2 _11926_ (.B1(_00558_),
    .Y(_01564_),
    .A2(_00559_),
    .A1(_00552_));
 sg13g2_nand2_1 _11927_ (.Y(_01565_),
    .A(_07354_),
    .B(_01564_));
 sg13g2_nor2_1 _11928_ (.A(_07354_),
    .B(_01564_),
    .Y(_01566_));
 sg13g2_a21oi_1 _11929_ (.A1(_07189_),
    .A2(_01565_),
    .Y(_01567_),
    .B1(_01566_));
 sg13g2_nand3_1 _11930_ (.B(_01563_),
    .C(_01567_),
    .A(_01560_),
    .Y(_01568_));
 sg13g2_a21o_1 _11931_ (.A2(_01563_),
    .A1(_01560_),
    .B1(_01567_),
    .X(_01569_));
 sg13g2_nand2_1 _11932_ (.Y(_01570_),
    .A(_01568_),
    .B(_01569_));
 sg13g2_nand2_1 _11933_ (.Y(_01571_),
    .A(_07739_),
    .B(_07783_));
 sg13g2_nand2_1 _11934_ (.Y(_01572_),
    .A(_07959_),
    .B(_08003_));
 sg13g2_a22oi_1 _11935_ (.Y(_01573_),
    .B1(_01572_),
    .B2(_07992_),
    .A2(_01571_),
    .A1(_07728_));
 sg13g2_nand4_1 _11936_ (.B(_07992_),
    .C(_01571_),
    .A(_07728_),
    .Y(_01574_),
    .D(_01572_));
 sg13g2_o21ai_1 _11937_ (.B1(_07860_),
    .Y(_01575_),
    .A1(_07882_),
    .A2(_07904_));
 sg13g2_nand2_2 _11938_ (.Y(_01576_),
    .A(_07915_),
    .B(_01575_));
 sg13g2_o21ai_1 _11939_ (.B1(_01574_),
    .Y(_01577_),
    .A1(_01573_),
    .A2(_01576_));
 sg13g2_xnor2_1 _11940_ (.Y(_01578_),
    .A(_01570_),
    .B(_01577_));
 sg13g2_or2_1 _11941_ (.X(_01579_),
    .B(_01578_),
    .A(_01556_));
 sg13g2_nand2_1 _11942_ (.Y(_01580_),
    .A(_01556_),
    .B(_01578_));
 sg13g2_a21o_2 _11943_ (.A2(_06276_),
    .A1(_06221_),
    .B1(_06232_),
    .X(_01581_));
 sg13g2_a21oi_2 _11944_ (.B1(_06881_),
    .Y(_01582_),
    .A2(_06870_),
    .A1(_06815_));
 sg13g2_nand2_1 _11945_ (.Y(_01583_),
    .A(_01581_),
    .B(_01582_));
 sg13g2_nor2_1 _11946_ (.A(_01581_),
    .B(_01582_),
    .Y(_01584_));
 sg13g2_nor2_1 _11947_ (.A(_06298_),
    .B(_06353_),
    .Y(_01585_));
 sg13g2_nor2_2 _11948_ (.A(_06364_),
    .B(_01585_),
    .Y(_01586_));
 sg13g2_a21oi_1 _11949_ (.A1(_01583_),
    .A2(_01586_),
    .Y(_01587_),
    .B1(_01584_));
 sg13g2_nand2_1 _11950_ (.Y(_01588_),
    .A(_01580_),
    .B(_01587_));
 sg13g2_nand2_2 _11951_ (.Y(_01589_),
    .A(_01579_),
    .B(_01588_));
 sg13g2_a21oi_1 _11952_ (.A1(_08223_),
    .A2(_00642_),
    .Y(_01590_),
    .B1(_08212_));
 sg13g2_nand2_1 _11953_ (.Y(_01591_),
    .A(_00523_),
    .B(_00641_));
 sg13g2_nor2_1 _11954_ (.A(_01590_),
    .B(_01591_),
    .Y(_01592_));
 sg13g2_xnor2_1 _11955_ (.Y(_01593_),
    .A(_07354_),
    .B(_01564_));
 sg13g2_xnor2_1 _11956_ (.Y(_01594_),
    .A(_07189_),
    .B(_01593_));
 sg13g2_o21ai_1 _11957_ (.B1(_00545_),
    .Y(_01595_),
    .A1(_00538_),
    .A2(_00546_));
 sg13g2_o21ai_1 _11958_ (.B1(_00632_),
    .Y(_01596_),
    .A1(_00627_),
    .A2(_00633_));
 sg13g2_nand2_1 _11959_ (.Y(_01597_),
    .A(_01595_),
    .B(_01596_));
 sg13g2_xor2_1 _11960_ (.B(_01596_),
    .A(_01595_),
    .X(_01598_));
 sg13g2_xnor2_1 _11961_ (.Y(_01599_),
    .A(_00534_),
    .B(_01598_));
 sg13g2_nor2_1 _11962_ (.A(_01594_),
    .B(_01599_),
    .Y(_01600_));
 sg13g2_nand2_1 _11963_ (.Y(_01601_),
    .A(_01594_),
    .B(_01599_));
 sg13g2_nor2b_1 _11964_ (.A(_01559_),
    .B_N(_01560_),
    .Y(_01602_));
 sg13g2_xnor2_1 _11965_ (.Y(_01603_),
    .A(_01562_),
    .B(_01602_));
 sg13g2_o21ai_1 _11966_ (.B1(_01601_),
    .Y(_01604_),
    .A1(_01600_),
    .A2(_01603_));
 sg13g2_nand2b_1 _11967_ (.Y(_01605_),
    .B(_01574_),
    .A_N(_01573_));
 sg13g2_xor2_1 _11968_ (.B(_01605_),
    .A(_01576_),
    .X(_01606_));
 sg13g2_and2_1 _11969_ (.A(_01552_),
    .B(_01553_),
    .X(_01607_));
 sg13g2_xnor2_1 _11970_ (.Y(_01608_),
    .A(_01554_),
    .B(_01607_));
 sg13g2_nand2_1 _11971_ (.Y(_01609_),
    .A(_01606_),
    .B(_01608_));
 sg13g2_nor2_1 _11972_ (.A(_01606_),
    .B(_01608_),
    .Y(_01610_));
 sg13g2_xor2_1 _11973_ (.B(_01582_),
    .A(_01581_),
    .X(_01611_));
 sg13g2_xnor2_1 _11974_ (.Y(_01612_),
    .A(_01586_),
    .B(_01611_));
 sg13g2_a21oi_1 _11975_ (.A1(_01609_),
    .A2(_01612_),
    .Y(_01613_),
    .B1(_01610_));
 sg13g2_nor2_1 _11976_ (.A(_01604_),
    .B(_01613_),
    .Y(_01614_));
 sg13g2_inv_1 _11977_ (.Y(_01615_),
    .A(_01614_));
 sg13g2_and2_1 _11978_ (.A(_01604_),
    .B(_01613_),
    .X(_01616_));
 sg13g2_nor2_1 _11979_ (.A(_01614_),
    .B(_01616_),
    .Y(_01617_));
 sg13g2_xnor2_1 _11980_ (.Y(_01618_),
    .A(_01592_),
    .B(_01617_));
 sg13g2_nand2_1 _11981_ (.Y(_01619_),
    .A(_00301_),
    .B(_00519_));
 sg13g2_nand2_1 _11982_ (.Y(_01620_),
    .A(_00520_),
    .B(_01619_));
 sg13g2_nand2b_1 _11983_ (.Y(_01621_),
    .B(_01620_),
    .A_N(_09554_));
 sg13g2_nor2b_1 _11984_ (.A(_01620_),
    .B_N(_09554_),
    .Y(_01622_));
 sg13g2_nor2_1 _11985_ (.A(_00562_),
    .B(_00637_),
    .Y(_01623_));
 sg13g2_nor2_1 _11986_ (.A(_00638_),
    .B(_01623_),
    .Y(_01624_));
 sg13g2_a21oi_1 _11987_ (.A1(_01621_),
    .A2(_01624_),
    .Y(_01625_),
    .B1(_01622_));
 sg13g2_nand2b_1 _11988_ (.Y(_01626_),
    .B(_07816_),
    .A_N(_08190_));
 sg13g2_nand2_1 _11989_ (.Y(_01627_),
    .A(_06155_),
    .B(_06936_));
 sg13g2_nand4_1 _11990_ (.B(_07827_),
    .C(_01626_),
    .A(_06925_),
    .Y(_01628_),
    .D(_01627_));
 sg13g2_inv_1 _11991_ (.Y(_01629_),
    .A(_01628_));
 sg13g2_a22oi_1 _11992_ (.Y(_01630_),
    .B1(_01627_),
    .B2(_06925_),
    .A2(_01626_),
    .A1(_07827_));
 sg13g2_o21ai_1 _11993_ (.B1(_09367_),
    .Y(_01631_),
    .A1(_09356_),
    .A2(_09499_));
 sg13g2_a21oi_1 _11994_ (.A1(_01628_),
    .A2(_01631_),
    .Y(_01632_),
    .B1(_01630_));
 sg13g2_and2_1 _11995_ (.A(_01625_),
    .B(_01632_),
    .X(_01633_));
 sg13g2_nor2_1 _11996_ (.A(_01625_),
    .B(_01632_),
    .Y(_01634_));
 sg13g2_nor2_1 _11997_ (.A(_01633_),
    .B(_01634_),
    .Y(_01635_));
 sg13g2_nand3_1 _11998_ (.B(_08927_),
    .C(_09081_),
    .A(_08652_),
    .Y(_01636_));
 sg13g2_inv_1 _11999_ (.Y(_01637_),
    .A(_01636_));
 sg13g2_a21oi_1 _12000_ (.A1(_08927_),
    .A2(_09081_),
    .Y(_01638_),
    .B1(_08652_));
 sg13g2_a21oi_2 _12001_ (.B1(_01638_),
    .Y(_01639_),
    .A2(_01636_),
    .A1(_00517_));
 sg13g2_nor2_1 _12002_ (.A(_01633_),
    .B(_01639_),
    .Y(_01640_));
 sg13g2_nor2_1 _12003_ (.A(_01634_),
    .B(_01640_),
    .Y(_01641_));
 sg13g2_xor2_1 _12004_ (.B(_01639_),
    .A(_01635_),
    .X(_01642_));
 sg13g2_or2_1 _12005_ (.X(_01643_),
    .B(_01642_),
    .A(_01618_));
 sg13g2_nand2_1 _12006_ (.Y(_01644_),
    .A(_01618_),
    .B(_01642_));
 sg13g2_o21ai_1 _12007_ (.B1(_07651_),
    .Y(_01645_),
    .A1(_07662_),
    .A2(_07794_));
 sg13g2_nand2_1 _12008_ (.Y(_01646_),
    .A(_08036_),
    .B(_08179_));
 sg13g2_nand2_1 _12009_ (.Y(_01647_),
    .A(_08047_),
    .B(_01646_));
 sg13g2_nand3_1 _12010_ (.B(_01645_),
    .C(_01646_),
    .A(_08047_),
    .Y(_01648_));
 sg13g2_a21oi_1 _12011_ (.A1(_08047_),
    .A2(_01646_),
    .Y(_01649_),
    .B1(_01645_));
 sg13g2_nor2_1 _12012_ (.A(_06793_),
    .B(_06903_),
    .Y(_01650_));
 sg13g2_a21oi_2 _12013_ (.B1(_01650_),
    .Y(_01651_),
    .A2(_06782_),
    .A1(_06683_));
 sg13g2_inv_1 _12014_ (.Y(_01652_),
    .A(_01651_));
 sg13g2_a21oi_2 _12015_ (.B1(_01649_),
    .Y(_01653_),
    .A2(_01652_),
    .A1(_01648_));
 sg13g2_a21oi_1 _12016_ (.A1(_09774_),
    .A2(_00297_),
    .Y(_01654_),
    .B1(_09785_));
 sg13g2_o21ai_1 _12017_ (.B1(_00464_),
    .Y(_01655_),
    .A1(_00348_),
    .A2(_00405_));
 sg13g2_nand2_1 _12018_ (.Y(_01656_),
    .A(_00411_),
    .B(_01655_));
 sg13g2_nand2_1 _12019_ (.Y(_01657_),
    .A(_01654_),
    .B(_01656_));
 sg13g2_or2_1 _12020_ (.X(_01658_),
    .B(_01656_),
    .A(_01654_));
 sg13g2_nand2_1 _12021_ (.Y(_01659_),
    .A(_00596_),
    .B(_01657_));
 sg13g2_nand2_1 _12022_ (.Y(_01660_),
    .A(_00622_),
    .B(_00635_));
 sg13g2_nand2_1 _12023_ (.Y(_01661_),
    .A(_00549_),
    .B(_00561_));
 sg13g2_nand2_2 _12024_ (.Y(_01662_),
    .A(_00550_),
    .B(_01661_));
 sg13g2_nand3_1 _12025_ (.B(_01660_),
    .C(_01662_),
    .A(_00623_),
    .Y(_01663_));
 sg13g2_a21o_1 _12026_ (.A2(_01660_),
    .A1(_00623_),
    .B1(_01662_),
    .X(_01664_));
 sg13g2_a21oi_2 _12027_ (.B1(_07387_),
    .Y(_01665_),
    .A2(_07398_),
    .A1(_07090_));
 sg13g2_nand2_1 _12028_ (.Y(_01666_),
    .A(_01664_),
    .B(_01665_));
 sg13g2_nand2_1 _12029_ (.Y(_01667_),
    .A(_01663_),
    .B(_01666_));
 sg13g2_a21o_1 _12030_ (.A2(_01659_),
    .A1(_01658_),
    .B1(_01667_),
    .X(_01668_));
 sg13g2_nand3_1 _12031_ (.B(_01659_),
    .C(_01667_),
    .A(_01658_),
    .Y(_01669_));
 sg13g2_inv_1 _12032_ (.Y(_01670_),
    .A(_01669_));
 sg13g2_nand2_1 _12033_ (.Y(_01671_),
    .A(_01668_),
    .B(_01669_));
 sg13g2_xor2_1 _12034_ (.B(_01671_),
    .A(_01653_),
    .X(_01672_));
 sg13g2_nand2_1 _12035_ (.Y(_01673_),
    .A(_01644_),
    .B(_01672_));
 sg13g2_nand2_1 _12036_ (.Y(_01674_),
    .A(_01643_),
    .B(_01673_));
 sg13g2_nand2_1 _12037_ (.Y(_01675_),
    .A(_06397_),
    .B(_06529_));
 sg13g2_o21ai_1 _12038_ (.B1(_09334_),
    .Y(_01676_),
    .A1(_09268_),
    .A2(_09301_));
 sg13g2_nand4_1 _12039_ (.B(_09312_),
    .C(_01675_),
    .A(_06408_),
    .Y(_01677_),
    .D(_01676_));
 sg13g2_inv_1 _12040_ (.Y(_01678_),
    .A(_01677_));
 sg13g2_a22oi_1 _12041_ (.Y(_01679_),
    .B1(_01676_),
    .B2(_09312_),
    .A2(_01675_),
    .A1(_06408_));
 sg13g2_o21ai_1 _12042_ (.B1(_09202_),
    .Y(_01680_),
    .A1(_09114_),
    .A2(_09213_));
 sg13g2_a21oi_1 _12043_ (.A1(_01677_),
    .A2(_01680_),
    .Y(_01681_),
    .B1(_01679_));
 sg13g2_nand2_1 _12044_ (.Y(_01682_),
    .A(_09400_),
    .B(_09477_));
 sg13g2_nand2_1 _12045_ (.Y(_01683_),
    .A(_08828_),
    .B(_08894_));
 sg13g2_o21ai_1 _12046_ (.B1(_01683_),
    .Y(_01684_),
    .A1(_08861_),
    .A2(_08883_));
 sg13g2_and3_2 _12047_ (.X(_01685_),
    .A(_09466_),
    .B(_01682_),
    .C(_01684_));
 sg13g2_a21oi_2 _12048_ (.B1(_01684_),
    .Y(_01686_),
    .A2(_01682_),
    .A1(_09466_));
 sg13g2_o21ai_1 _12049_ (.B1(_08773_),
    .Y(_01687_),
    .A1(_08707_),
    .A2(_08784_));
 sg13g2_nor2_1 _12050_ (.A(_01686_),
    .B(_01687_),
    .Y(_01688_));
 sg13g2_o21ai_1 _12051_ (.B1(_01681_),
    .Y(_01689_),
    .A1(_01685_),
    .A2(_01688_));
 sg13g2_or3_1 _12052_ (.A(_01681_),
    .B(_01685_),
    .C(_01688_),
    .X(_01690_));
 sg13g2_and2_1 _12053_ (.A(_01689_),
    .B(_01690_),
    .X(_01691_));
 sg13g2_a21oi_2 _12054_ (.B1(_08454_),
    .Y(_01692_),
    .A2(_08465_),
    .A1(_08355_));
 sg13g2_and2_1 _12055_ (.A(_09059_),
    .B(_01692_),
    .X(_01693_));
 sg13g2_or2_1 _12056_ (.X(_01694_),
    .B(_01692_),
    .A(_09059_));
 sg13g2_o21ai_1 _12057_ (.B1(_01694_),
    .Y(_01695_),
    .A1(_08608_),
    .A2(_01693_));
 sg13g2_xor2_1 _12058_ (.B(_01695_),
    .A(_01691_),
    .X(_01696_));
 sg13g2_a21o_1 _12059_ (.A2(_08311_),
    .A1(_08245_),
    .B1(_08300_),
    .X(_01697_));
 sg13g2_inv_1 _12060_ (.Y(_01698_),
    .A(_01697_));
 sg13g2_nor2_1 _12061_ (.A(_00512_),
    .B(_01698_),
    .Y(_01699_));
 sg13g2_nand2_1 _12062_ (.Y(_01700_),
    .A(_00512_),
    .B(_01698_));
 sg13g2_a21oi_1 _12063_ (.A1(_00488_),
    .A2(_00492_),
    .Y(_01701_),
    .B1(_00497_));
 sg13g2_nor2_2 _12064_ (.A(_00493_),
    .B(_01701_),
    .Y(_01702_));
 sg13g2_o21ai_1 _12065_ (.B1(_01700_),
    .Y(_01703_),
    .A1(_01699_),
    .A2(_01702_));
 sg13g2_nand2_1 _12066_ (.Y(_01704_),
    .A(_00475_),
    .B(_00481_));
 sg13g2_nand2_2 _12067_ (.Y(_01705_),
    .A(_00480_),
    .B(_01704_));
 sg13g2_nand2_1 _12068_ (.Y(_01706_),
    .A(_00305_),
    .B(_00338_));
 sg13g2_o21ai_1 _12069_ (.B1(_01706_),
    .Y(_01707_),
    .A1(_00320_),
    .A2(_00333_));
 sg13g2_or2_1 _12070_ (.X(_01708_),
    .B(_01707_),
    .A(_01705_));
 sg13g2_and2_1 _12071_ (.A(_01705_),
    .B(_01707_),
    .X(_01709_));
 sg13g2_a21o_2 _12072_ (.A2(_00400_),
    .A1(_00384_),
    .B1(_00378_),
    .X(_01710_));
 sg13g2_a21oi_1 _12073_ (.A1(_01708_),
    .A2(_01710_),
    .Y(_01711_),
    .B1(_01709_));
 sg13g2_nand2_1 _12074_ (.Y(_01712_),
    .A(_01703_),
    .B(_01711_));
 sg13g2_or2_1 _12075_ (.X(_01713_),
    .B(_01711_),
    .A(_01703_));
 sg13g2_and2_1 _12076_ (.A(_01712_),
    .B(_01713_),
    .X(_01714_));
 sg13g2_a21o_1 _12077_ (.A2(_09609_),
    .A1(_06705_),
    .B1(_09642_),
    .X(_01715_));
 sg13g2_nand2b_1 _12078_ (.Y(_01716_),
    .B(_00450_),
    .A_N(_00425_));
 sg13g2_a22oi_1 _12079_ (.Y(_01717_),
    .B1(_01716_),
    .B2(_00454_),
    .A2(_01715_),
    .A1(_09620_));
 sg13g2_nand4_1 _12080_ (.B(_00454_),
    .C(_01715_),
    .A(_09620_),
    .Y(_01718_),
    .D(_01716_));
 sg13g2_nor2b_1 _12081_ (.A(_09741_),
    .B_N(_09675_),
    .Y(_01719_));
 sg13g2_a21oi_2 _12082_ (.B1(_01719_),
    .Y(_01720_),
    .A2(_09730_),
    .A1(_09697_));
 sg13g2_o21ai_1 _12083_ (.B1(_01718_),
    .Y(_01721_),
    .A1(_01717_),
    .A2(_01720_));
 sg13g2_xor2_1 _12084_ (.B(_01721_),
    .A(_01714_),
    .X(_01722_));
 sg13g2_nor2_1 _12085_ (.A(_01696_),
    .B(_01722_),
    .Y(_01723_));
 sg13g2_and2_1 _12086_ (.A(_01696_),
    .B(_01722_),
    .X(_01724_));
 sg13g2_nand2_1 _12087_ (.Y(_01725_),
    .A(_00534_),
    .B(_01597_));
 sg13g2_o21ai_1 _12088_ (.B1(_01725_),
    .Y(_01726_),
    .A1(_01595_),
    .A2(_01596_));
 sg13g2_or2_1 _12089_ (.X(_01727_),
    .B(_00580_),
    .A(_00575_));
 sg13g2_or2_1 _12090_ (.X(_01728_),
    .B(_00287_),
    .A(_09840_));
 sg13g2_a22oi_1 _12091_ (.Y(_01729_),
    .B1(_01728_),
    .B2(_00290_),
    .A2(_01727_),
    .A1(_00579_));
 sg13g2_nand4_1 _12092_ (.B(_00579_),
    .C(_01727_),
    .A(_00290_),
    .Y(_01730_),
    .D(_01728_));
 sg13g2_a21oi_1 _12093_ (.A1(_00585_),
    .A2(_00591_),
    .Y(_01731_),
    .B1(_00590_));
 sg13g2_o21ai_1 _12094_ (.B1(_01730_),
    .Y(_01732_),
    .A1(_01729_),
    .A2(_01731_));
 sg13g2_or2_1 _12095_ (.X(_01733_),
    .B(_00572_),
    .A(_00568_));
 sg13g2_a21oi_1 _12096_ (.A1(_00569_),
    .A2(_01733_),
    .Y(_01734_),
    .B1(_00620_));
 sg13g2_and3_1 _12097_ (.X(_01735_),
    .A(_00569_),
    .B(_00620_),
    .C(_01733_));
 sg13g2_a21o_1 _12098_ (.A2(_00607_),
    .A1(_00601_),
    .B1(_00606_),
    .X(_01736_));
 sg13g2_nor2_1 _12099_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sg13g2_or2_1 _12100_ (.X(_01738_),
    .B(_01737_),
    .A(_01734_));
 sg13g2_inv_1 _12101_ (.Y(_01739_),
    .A(_01738_));
 sg13g2_nand2b_1 _12102_ (.Y(_01740_),
    .B(_01738_),
    .A_N(_01732_));
 sg13g2_inv_1 _12103_ (.Y(_01741_),
    .A(_01740_));
 sg13g2_nand2_1 _12104_ (.Y(_01742_),
    .A(_01732_),
    .B(_01739_));
 sg13g2_o21ai_1 _12105_ (.B1(_01742_),
    .Y(_01743_),
    .A1(_01726_),
    .A2(_01741_));
 sg13g2_or2_1 _12106_ (.X(_01744_),
    .B(_01742_),
    .A(_01726_));
 sg13g2_a22oi_1 _12107_ (.Y(_01745_),
    .B1(_01743_),
    .B2(_01744_),
    .A2(_01741_),
    .A1(_01726_));
 sg13g2_nor2b_1 _12108_ (.A(_01723_),
    .B_N(_01745_),
    .Y(_01746_));
 sg13g2_nor3_1 _12109_ (.A(_01674_),
    .B(_01724_),
    .C(_01746_),
    .Y(_01747_));
 sg13g2_o21ai_1 _12110_ (.B1(_01674_),
    .Y(_01748_),
    .A1(_01724_),
    .A2(_01746_));
 sg13g2_o21ai_1 _12111_ (.B1(_01748_),
    .Y(_01749_),
    .A1(_01589_),
    .A2(_01747_));
 sg13g2_nand2b_1 _12112_ (.Y(_01750_),
    .B(_01748_),
    .A_N(_01747_));
 sg13g2_xnor2_1 _12113_ (.Y(_01751_),
    .A(_01589_),
    .B(_01750_));
 sg13g2_xor2_1 _12114_ (.B(_01591_),
    .A(_01590_),
    .X(_01752_));
 sg13g2_xnor2_1 _12115_ (.Y(_01753_),
    .A(_09554_),
    .B(_01620_));
 sg13g2_xnor2_1 _12116_ (.Y(_01754_),
    .A(_01624_),
    .B(_01753_));
 sg13g2_nand2b_1 _12117_ (.Y(_01755_),
    .B(_01752_),
    .A_N(_01754_));
 sg13g2_nand2b_1 _12118_ (.Y(_01756_),
    .B(_01754_),
    .A_N(_01752_));
 sg13g2_nor2_1 _12119_ (.A(_01629_),
    .B(_01630_),
    .Y(_01757_));
 sg13g2_xor2_1 _12120_ (.B(_01757_),
    .A(_01631_),
    .X(_01758_));
 sg13g2_nand2b_1 _12121_ (.Y(_01759_),
    .B(_01755_),
    .A_N(_01758_));
 sg13g2_nand2b_1 _12122_ (.Y(_01760_),
    .B(_01718_),
    .A_N(_01717_));
 sg13g2_xor2_1 _12123_ (.B(_01760_),
    .A(_01720_),
    .X(_01761_));
 sg13g2_nor2b_1 _12124_ (.A(_01729_),
    .B_N(_01730_),
    .Y(_01762_));
 sg13g2_xnor2_1 _12125_ (.Y(_01763_),
    .A(_01731_),
    .B(_01762_));
 sg13g2_xnor2_1 _12126_ (.Y(_01764_),
    .A(_01761_),
    .B(_01763_));
 sg13g2_nor2_1 _12127_ (.A(_01734_),
    .B(_01735_),
    .Y(_01765_));
 sg13g2_xor2_1 _12128_ (.B(_01765_),
    .A(_01736_),
    .X(_01766_));
 sg13g2_xnor2_1 _12129_ (.Y(_01767_),
    .A(_01764_),
    .B(_01766_));
 sg13g2_nor2b_1 _12130_ (.A(_01693_),
    .B_N(_01694_),
    .Y(_01768_));
 sg13g2_xnor2_1 _12131_ (.Y(_01769_),
    .A(_08608_),
    .B(_01768_));
 sg13g2_nor2b_1 _12132_ (.A(_01699_),
    .B_N(_01700_),
    .Y(_01770_));
 sg13g2_xnor2_1 _12133_ (.Y(_01771_),
    .A(_01702_),
    .B(_01770_));
 sg13g2_nand2b_1 _12134_ (.Y(_01772_),
    .B(_01769_),
    .A_N(_01771_));
 sg13g2_nor2b_1 _12135_ (.A(_01769_),
    .B_N(_01771_),
    .Y(_01773_));
 sg13g2_xnor2_1 _12136_ (.Y(_01774_),
    .A(_01769_),
    .B(_01771_));
 sg13g2_xor2_1 _12137_ (.B(_01707_),
    .A(_01705_),
    .X(_01775_));
 sg13g2_xnor2_1 _12138_ (.Y(_01776_),
    .A(_01710_),
    .B(_01775_));
 sg13g2_xnor2_1 _12139_ (.Y(_01777_),
    .A(_01774_),
    .B(_01776_));
 sg13g2_or2_1 _12140_ (.X(_01778_),
    .B(_01777_),
    .A(_01767_));
 sg13g2_nand2_1 _12141_ (.Y(_01779_),
    .A(_01767_),
    .B(_01777_));
 sg13g2_a21o_1 _12142_ (.A2(_01603_),
    .A1(_01600_),
    .B1(_01604_),
    .X(_01780_));
 sg13g2_o21ai_1 _12143_ (.B1(_01780_),
    .Y(_01781_),
    .A1(_01601_),
    .A2(_01603_));
 sg13g2_nand2_1 _12144_ (.Y(_01782_),
    .A(_01778_),
    .B(_01781_));
 sg13g2_nand2_1 _12145_ (.Y(_01783_),
    .A(_01779_),
    .B(_01782_));
 sg13g2_a21oi_1 _12146_ (.A1(_01756_),
    .A2(_01759_),
    .Y(_01784_),
    .B1(_01783_));
 sg13g2_and3_1 _12147_ (.X(_01785_),
    .A(_01756_),
    .B(_01759_),
    .C(_01783_));
 sg13g2_nor2_1 _12148_ (.A(_01784_),
    .B(_01785_),
    .Y(_01786_));
 sg13g2_nand2_1 _12149_ (.Y(_01787_),
    .A(_01657_),
    .B(_01658_));
 sg13g2_xor2_1 _12150_ (.B(_01787_),
    .A(_00596_),
    .X(_01788_));
 sg13g2_inv_1 _12151_ (.Y(_01789_),
    .A(_01788_));
 sg13g2_nor2_1 _12152_ (.A(_01637_),
    .B(_01638_),
    .Y(_01790_));
 sg13g2_xor2_1 _12153_ (.B(_01790_),
    .A(_00517_),
    .X(_01791_));
 sg13g2_nand2_1 _12154_ (.Y(_01792_),
    .A(_01789_),
    .B(_01791_));
 sg13g2_nand2_1 _12155_ (.Y(_01793_),
    .A(_01663_),
    .B(_01664_));
 sg13g2_xor2_1 _12156_ (.B(_01793_),
    .A(_01665_),
    .X(_01794_));
 sg13g2_o21ai_1 _12157_ (.B1(_01794_),
    .Y(_01795_),
    .A1(_01789_),
    .A2(_01791_));
 sg13g2_nand2_1 _12158_ (.Y(_01796_),
    .A(_01792_),
    .B(_01795_));
 sg13g2_xnor2_1 _12159_ (.Y(_01797_),
    .A(_01786_),
    .B(_01796_));
 sg13g2_xnor2_1 _12160_ (.Y(_01798_),
    .A(_01788_),
    .B(_01791_));
 sg13g2_xnor2_1 _12161_ (.Y(_01799_),
    .A(_01794_),
    .B(_01798_));
 sg13g2_xnor2_1 _12162_ (.Y(_01800_),
    .A(_01752_),
    .B(_01754_));
 sg13g2_xnor2_1 _12163_ (.Y(_01801_),
    .A(_01758_),
    .B(_01800_));
 sg13g2_xnor2_1 _12164_ (.Y(_01802_),
    .A(_01645_),
    .B(_01647_));
 sg13g2_xnor2_1 _12165_ (.Y(_01803_),
    .A(_01651_),
    .B(_01802_));
 sg13g2_nor2_1 _12166_ (.A(_01678_),
    .B(_01679_),
    .Y(_01804_));
 sg13g2_xor2_1 _12167_ (.B(_01804_),
    .A(_01680_),
    .X(_01805_));
 sg13g2_nand2_1 _12168_ (.Y(_01806_),
    .A(_01803_),
    .B(_01805_));
 sg13g2_xor2_1 _12169_ (.B(_01805_),
    .A(_01803_),
    .X(_01807_));
 sg13g2_nor2_1 _12170_ (.A(_01685_),
    .B(_01686_),
    .Y(_01808_));
 sg13g2_xor2_1 _12171_ (.B(_01808_),
    .A(_01687_),
    .X(_01809_));
 sg13g2_xnor2_1 _12172_ (.Y(_01810_),
    .A(_01807_),
    .B(_01809_));
 sg13g2_a21o_1 _12173_ (.A2(_01801_),
    .A1(_01799_),
    .B1(_01810_),
    .X(_01811_));
 sg13g2_o21ai_1 _12174_ (.B1(_01811_),
    .Y(_01812_),
    .A1(_01799_),
    .A2(_01801_));
 sg13g2_inv_1 _12175_ (.Y(_01813_),
    .A(_01812_));
 sg13g2_o21ai_1 _12176_ (.B1(_06485_),
    .Y(_01814_),
    .A1(_06474_),
    .A2(_06518_));
 sg13g2_inv_1 _12177_ (.Y(_01815_),
    .A(_01814_));
 sg13g2_nand2_1 _12178_ (.Y(_01816_),
    .A(_01778_),
    .B(_01779_));
 sg13g2_xor2_1 _12179_ (.B(_01816_),
    .A(_01781_),
    .X(_01817_));
 sg13g2_xnor2_1 _12180_ (.Y(_01818_),
    .A(_01799_),
    .B(_01801_));
 sg13g2_xnor2_1 _12181_ (.Y(_01819_),
    .A(_01810_),
    .B(_01818_));
 sg13g2_nor2_1 _12182_ (.A(_01817_),
    .B(_01819_),
    .Y(_01820_));
 sg13g2_a21o_1 _12183_ (.A2(_01612_),
    .A1(_01610_),
    .B1(_01613_),
    .X(_01821_));
 sg13g2_o21ai_1 _12184_ (.B1(_01821_),
    .Y(_01822_),
    .A1(_01609_),
    .A2(_01612_));
 sg13g2_and2_1 _12185_ (.A(_01820_),
    .B(_01822_),
    .X(_01823_));
 sg13g2_nand2_1 _12186_ (.Y(_01824_),
    .A(_01817_),
    .B(_01819_));
 sg13g2_o21ai_1 _12187_ (.B1(_01824_),
    .Y(_01825_),
    .A1(_01820_),
    .A2(_01822_));
 sg13g2_nor2_1 _12188_ (.A(_01823_),
    .B(_01825_),
    .Y(_01826_));
 sg13g2_nor2_1 _12189_ (.A(_01822_),
    .B(_01824_),
    .Y(_01827_));
 sg13g2_or2_1 _12190_ (.X(_01828_),
    .B(_01827_),
    .A(_01826_));
 sg13g2_nand2_1 _12191_ (.Y(_01829_),
    .A(_01814_),
    .B(_01823_));
 sg13g2_o21ai_1 _12192_ (.B1(_01825_),
    .Y(_01830_),
    .A1(_01815_),
    .A2(_01827_));
 sg13g2_a22oi_1 _12193_ (.Y(_01831_),
    .B1(_01830_),
    .B2(_01812_),
    .A2(_01823_),
    .A1(_01814_));
 sg13g2_nand3_1 _12194_ (.B(_01829_),
    .C(_01830_),
    .A(_01813_),
    .Y(_01832_));
 sg13g2_a21o_1 _12195_ (.A2(_01830_),
    .A1(_01829_),
    .B1(_01813_),
    .X(_01833_));
 sg13g2_nand3_1 _12196_ (.B(_01832_),
    .C(_01833_),
    .A(_01797_),
    .Y(_01834_));
 sg13g2_a21o_1 _12197_ (.A2(_01833_),
    .A1(_01832_),
    .B1(_01797_),
    .X(_01835_));
 sg13g2_a21o_1 _12198_ (.A2(_01776_),
    .A1(_01772_),
    .B1(_01773_),
    .X(_01836_));
 sg13g2_o21ai_1 _12199_ (.B1(_01809_),
    .Y(_01837_),
    .A1(_01803_),
    .A2(_01805_));
 sg13g2_and3_1 _12200_ (.X(_01838_),
    .A(_01806_),
    .B(_01836_),
    .C(_01837_));
 sg13g2_a21oi_1 _12201_ (.A1(_01806_),
    .A2(_01837_),
    .Y(_01839_),
    .B1(_01836_));
 sg13g2_nor2_1 _12202_ (.A(_01838_),
    .B(_01839_),
    .Y(_01840_));
 sg13g2_a21o_1 _12203_ (.A2(_01763_),
    .A1(_01761_),
    .B1(_01766_),
    .X(_01841_));
 sg13g2_o21ai_1 _12204_ (.B1(_01841_),
    .Y(_01842_),
    .A1(_01761_),
    .A2(_01763_));
 sg13g2_xor2_1 _12205_ (.B(_01842_),
    .A(_01840_),
    .X(_01843_));
 sg13g2_nand2_1 _12206_ (.Y(_01844_),
    .A(_01835_),
    .B(_01843_));
 sg13g2_nand2_1 _12207_ (.Y(_01845_),
    .A(_01834_),
    .B(_01844_));
 sg13g2_and3_1 _12208_ (.X(_01846_),
    .A(_01834_),
    .B(_01835_),
    .C(_01843_));
 sg13g2_a21oi_1 _12209_ (.A1(_01834_),
    .A2(_01835_),
    .Y(_01847_),
    .B1(_01843_));
 sg13g2_nand2_1 _12210_ (.Y(_01848_),
    .A(_01643_),
    .B(_01644_));
 sg13g2_xnor2_1 _12211_ (.Y(_01849_),
    .A(_01672_),
    .B(_01848_));
 sg13g2_o21ai_1 _12212_ (.B1(_01849_),
    .Y(_01850_),
    .A1(_01846_),
    .A2(_01847_));
 sg13g2_nor3_1 _12213_ (.A(_01846_),
    .B(_01847_),
    .C(_01849_),
    .Y(_01851_));
 sg13g2_nor2_1 _12214_ (.A(_01723_),
    .B(_01724_),
    .Y(_01852_));
 sg13g2_xnor2_1 _12215_ (.Y(_01853_),
    .A(_01745_),
    .B(_01852_));
 sg13g2_a21oi_2 _12216_ (.B1(_01851_),
    .Y(_01854_),
    .A2(_01853_),
    .A1(_01850_));
 sg13g2_or2_1 _12217_ (.X(_01855_),
    .B(_01853_),
    .A(_01850_));
 sg13g2_and2_1 _12218_ (.A(_01851_),
    .B(_01853_),
    .X(_01856_));
 sg13g2_a21o_1 _12219_ (.A2(_01855_),
    .A1(_01854_),
    .B1(_01856_),
    .X(_01857_));
 sg13g2_a21oi_1 _12220_ (.A1(_01579_),
    .A2(_01580_),
    .Y(_01858_),
    .B1(_01587_));
 sg13g2_a21o_1 _12221_ (.A2(_01589_),
    .A1(_01579_),
    .B1(_01858_),
    .X(_01859_));
 sg13g2_inv_1 _12222_ (.Y(_01860_),
    .A(_01859_));
 sg13g2_nor2_1 _12223_ (.A(_01857_),
    .B(_01860_),
    .Y(_01861_));
 sg13g2_nor2_1 _12224_ (.A(_01854_),
    .B(_01861_),
    .Y(_01862_));
 sg13g2_nor2_1 _12225_ (.A(_01855_),
    .B(_01860_),
    .Y(_01863_));
 sg13g2_nand2b_1 _12226_ (.Y(_01864_),
    .B(_01859_),
    .A_N(_01855_));
 sg13g2_o21ai_1 _12227_ (.B1(_01864_),
    .Y(_01865_),
    .A1(_01854_),
    .A2(_01861_));
 sg13g2_xnor2_1 _12228_ (.Y(_01866_),
    .A(_01845_),
    .B(_01865_));
 sg13g2_nand2_1 _12229_ (.Y(_01867_),
    .A(_01751_),
    .B(_01866_));
 sg13g2_nor2_1 _12230_ (.A(_01751_),
    .B(_01866_),
    .Y(_01868_));
 sg13g2_xor2_1 _12231_ (.B(_01866_),
    .A(_01751_),
    .X(_01869_));
 sg13g2_nor2_1 _12232_ (.A(_01785_),
    .B(_01796_),
    .Y(_01870_));
 sg13g2_or2_1 _12233_ (.X(_01871_),
    .B(_01870_),
    .A(_01784_));
 sg13g2_nand2_1 _12234_ (.Y(_01872_),
    .A(_01831_),
    .B(_01871_));
 sg13g2_xor2_1 _12235_ (.B(_01871_),
    .A(_01831_),
    .X(_01873_));
 sg13g2_nor2_1 _12236_ (.A(_01838_),
    .B(_01842_),
    .Y(_01874_));
 sg13g2_nor2_2 _12237_ (.A(_01839_),
    .B(_01874_),
    .Y(_01875_));
 sg13g2_xnor2_1 _12238_ (.Y(_01876_),
    .A(_01873_),
    .B(_01875_));
 sg13g2_xnor2_1 _12239_ (.Y(_01877_),
    .A(_01869_),
    .B(_01876_));
 sg13g2_nand2_1 _12240_ (.Y(_01878_),
    .A(_01689_),
    .B(_01695_));
 sg13g2_nand2_2 _12241_ (.Y(_01879_),
    .A(_01690_),
    .B(_01878_));
 sg13g2_nand2_1 _12242_ (.Y(_01880_),
    .A(_01712_),
    .B(_01721_));
 sg13g2_nand2_2 _12243_ (.Y(_01881_),
    .A(_01713_),
    .B(_01880_));
 sg13g2_xor2_1 _12244_ (.B(_01881_),
    .A(_01879_),
    .X(_01882_));
 sg13g2_xnor2_1 _12245_ (.Y(_01883_),
    .A(_01743_),
    .B(_01882_));
 sg13g2_o21ai_1 _12246_ (.B1(_01668_),
    .Y(_01884_),
    .A1(_01653_),
    .A2(_01670_));
 sg13g2_a21oi_1 _12247_ (.A1(_01592_),
    .A2(_01615_),
    .Y(_01885_),
    .B1(_01616_));
 sg13g2_nand2_1 _12248_ (.Y(_01886_),
    .A(_01641_),
    .B(_01885_));
 sg13g2_nor2_1 _12249_ (.A(_01641_),
    .B(_01885_),
    .Y(_01887_));
 sg13g2_a21oi_2 _12250_ (.B1(_01887_),
    .Y(_01888_),
    .A2(_01886_),
    .A1(_01884_));
 sg13g2_o21ai_1 _12251_ (.B1(_01888_),
    .Y(_01889_),
    .A1(_01884_),
    .A2(_01886_));
 sg13g2_nand2_1 _12252_ (.Y(_01890_),
    .A(_01884_),
    .B(_01887_));
 sg13g2_nand2_1 _12253_ (.Y(_01891_),
    .A(_01889_),
    .B(_01890_));
 sg13g2_nor2b_1 _12254_ (.A(_01883_),
    .B_N(_01891_),
    .Y(_01892_));
 sg13g2_nand2b_1 _12255_ (.Y(_01893_),
    .B(_01883_),
    .A_N(_01891_));
 sg13g2_nor2b_1 _12256_ (.A(_01892_),
    .B_N(_01893_),
    .Y(_01894_));
 sg13g2_nand2_1 _12257_ (.Y(_01895_),
    .A(_01568_),
    .B(_01577_));
 sg13g2_nand2_2 _12258_ (.Y(_01896_),
    .A(_01569_),
    .B(_01895_));
 sg13g2_xnor2_1 _12259_ (.Y(_01897_),
    .A(_01894_),
    .B(_01896_));
 sg13g2_a21oi_1 _12260_ (.A1(_01867_),
    .A2(_01876_),
    .Y(_01898_),
    .B1(_01868_));
 sg13g2_o21ai_1 _12261_ (.B1(_01898_),
    .Y(_01899_),
    .A1(_01877_),
    .A2(_01897_));
 sg13g2_nand3b_1 _12262_ (.B(_01876_),
    .C(_01868_),
    .Y(_01900_),
    .A_N(_01897_));
 sg13g2_nand2_1 _12263_ (.Y(_01901_),
    .A(_01899_),
    .B(_01900_));
 sg13g2_o21ai_1 _12264_ (.B1(_01893_),
    .Y(_01902_),
    .A1(_01892_),
    .A2(_01896_));
 sg13g2_xor2_1 _12265_ (.B(_01902_),
    .A(_01901_),
    .X(_01903_));
 sg13g2_nor2_1 _12266_ (.A(_01845_),
    .B(_01862_),
    .Y(_01904_));
 sg13g2_nor2_1 _12267_ (.A(_01863_),
    .B(_01904_),
    .Y(_01905_));
 sg13g2_o21ai_1 _12268_ (.B1(_01749_),
    .Y(_01906_),
    .A1(_01863_),
    .A2(_01904_));
 sg13g2_nor3_1 _12269_ (.A(_01749_),
    .B(_01863_),
    .C(_01904_),
    .Y(_01907_));
 sg13g2_xnor2_1 _12270_ (.Y(_01908_),
    .A(_01749_),
    .B(_01905_));
 sg13g2_o21ai_1 _12271_ (.B1(_01875_),
    .Y(_01909_),
    .A1(_01831_),
    .A2(_01871_));
 sg13g2_nand2_1 _12272_ (.Y(_01910_),
    .A(_01872_),
    .B(_01909_));
 sg13g2_xnor2_1 _12273_ (.Y(_01911_),
    .A(_01908_),
    .B(_01910_));
 sg13g2_nor2_1 _12274_ (.A(_01903_),
    .B(_01911_),
    .Y(_01912_));
 sg13g2_nand2_1 _12275_ (.Y(_01913_),
    .A(_01903_),
    .B(_01911_));
 sg13g2_o21ai_1 _12276_ (.B1(_01913_),
    .Y(_01914_),
    .A1(_01888_),
    .A2(_01912_));
 sg13g2_or2_1 _12277_ (.X(_01915_),
    .B(_01913_),
    .A(_01888_));
 sg13g2_nand2_1 _12278_ (.Y(_01916_),
    .A(_01888_),
    .B(_01912_));
 sg13g2_a22oi_1 _12279_ (.Y(_01917_),
    .B1(_01914_),
    .B2(_01915_),
    .A2(_01912_),
    .A1(_01888_));
 sg13g2_a21o_1 _12280_ (.A2(_01881_),
    .A1(_01879_),
    .B1(_01743_),
    .X(_01918_));
 sg13g2_o21ai_1 _12281_ (.B1(_01918_),
    .Y(_01919_),
    .A1(_01879_),
    .A2(_01881_));
 sg13g2_inv_1 _12282_ (.Y(_01920_),
    .A(_01919_));
 sg13g2_a21oi_1 _12283_ (.A1(_01916_),
    .A2(_01920_),
    .Y(_01921_),
    .B1(_01914_));
 sg13g2_nor2_1 _12284_ (.A(_01915_),
    .B(_01919_),
    .Y(_01922_));
 sg13g2_nand2_1 _12285_ (.Y(_01923_),
    .A(_01900_),
    .B(_01902_));
 sg13g2_nand2_1 _12286_ (.Y(_01924_),
    .A(_01899_),
    .B(_01923_));
 sg13g2_nor2b_1 _12287_ (.A(_01922_),
    .B_N(_01924_),
    .Y(_01925_));
 sg13g2_o21ai_1 _12288_ (.B1(_01906_),
    .Y(_01926_),
    .A1(_01907_),
    .A2(_01910_));
 sg13g2_nor2_1 _12289_ (.A(_01921_),
    .B(_01922_),
    .Y(_01927_));
 sg13g2_xnor2_1 _12290_ (.Y(_01928_),
    .A(_01924_),
    .B(_01927_));
 sg13g2_nand2_1 _12291_ (.Y(_01929_),
    .A(_01926_),
    .B(_01928_));
 sg13g2_o21ai_1 _12292_ (.B1(_01929_),
    .Y(_01930_),
    .A1(_01921_),
    .A2(_01925_));
 sg13g2_xnor2_1 _12293_ (.Y(_01931_),
    .A(_01926_),
    .B(_01928_));
 sg13g2_xnor2_1 _12294_ (.Y(_01932_),
    .A(_01492_),
    .B(_01545_));
 sg13g2_xor2_1 _12295_ (.B(_01529_),
    .A(_01527_),
    .X(_01933_));
 sg13g2_xor2_1 _12296_ (.B(_01897_),
    .A(_01877_),
    .X(_01934_));
 sg13g2_xnor2_1 _12297_ (.Y(_01935_),
    .A(_01217_),
    .B(_01287_));
 sg13g2_nand2b_1 _12298_ (.Y(_01936_),
    .B(_00643_),
    .A_N(_01935_));
 sg13g2_xnor2_1 _12299_ (.Y(_01937_),
    .A(_01380_),
    .B(_01382_));
 sg13g2_xnor2_1 _12300_ (.Y(_01938_),
    .A(_01815_),
    .B(_01828_));
 sg13g2_nor2_1 _12301_ (.A(_01936_),
    .B(_01937_),
    .Y(_01939_));
 sg13g2_nor2_1 _12302_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sg13g2_a21oi_2 _12303_ (.B1(_01940_),
    .Y(_01941_),
    .A2(_01937_),
    .A1(_01936_));
 sg13g2_xor2_1 _12304_ (.B(_01469_),
    .A(_01456_),
    .X(_01942_));
 sg13g2_xnor2_1 _12305_ (.Y(_01943_),
    .A(_01857_),
    .B(_01860_));
 sg13g2_nor2_1 _12306_ (.A(_01941_),
    .B(_01943_),
    .Y(_01944_));
 sg13g2_nand2_1 _12307_ (.Y(_01945_),
    .A(_01941_),
    .B(_01943_));
 sg13g2_a21oi_1 _12308_ (.A1(_01942_),
    .A2(_01945_),
    .Y(_01946_),
    .B1(_01944_));
 sg13g2_nand2_1 _12309_ (.Y(_01947_),
    .A(_01933_),
    .B(_01946_));
 sg13g2_nand2_1 _12310_ (.Y(_01948_),
    .A(_01934_),
    .B(_01947_));
 sg13g2_o21ai_1 _12311_ (.B1(_01948_),
    .Y(_01949_),
    .A1(_01933_),
    .A2(_01946_));
 sg13g2_xnor2_1 _12312_ (.Y(_01950_),
    .A(_01509_),
    .B(_01539_));
 sg13g2_xnor2_1 _12313_ (.Y(_01951_),
    .A(_01917_),
    .B(_01920_));
 sg13g2_nand2_1 _12314_ (.Y(_01952_),
    .A(_01949_),
    .B(_01950_));
 sg13g2_nor2_1 _12315_ (.A(_01949_),
    .B(_01950_),
    .Y(_01953_));
 sg13g2_a21oi_1 _12316_ (.A1(_01951_),
    .A2(_01952_),
    .Y(_01954_),
    .B1(_01953_));
 sg13g2_nand2_1 _12317_ (.Y(_01955_),
    .A(_01932_),
    .B(_01954_));
 sg13g2_nand2_1 _12318_ (.Y(_01956_),
    .A(_01931_),
    .B(_01955_));
 sg13g2_nor2_1 _12319_ (.A(_01547_),
    .B(_01930_),
    .Y(_01957_));
 sg13g2_nor2_1 _12320_ (.A(_01932_),
    .B(_01954_),
    .Y(_01958_));
 sg13g2_nor2_1 _12321_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sg13g2_a22oi_1 _12322_ (.Y(_01960_),
    .B1(_01956_),
    .B2(_01959_),
    .A2(_01930_),
    .A1(_01547_));
 sg13g2_inv_4 _12323_ (.A(_01960_),
    .Y(_01961_));
 sg13g2_mux2_2 _12324_ (.A0(_00643_),
    .A1(_01935_),
    .S(_01960_),
    .X(_01962_));
 sg13g2_a22oi_1 _12325_ (.Y(_01963_),
    .B1(_05528_),
    .B2(net2417),
    .A2(net2612),
    .A1(net2555));
 sg13g2_o21ai_1 _12326_ (.B1(net2693),
    .Y(_01964_),
    .A1(net2741),
    .A2(net2608));
 sg13g2_nor2_1 _12327_ (.A(net2782),
    .B(_01964_),
    .Y(_01965_));
 sg13g2_xor2_1 _12328_ (.B(net2427),
    .A(net2297),
    .X(_01966_));
 sg13g2_nor2b_1 _12329_ (.A(_01965_),
    .B_N(_01966_),
    .Y(_01967_));
 sg13g2_nor3_1 _12330_ (.A(net2781),
    .B(_01964_),
    .C(_01966_),
    .Y(_01968_));
 sg13g2_inv_1 _12331_ (.Y(_01969_),
    .A(_01968_));
 sg13g2_nor2_1 _12332_ (.A(_01967_),
    .B(_01968_),
    .Y(_01970_));
 sg13g2_xnor2_1 _12333_ (.Y(_01971_),
    .A(_01963_),
    .B(_01970_));
 sg13g2_xnor2_1 _12334_ (.Y(_01972_),
    .A(net2297),
    .B(net2386));
 sg13g2_xnor2_1 _12335_ (.Y(_01973_),
    .A(net2789),
    .B(net2798));
 sg13g2_nand2_2 _12336_ (.Y(_01974_),
    .A(_01972_),
    .B(_01973_));
 sg13g2_nor2b_1 _12337_ (.A(net2454),
    .B_N(net2474),
    .Y(_01975_));
 sg13g2_nand2b_1 _12338_ (.Y(_01976_),
    .B(net2474),
    .A_N(net2456));
 sg13g2_nand2_2 _12339_ (.Y(_01977_),
    .A(_05242_),
    .B(\net.in[59] ));
 sg13g2_xnor2_1 _12340_ (.Y(_01978_),
    .A(net2331),
    .B(\net.in[242] ));
 sg13g2_nand3_1 _12341_ (.B(_01977_),
    .C(_01978_),
    .A(_01975_),
    .Y(_01979_));
 sg13g2_a21o_1 _12342_ (.A2(_01977_),
    .A1(_01975_),
    .B1(_01978_),
    .X(_01980_));
 sg13g2_nand2_1 _12343_ (.Y(_01981_),
    .A(_01979_),
    .B(_01980_));
 sg13g2_xor2_1 _12344_ (.B(_01981_),
    .A(_01974_),
    .X(_01982_));
 sg13g2_nor2_1 _12345_ (.A(_01971_),
    .B(_01982_),
    .Y(_01983_));
 sg13g2_xor2_1 _12346_ (.B(_01982_),
    .A(_01971_),
    .X(_01984_));
 sg13g2_nand2b_2 _12347_ (.Y(_01985_),
    .B(net2479),
    .A_N(\net.in[140] ));
 sg13g2_xnor2_1 _12348_ (.Y(_01986_),
    .A(net2487),
    .B(net2528));
 sg13g2_o21ai_1 _12349_ (.B1(_01986_),
    .Y(_01987_),
    .A1(net2331),
    .A2(net2693));
 sg13g2_nor2b_1 _12350_ (.A(net2339),
    .B_N(net2321),
    .Y(_01988_));
 sg13g2_xnor2_1 _12351_ (.Y(_01989_),
    .A(net2420),
    .B(_01988_));
 sg13g2_nand2_1 _12352_ (.Y(_01990_),
    .A(_01987_),
    .B(_01989_));
 sg13g2_or2_1 _12353_ (.X(_01991_),
    .B(_01989_),
    .A(_01987_));
 sg13g2_nand2_1 _12354_ (.Y(_01992_),
    .A(_01990_),
    .B(_01991_));
 sg13g2_xnor2_1 _12355_ (.Y(_01993_),
    .A(_01985_),
    .B(_01992_));
 sg13g2_xnor2_1 _12356_ (.Y(_01994_),
    .A(_01984_),
    .B(_01993_));
 sg13g2_xnor2_1 _12357_ (.Y(_01995_),
    .A(net2313),
    .B(net2239));
 sg13g2_xnor2_1 _12358_ (.Y(_01996_),
    .A(net2273),
    .B(net2238));
 sg13g2_nand2_1 _12359_ (.Y(_01997_),
    .A(_01995_),
    .B(_01996_));
 sg13g2_and2_1 _12360_ (.A(net2518),
    .B(net2676),
    .X(_01998_));
 sg13g2_nor2_1 _12361_ (.A(net2518),
    .B(net2676),
    .Y(_01999_));
 sg13g2_nor2b_1 _12362_ (.A(net2569),
    .B_N(net2433),
    .Y(_02000_));
 sg13g2_nor3_2 _12363_ (.A(_01998_),
    .B(_01999_),
    .C(_02000_),
    .Y(_02001_));
 sg13g2_and2_1 _12364_ (.A(_01976_),
    .B(_02001_),
    .X(_02002_));
 sg13g2_nor2_1 _12365_ (.A(_01976_),
    .B(_02001_),
    .Y(_02003_));
 sg13g2_nor2_1 _12366_ (.A(_02002_),
    .B(_02003_),
    .Y(_02004_));
 sg13g2_xor2_1 _12367_ (.B(_02004_),
    .A(_01997_),
    .X(_02005_));
 sg13g2_nor2_1 _12368_ (.A(net2654),
    .B(net2739),
    .Y(_02006_));
 sg13g2_xnor2_1 _12369_ (.Y(_02007_),
    .A(net2653),
    .B(net2739));
 sg13g2_nand2b_1 _12370_ (.Y(_02008_),
    .B(net2522),
    .A_N(net2504));
 sg13g2_xnor2_1 _12371_ (.Y(_02009_),
    .A(net2234),
    .B(net2343));
 sg13g2_and2_1 _12372_ (.A(_02008_),
    .B(_02009_),
    .X(_02010_));
 sg13g2_nor2_2 _12373_ (.A(net2759),
    .B(net2778),
    .Y(_02011_));
 sg13g2_nand2_1 _12374_ (.Y(_02012_),
    .A(_02010_),
    .B(_02011_));
 sg13g2_nor2_1 _12375_ (.A(_02010_),
    .B(_02011_),
    .Y(_02013_));
 sg13g2_xnor2_1 _12376_ (.Y(_02014_),
    .A(_02010_),
    .B(_02011_));
 sg13g2_xnor2_1 _12377_ (.Y(_02015_),
    .A(_02007_),
    .B(_02014_));
 sg13g2_xnor2_1 _12378_ (.Y(_02016_),
    .A(net2518),
    .B(net2427));
 sg13g2_xnor2_1 _12379_ (.Y(_02017_),
    .A(net2356),
    .B(\net.in[237] ));
 sg13g2_nand2_2 _12380_ (.Y(_02018_),
    .A(_02016_),
    .B(_02017_));
 sg13g2_nor2_1 _12381_ (.A(net2582),
    .B(net2592),
    .Y(_02019_));
 sg13g2_xnor2_1 _12382_ (.Y(_02020_),
    .A(net2584),
    .B(net2595));
 sg13g2_xor2_1 _12383_ (.B(net2378),
    .A(net2443),
    .X(_02021_));
 sg13g2_nand2_1 _12384_ (.Y(_02022_),
    .A(_02020_),
    .B(_02021_));
 sg13g2_nor2_1 _12385_ (.A(_02020_),
    .B(_02021_),
    .Y(_02023_));
 sg13g2_xor2_1 _12386_ (.B(_02021_),
    .A(_02020_),
    .X(_02024_));
 sg13g2_xnor2_1 _12387_ (.Y(_02025_),
    .A(_02018_),
    .B(_02024_));
 sg13g2_nor2b_1 _12388_ (.A(_02025_),
    .B_N(_02015_),
    .Y(_02026_));
 sg13g2_nand2b_1 _12389_ (.Y(_02027_),
    .B(_02025_),
    .A_N(_02015_));
 sg13g2_xnor2_1 _12390_ (.Y(_02028_),
    .A(_02015_),
    .B(_02025_));
 sg13g2_xnor2_1 _12391_ (.Y(_02029_),
    .A(_02005_),
    .B(_02028_));
 sg13g2_nor2b_1 _12392_ (.A(\net.in[23] ),
    .B_N(net2678),
    .Y(_02030_));
 sg13g2_xnor2_1 _12393_ (.Y(_02031_),
    .A(net2693),
    .B(_02030_));
 sg13g2_nand2_1 _12394_ (.Y(_02032_),
    .A(net2644),
    .B(_02009_));
 sg13g2_nand2b_1 _12395_ (.Y(_02033_),
    .B(net2417),
    .A_N(net2781));
 sg13g2_xnor2_1 _12396_ (.Y(_02034_),
    .A(_06188_),
    .B(_02033_));
 sg13g2_o21ai_1 _12397_ (.B1(_02034_),
    .Y(_02035_),
    .A1(net2429),
    .A2(_02032_));
 sg13g2_or3_1 _12398_ (.A(net2425),
    .B(_02032_),
    .C(_02034_),
    .X(_02036_));
 sg13g2_nand2_1 _12399_ (.Y(_02037_),
    .A(_02035_),
    .B(_02036_));
 sg13g2_xor2_1 _12400_ (.B(_02037_),
    .A(_02031_),
    .X(_02038_));
 sg13g2_xnor2_1 _12401_ (.Y(_02039_),
    .A(net2297),
    .B(net2228));
 sg13g2_nor2_1 _12402_ (.A(net2612),
    .B(net2684),
    .Y(_02040_));
 sg13g2_nor3_1 _12403_ (.A(net2242),
    .B(net2778),
    .C(_02040_),
    .Y(_02041_));
 sg13g2_nor2_1 _12404_ (.A(net2275),
    .B(net2319),
    .Y(_02042_));
 sg13g2_nand2b_1 _12405_ (.Y(_02043_),
    .B(net2414),
    .A_N(net2308));
 sg13g2_xnor2_1 _12406_ (.Y(_02044_),
    .A(_02042_),
    .B(_02043_));
 sg13g2_nor4_1 _12407_ (.A(net2242),
    .B(net2779),
    .C(_02040_),
    .D(_02044_),
    .Y(_02045_));
 sg13g2_nand2b_1 _12408_ (.Y(_02046_),
    .B(_02044_),
    .A_N(_02041_));
 sg13g2_xnor2_1 _12409_ (.Y(_02047_),
    .A(_02041_),
    .B(_02044_));
 sg13g2_xnor2_1 _12410_ (.Y(_02048_),
    .A(_02039_),
    .B(_02047_));
 sg13g2_inv_1 _12411_ (.Y(_02049_),
    .A(_02048_));
 sg13g2_nor2_1 _12412_ (.A(net2486),
    .B(_05374_),
    .Y(_02050_));
 sg13g2_nor2_1 _12413_ (.A(net2443),
    .B(net2577),
    .Y(_02051_));
 sg13g2_xnor2_1 _12414_ (.Y(_02052_),
    .A(_02050_),
    .B(_02051_));
 sg13g2_nor2b_1 _12415_ (.A(net2788),
    .B_N(net2778),
    .Y(_02053_));
 sg13g2_nor2b_1 _12416_ (.A(net2778),
    .B_N(net2788),
    .Y(_02054_));
 sg13g2_nor2_1 _12417_ (.A(net2712),
    .B(net2704),
    .Y(_02055_));
 sg13g2_nor3_2 _12418_ (.A(_02053_),
    .B(_02054_),
    .C(_02055_),
    .Y(_02056_));
 sg13g2_xor2_1 _12419_ (.B(net2247),
    .A(net2185),
    .X(_02057_));
 sg13g2_xnor2_1 _12420_ (.Y(_02058_),
    .A(net2185),
    .B(net2247));
 sg13g2_nor3_2 _12421_ (.A(net2810),
    .B(net2778),
    .C(_02057_),
    .Y(_02059_));
 sg13g2_nor2_1 _12422_ (.A(_02056_),
    .B(_02059_),
    .Y(_02060_));
 sg13g2_xnor2_1 _12423_ (.Y(_02061_),
    .A(_02056_),
    .B(_02059_));
 sg13g2_xnor2_1 _12424_ (.Y(_02062_),
    .A(_02052_),
    .B(_02061_));
 sg13g2_nor2_1 _12425_ (.A(_02049_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_nand2_1 _12426_ (.Y(_02064_),
    .A(_02049_),
    .B(_02062_));
 sg13g2_a21oi_2 _12427_ (.B1(_02063_),
    .Y(_02065_),
    .A2(_02064_),
    .A1(_02038_));
 sg13g2_xnor2_1 _12428_ (.Y(_02066_),
    .A(_02048_),
    .B(_02062_));
 sg13g2_xnor2_1 _12429_ (.Y(_02067_),
    .A(_02038_),
    .B(_02066_));
 sg13g2_nand2_1 _12430_ (.Y(_02068_),
    .A(_02029_),
    .B(_02067_));
 sg13g2_nor2_1 _12431_ (.A(_02029_),
    .B(_02067_),
    .Y(_02069_));
 sg13g2_xor2_1 _12432_ (.B(_02067_),
    .A(_02029_),
    .X(_02070_));
 sg13g2_xnor2_1 _12433_ (.Y(_02071_),
    .A(_01994_),
    .B(_02070_));
 sg13g2_inv_1 _12434_ (.Y(_02072_),
    .A(_02071_));
 sg13g2_nor2_1 _12435_ (.A(net2433),
    .B(net2785),
    .Y(_02073_));
 sg13g2_xor2_1 _12436_ (.B(net2735),
    .A(net2353),
    .X(_02074_));
 sg13g2_xnor2_1 _12437_ (.Y(_02075_),
    .A(_02073_),
    .B(_02074_));
 sg13g2_xor2_1 _12438_ (.B(net2578),
    .A(net2718),
    .X(_02076_));
 sg13g2_or2_1 _12439_ (.X(_02077_),
    .B(\net.in[177] ),
    .A(net2474));
 sg13g2_xnor2_1 _12440_ (.Y(_02078_),
    .A(net2494),
    .B(net2377));
 sg13g2_nor3_1 _12441_ (.A(_08377_),
    .B(_02077_),
    .C(_02078_),
    .Y(_02079_));
 sg13g2_o21ai_1 _12442_ (.B1(_08377_),
    .Y(_02080_),
    .A1(_02077_),
    .A2(_02078_));
 sg13g2_nand2b_1 _12443_ (.Y(_02081_),
    .B(_02080_),
    .A_N(_02079_));
 sg13g2_xor2_1 _12444_ (.B(_02081_),
    .A(_02076_),
    .X(_02082_));
 sg13g2_nor2_1 _12445_ (.A(\net.in[38] ),
    .B(\net.in[242] ),
    .Y(_02083_));
 sg13g2_xnor2_1 _12446_ (.Y(_02084_),
    .A(net2698),
    .B(net2599));
 sg13g2_xnor2_1 _12447_ (.Y(_02085_),
    .A(_02083_),
    .B(_02084_));
 sg13g2_xor2_1 _12448_ (.B(net2703),
    .A(net2772),
    .X(_02086_));
 sg13g2_or2_1 _12449_ (.X(_02087_),
    .B(net2210),
    .A(\net.in[112] ));
 sg13g2_xnor2_1 _12450_ (.Y(_02088_),
    .A(net2584),
    .B(\net.in[97] ));
 sg13g2_o21ai_1 _12451_ (.B1(_02088_),
    .Y(_02089_),
    .A1(_02086_),
    .A2(_02087_));
 sg13g2_or3_1 _12452_ (.A(_02086_),
    .B(_02087_),
    .C(_02088_),
    .X(_02090_));
 sg13g2_nand2_1 _12453_ (.Y(_02091_),
    .A(_02089_),
    .B(_02090_));
 sg13g2_xnor2_1 _12454_ (.Y(_02092_),
    .A(_02085_),
    .B(_02091_));
 sg13g2_nand2_1 _12455_ (.Y(_02093_),
    .A(_02082_),
    .B(_02092_));
 sg13g2_xor2_1 _12456_ (.B(_02092_),
    .A(_02082_),
    .X(_02094_));
 sg13g2_nand2_1 _12457_ (.Y(_02095_),
    .A(_05770_),
    .B(net2286));
 sg13g2_o21ai_1 _12458_ (.B1(_02095_),
    .Y(_02096_),
    .A1(net2181),
    .A2(net2386));
 sg13g2_a21oi_2 _12459_ (.B1(_02096_),
    .Y(_02097_),
    .A2(net2386),
    .A1(net2181));
 sg13g2_xor2_1 _12460_ (.B(net2284),
    .A(\net.in[252] ),
    .X(_02098_));
 sg13g2_nor3_2 _12461_ (.A(_05715_),
    .B(net2546),
    .C(_02098_),
    .Y(_02099_));
 sg13g2_nor2b_1 _12462_ (.A(net2278),
    .B_N(net2640),
    .Y(_02100_));
 sg13g2_nor2b_1 _12463_ (.A(net2594),
    .B_N(net2297),
    .Y(_02101_));
 sg13g2_xnor2_1 _12464_ (.Y(_02102_),
    .A(_02100_),
    .B(_02101_));
 sg13g2_nor2b_1 _12465_ (.A(_02102_),
    .B_N(_02099_),
    .Y(_02103_));
 sg13g2_nor2b_1 _12466_ (.A(_02099_),
    .B_N(_02102_),
    .Y(_02104_));
 sg13g2_inv_1 _12467_ (.Y(_02105_),
    .A(_02104_));
 sg13g2_nor2_1 _12468_ (.A(_02103_),
    .B(_02104_),
    .Y(_02106_));
 sg13g2_xnor2_1 _12469_ (.Y(_02107_),
    .A(_02097_),
    .B(_02106_));
 sg13g2_xnor2_1 _12470_ (.Y(_02108_),
    .A(_02094_),
    .B(_02107_));
 sg13g2_xor2_1 _12471_ (.B(net2396),
    .A(net2474),
    .X(_02109_));
 sg13g2_a21oi_2 _12472_ (.B1(_02109_),
    .Y(_02110_),
    .A2(_05638_),
    .A1(_05583_));
 sg13g2_nor2b_1 _12473_ (.A(\net.in[81] ),
    .B_N(net2250),
    .Y(_02111_));
 sg13g2_nor2_1 _12474_ (.A(net2617),
    .B(\net.in[247] ),
    .Y(_02112_));
 sg13g2_xnor2_1 _12475_ (.Y(_02113_),
    .A(net2188),
    .B(net2196));
 sg13g2_o21ai_1 _12476_ (.B1(_02113_),
    .Y(_02114_),
    .A1(_02111_),
    .A2(_02112_));
 sg13g2_nor3_1 _12477_ (.A(_02111_),
    .B(_02112_),
    .C(_02113_),
    .Y(_02115_));
 sg13g2_inv_1 _12478_ (.Y(_02116_),
    .A(_02115_));
 sg13g2_nand2_1 _12479_ (.Y(_02117_),
    .A(_02114_),
    .B(_02116_));
 sg13g2_xnor2_1 _12480_ (.Y(_02118_),
    .A(_02110_),
    .B(_02117_));
 sg13g2_xnor2_1 _12481_ (.Y(_02119_),
    .A(net2425),
    .B(_00019_));
 sg13g2_xnor2_1 _12482_ (.Y(_02120_),
    .A(net2303),
    .B(_02119_));
 sg13g2_nand2b_1 _12483_ (.Y(_02121_),
    .B(net2284),
    .A_N(\net.in[80] ));
 sg13g2_nor2b_1 _12484_ (.A(net2353),
    .B_N(net2631),
    .Y(_02122_));
 sg13g2_xnor2_1 _12485_ (.Y(_02123_),
    .A(net2811),
    .B(net2778));
 sg13g2_nor2_2 _12486_ (.A(net2313),
    .B(\net.in[222] ),
    .Y(_02124_));
 sg13g2_a22oi_1 _12487_ (.Y(_02125_),
    .B1(_02123_),
    .B2(_02124_),
    .A2(_02122_),
    .A1(_02121_));
 sg13g2_and4_2 _12488_ (.A(_02121_),
    .B(_02122_),
    .C(_02123_),
    .D(_02124_),
    .X(_02126_));
 sg13g2_or3_1 _12489_ (.A(_02120_),
    .B(_02125_),
    .C(_02126_),
    .X(_02127_));
 sg13g2_o21ai_1 _12490_ (.B1(_02120_),
    .Y(_02128_),
    .A1(_02125_),
    .A2(_02126_));
 sg13g2_nor2_1 _12491_ (.A(net2744),
    .B(\net.in[81] ),
    .Y(_02129_));
 sg13g2_xnor2_1 _12492_ (.Y(_02130_),
    .A(net2427),
    .B(net2273));
 sg13g2_xnor2_1 _12493_ (.Y(_02131_),
    .A(net2474),
    .B(net2391));
 sg13g2_a21o_1 _12494_ (.A2(_02131_),
    .A1(_02130_),
    .B1(_02016_),
    .X(_02132_));
 sg13g2_nand3_1 _12495_ (.B(_02130_),
    .C(_02131_),
    .A(_02016_),
    .Y(_02133_));
 sg13g2_a21o_1 _12496_ (.A2(_02133_),
    .A1(_02132_),
    .B1(_02129_),
    .X(_02134_));
 sg13g2_nand3_1 _12497_ (.B(_02132_),
    .C(_02133_),
    .A(_02129_),
    .Y(_02135_));
 sg13g2_a22oi_1 _12498_ (.Y(_02136_),
    .B1(_02134_),
    .B2(_02135_),
    .A2(_02128_),
    .A1(_02127_));
 sg13g2_nand4_1 _12499_ (.B(_02128_),
    .C(_02134_),
    .A(_02127_),
    .Y(_02137_),
    .D(_02135_));
 sg13g2_nand2b_1 _12500_ (.Y(_02138_),
    .B(_02137_),
    .A_N(_02136_));
 sg13g2_o21ai_1 _12501_ (.B1(_02137_),
    .Y(_02139_),
    .A1(_02118_),
    .A2(_02136_));
 sg13g2_xnor2_1 _12502_ (.Y(_02140_),
    .A(_02118_),
    .B(_02138_));
 sg13g2_nor2_1 _12503_ (.A(_02108_),
    .B(_02140_),
    .Y(_02141_));
 sg13g2_nand2_1 _12504_ (.Y(_02142_),
    .A(_02108_),
    .B(_02140_));
 sg13g2_xnor2_1 _12505_ (.Y(_02143_),
    .A(_02108_),
    .B(_02140_));
 sg13g2_a21oi_1 _12506_ (.A1(_02075_),
    .A2(_02142_),
    .Y(_02144_),
    .B1(_02141_));
 sg13g2_xnor2_1 _12507_ (.Y(_02145_),
    .A(_02075_),
    .B(_02143_));
 sg13g2_nor2_1 _12508_ (.A(_02072_),
    .B(_02145_),
    .Y(_02146_));
 sg13g2_xnor2_1 _12509_ (.Y(_02147_),
    .A(_02071_),
    .B(_02145_));
 sg13g2_nand2_2 _12510_ (.Y(_02148_),
    .A(net2183),
    .B(net2621));
 sg13g2_o21ai_1 _12511_ (.B1(_02148_),
    .Y(_02149_),
    .A1(_05946_),
    .A2(\net.in[81] ));
 sg13g2_a21oi_2 _12512_ (.B1(_02149_),
    .Y(_02150_),
    .A2(\net.in[81] ),
    .A1(_05946_));
 sg13g2_nor2b_1 _12513_ (.A(net2578),
    .B_N(net2693),
    .Y(_02151_));
 sg13g2_xnor2_1 _12514_ (.Y(_02152_),
    .A(net2698),
    .B(_02151_));
 sg13g2_nor2_1 _12515_ (.A(net2794),
    .B(net2584),
    .Y(_02153_));
 sg13g2_xnor2_1 _12516_ (.Y(_02154_),
    .A(net2735),
    .B(_02153_));
 sg13g2_nand2_1 _12517_ (.Y(_02155_),
    .A(_02152_),
    .B(_02154_));
 sg13g2_nor2_1 _12518_ (.A(_02152_),
    .B(_02154_),
    .Y(_02156_));
 sg13g2_xnor2_1 _12519_ (.Y(_02157_),
    .A(_02152_),
    .B(_02154_));
 sg13g2_o21ai_1 _12520_ (.B1(_02155_),
    .Y(_02158_),
    .A1(_02150_),
    .A2(_02156_));
 sg13g2_xnor2_1 _12521_ (.Y(_02159_),
    .A(_02150_),
    .B(_02157_));
 sg13g2_xor2_1 _12522_ (.B(net2258),
    .A(net2384),
    .X(_02160_));
 sg13g2_a21oi_2 _12523_ (.B1(_09807_),
    .Y(_02161_),
    .A2(_07849_),
    .A1(net2535));
 sg13g2_nor2_1 _12524_ (.A(net2684),
    .B(net2459),
    .Y(_02162_));
 sg13g2_nor2_1 _12525_ (.A(net2356),
    .B(net2780),
    .Y(_02163_));
 sg13g2_xnor2_1 _12526_ (.Y(_02164_),
    .A(_02162_),
    .B(_02163_));
 sg13g2_xnor2_1 _12527_ (.Y(_02165_),
    .A(_02161_),
    .B(_02164_));
 sg13g2_xnor2_1 _12528_ (.Y(_02166_),
    .A(_02160_),
    .B(_02165_));
 sg13g2_nor2_1 _12529_ (.A(net2330),
    .B(net2644),
    .Y(_02167_));
 sg13g2_xnor2_1 _12530_ (.Y(_02168_),
    .A(_02006_),
    .B(_02167_));
 sg13g2_xor2_1 _12531_ (.B(net2644),
    .A(net2518),
    .X(_02169_));
 sg13g2_nand3_1 _12532_ (.B(_06056_),
    .C(_02169_),
    .A(_05121_),
    .Y(_02170_));
 sg13g2_nor2b_1 _12533_ (.A(net2318),
    .B_N(net2735),
    .Y(_02171_));
 sg13g2_xnor2_1 _12534_ (.Y(_02172_),
    .A(net2684),
    .B(_02171_));
 sg13g2_nand2b_1 _12535_ (.Y(_02173_),
    .B(_02172_),
    .A_N(_02170_));
 sg13g2_nand2b_1 _12536_ (.Y(_02174_),
    .B(_02170_),
    .A_N(_02172_));
 sg13g2_nand2_1 _12537_ (.Y(_02175_),
    .A(_02173_),
    .B(_02174_));
 sg13g2_xor2_1 _12538_ (.B(_02175_),
    .A(_02168_),
    .X(_02176_));
 sg13g2_nor2_1 _12539_ (.A(_02166_),
    .B(_02176_),
    .Y(_02177_));
 sg13g2_inv_1 _12540_ (.Y(_02178_),
    .A(_02177_));
 sg13g2_and2_1 _12541_ (.A(_02166_),
    .B(_02176_),
    .X(_02179_));
 sg13g2_nor2_1 _12542_ (.A(_02177_),
    .B(_02179_),
    .Y(_02180_));
 sg13g2_o21ai_1 _12543_ (.B1(_02178_),
    .Y(_02181_),
    .A1(_02159_),
    .A2(_02179_));
 sg13g2_xnor2_1 _12544_ (.Y(_02182_),
    .A(_02159_),
    .B(_02180_));
 sg13g2_xnor2_1 _12545_ (.Y(_02183_),
    .A(net2241),
    .B(net2185));
 sg13g2_xnor2_1 _12546_ (.Y(_02184_),
    .A(net2607),
    .B(net2704));
 sg13g2_nand2b_2 _12547_ (.Y(_02185_),
    .B(_02184_),
    .A_N(_02183_));
 sg13g2_xor2_1 _12548_ (.B(net2578),
    .A(net2723),
    .X(_02186_));
 sg13g2_nor2_2 _12549_ (.A(\net.in[191] ),
    .B(net2205),
    .Y(_02187_));
 sg13g2_nor2b_1 _12550_ (.A(net2262),
    .B_N(net2288),
    .Y(_02188_));
 sg13g2_xnor2_1 _12551_ (.Y(_02189_),
    .A(_02187_),
    .B(_02188_));
 sg13g2_nand2_1 _12552_ (.Y(_02190_),
    .A(_02186_),
    .B(_02189_));
 sg13g2_or2_1 _12553_ (.X(_02191_),
    .B(_02189_),
    .A(_02186_));
 sg13g2_nand2_1 _12554_ (.Y(_02192_),
    .A(_02190_),
    .B(_02191_));
 sg13g2_xor2_1 _12555_ (.B(_02192_),
    .A(_02185_),
    .X(_02193_));
 sg13g2_nor2b_2 _12556_ (.A(net2784),
    .B_N(net2672),
    .Y(_02194_));
 sg13g2_and3_2 _12557_ (.X(_02195_),
    .A(net2683),
    .B(net2621),
    .C(_02194_));
 sg13g2_and2_1 _12558_ (.A(net2377),
    .B(net2501),
    .X(_02196_));
 sg13g2_nor2_1 _12559_ (.A(net2376),
    .B(net2501),
    .Y(_02197_));
 sg13g2_nor4_2 _12560_ (.A(net2186),
    .B(net2273),
    .C(_02196_),
    .Y(_02198_),
    .D(_02197_));
 sg13g2_nor2_1 _12561_ (.A(net2678),
    .B(net2366),
    .Y(_02199_));
 sg13g2_nor2_2 _12562_ (.A(net2782),
    .B(_02199_),
    .Y(_02200_));
 sg13g2_xor2_1 _12563_ (.B(_02200_),
    .A(_02198_),
    .X(_02201_));
 sg13g2_xnor2_1 _12564_ (.Y(_02202_),
    .A(_02195_),
    .B(_02201_));
 sg13g2_xor2_1 _12565_ (.B(net2637),
    .A(net2303),
    .X(_02203_));
 sg13g2_xnor2_1 _12566_ (.Y(_02204_),
    .A(net2532),
    .B(net2446));
 sg13g2_nor2b_1 _12567_ (.A(net2247),
    .B_N(net2763),
    .Y(_02205_));
 sg13g2_nor2b_1 _12568_ (.A(net2352),
    .B_N(net2584),
    .Y(_02206_));
 sg13g2_xnor2_1 _12569_ (.Y(_02207_),
    .A(_02205_),
    .B(_02206_));
 sg13g2_nand2b_1 _12570_ (.Y(_02208_),
    .B(_02204_),
    .A_N(_02207_));
 sg13g2_nand2b_1 _12571_ (.Y(_02209_),
    .B(_02207_),
    .A_N(_02204_));
 sg13g2_xor2_1 _12572_ (.B(_02207_),
    .A(_02204_),
    .X(_02210_));
 sg13g2_xnor2_1 _12573_ (.Y(_02211_),
    .A(_02203_),
    .B(_02210_));
 sg13g2_nor2b_1 _12574_ (.A(_02202_),
    .B_N(_02211_),
    .Y(_02212_));
 sg13g2_nor2b_1 _12575_ (.A(_02211_),
    .B_N(_02202_),
    .Y(_02213_));
 sg13g2_xor2_1 _12576_ (.B(_02211_),
    .A(_02202_),
    .X(_02214_));
 sg13g2_xnor2_1 _12577_ (.Y(_02215_),
    .A(_02193_),
    .B(_02214_));
 sg13g2_xor2_1 _12578_ (.B(\net.in[80] ),
    .A(net2664),
    .X(_02216_));
 sg13g2_xor2_1 _12579_ (.B(net2739),
    .A(net2658),
    .X(_02217_));
 sg13g2_nor2_2 _12580_ (.A(_02216_),
    .B(_02217_),
    .Y(_02218_));
 sg13g2_o21ai_1 _12581_ (.B1(net2417),
    .Y(_02219_),
    .A1(net2771),
    .A2(net2701));
 sg13g2_nor2_2 _12582_ (.A(net2528),
    .B(_02219_),
    .Y(_02220_));
 sg13g2_nor2_1 _12583_ (.A(net2192),
    .B(\net.in[97] ),
    .Y(_02221_));
 sg13g2_xor2_1 _12584_ (.B(_02221_),
    .A(net2327),
    .X(_02222_));
 sg13g2_nand2_1 _12585_ (.Y(_02223_),
    .A(_02220_),
    .B(_02222_));
 sg13g2_or2_1 _12586_ (.X(_02224_),
    .B(_02222_),
    .A(_02220_));
 sg13g2_nand2_1 _12587_ (.Y(_02225_),
    .A(_02223_),
    .B(_02224_));
 sg13g2_xnor2_1 _12588_ (.Y(_02226_),
    .A(_02218_),
    .B(_02225_));
 sg13g2_xor2_1 _12589_ (.B(net2252),
    .A(net2258),
    .X(_02227_));
 sg13g2_xnor2_1 _12590_ (.Y(_02228_),
    .A(net2611),
    .B(net2254));
 sg13g2_xor2_1 _12591_ (.B(net2522),
    .A(net2432),
    .X(_02229_));
 sg13g2_nor2b_1 _12592_ (.A(net2272),
    .B_N(net2594),
    .Y(_02230_));
 sg13g2_xnor2_1 _12593_ (.Y(_02231_),
    .A(_02229_),
    .B(_02230_));
 sg13g2_or2_1 _12594_ (.X(_02232_),
    .B(_02231_),
    .A(_02228_));
 sg13g2_nand2_1 _12595_ (.Y(_02233_),
    .A(_02228_),
    .B(_02231_));
 sg13g2_xnor2_1 _12596_ (.Y(_02234_),
    .A(_02228_),
    .B(_02231_));
 sg13g2_xnor2_1 _12597_ (.Y(_02235_),
    .A(_02227_),
    .B(_02234_));
 sg13g2_xnor2_1 _12598_ (.Y(_02236_),
    .A(net2653),
    .B(net2735));
 sg13g2_xor2_1 _12599_ (.B(net2240),
    .A(net2267),
    .X(_02237_));
 sg13g2_nor2_2 _12600_ (.A(_02236_),
    .B(_02237_),
    .Y(_02238_));
 sg13g2_nor2b_1 _12601_ (.A(net2479),
    .B_N(net2709),
    .Y(_02239_));
 sg13g2_nor3_2 _12602_ (.A(\net.in[35] ),
    .B(net2703),
    .C(_02239_),
    .Y(_02240_));
 sg13g2_xnor2_1 _12603_ (.Y(_02241_),
    .A(net2736),
    .B(net2703));
 sg13g2_nor3_2 _12604_ (.A(net2794),
    .B(net2177),
    .C(_02241_),
    .Y(_02242_));
 sg13g2_nor2b_1 _12605_ (.A(_02240_),
    .B_N(_02242_),
    .Y(_02243_));
 sg13g2_nand2b_1 _12606_ (.Y(_02244_),
    .B(_02240_),
    .A_N(_02242_));
 sg13g2_xor2_1 _12607_ (.B(_02242_),
    .A(_02240_),
    .X(_02245_));
 sg13g2_xnor2_1 _12608_ (.Y(_02246_),
    .A(_02238_),
    .B(_02245_));
 sg13g2_nand2_1 _12609_ (.Y(_02247_),
    .A(_02235_),
    .B(_02246_));
 sg13g2_nor2_1 _12610_ (.A(_02235_),
    .B(_02246_),
    .Y(_02248_));
 sg13g2_xnor2_1 _12611_ (.Y(_02249_),
    .A(_02235_),
    .B(_02246_));
 sg13g2_xnor2_1 _12612_ (.Y(_02250_),
    .A(_02226_),
    .B(_02249_));
 sg13g2_nor2_1 _12613_ (.A(_02215_),
    .B(_02250_),
    .Y(_02251_));
 sg13g2_and2_1 _12614_ (.A(_02215_),
    .B(_02250_),
    .X(_02252_));
 sg13g2_inv_1 _12615_ (.Y(_02253_),
    .A(_02252_));
 sg13g2_nor2_1 _12616_ (.A(_02251_),
    .B(_02252_),
    .Y(_02254_));
 sg13g2_a21oi_1 _12617_ (.A1(_02182_),
    .A2(_02253_),
    .Y(_02255_),
    .B1(_02251_));
 sg13g2_xor2_1 _12618_ (.B(_02254_),
    .A(_02182_),
    .X(_02256_));
 sg13g2_a22oi_1 _12619_ (.Y(_02257_),
    .B1(net2549),
    .B2(net2183),
    .A2(net2178),
    .A1(\net.in[149] ));
 sg13g2_o21ai_1 _12620_ (.B1(_02257_),
    .Y(_02258_),
    .A1(net2183),
    .A2(net2549));
 sg13g2_or2_1 _12621_ (.X(_02259_),
    .B(net2631),
    .A(net2375));
 sg13g2_xnor2_1 _12622_ (.Y(_02260_),
    .A(net2185),
    .B(net2286));
 sg13g2_a22oi_1 _12623_ (.Y(_02261_),
    .B1(_02259_),
    .B2(_02260_),
    .A2(_02058_),
    .A1(net2631));
 sg13g2_nand3_1 _12624_ (.B(_02058_),
    .C(_02260_),
    .A(net2631),
    .Y(_02262_));
 sg13g2_nor2b_1 _12625_ (.A(_02261_),
    .B_N(_02262_),
    .Y(_02263_));
 sg13g2_xnor2_1 _12626_ (.Y(_02264_),
    .A(_02258_),
    .B(_02263_));
 sg13g2_xnor2_1 _12627_ (.Y(_02265_),
    .A(net2680),
    .B(net2603));
 sg13g2_o21ai_1 _12628_ (.B1(_02265_),
    .Y(_02266_),
    .A1(net2223),
    .A2(_06034_));
 sg13g2_nand2b_1 _12629_ (.Y(_02267_),
    .B(net2528),
    .A_N(net2504));
 sg13g2_nor2_1 _12630_ (.A(net2687),
    .B(net2612),
    .Y(_02268_));
 sg13g2_xor2_1 _12631_ (.B(net2236),
    .A(net2385),
    .X(_02269_));
 sg13g2_xnor2_1 _12632_ (.Y(_02270_),
    .A(_02268_),
    .B(_02269_));
 sg13g2_nor2_1 _12633_ (.A(_02267_),
    .B(_02270_),
    .Y(_02271_));
 sg13g2_xnor2_1 _12634_ (.Y(_02272_),
    .A(_02267_),
    .B(_02270_));
 sg13g2_xor2_1 _12635_ (.B(_02272_),
    .A(_02266_),
    .X(_02273_));
 sg13g2_nor2b_1 _12636_ (.A(net2780),
    .B_N(_02194_),
    .Y(_02274_));
 sg13g2_a22oi_1 _12637_ (.Y(_02275_),
    .B1(net2459),
    .B2(\net.in[80] ),
    .A2(_05572_),
    .A1(net2529));
 sg13g2_o21ai_1 _12638_ (.B1(_02275_),
    .Y(_02276_),
    .A1(net2528),
    .A2(_05572_));
 sg13g2_nand2_1 _12639_ (.Y(_02277_),
    .A(_05253_),
    .B(net2733));
 sg13g2_nor2b_1 _12640_ (.A(net2649),
    .B_N(net2719),
    .Y(_02278_));
 sg13g2_xnor2_1 _12641_ (.Y(_02279_),
    .A(_02277_),
    .B(_02278_));
 sg13g2_inv_1 _12642_ (.Y(_02280_),
    .A(_02279_));
 sg13g2_nand2_1 _12643_ (.Y(_02281_),
    .A(_02276_),
    .B(_02280_));
 sg13g2_xnor2_1 _12644_ (.Y(_02282_),
    .A(_02276_),
    .B(_02279_));
 sg13g2_xnor2_1 _12645_ (.Y(_02283_),
    .A(_02274_),
    .B(_02282_));
 sg13g2_nor2_1 _12646_ (.A(_02273_),
    .B(_02283_),
    .Y(_02284_));
 sg13g2_nand2_1 _12647_ (.Y(_02285_),
    .A(_02273_),
    .B(_02283_));
 sg13g2_xor2_1 _12648_ (.B(_02283_),
    .A(_02273_),
    .X(_02286_));
 sg13g2_xnor2_1 _12649_ (.Y(_02287_),
    .A(_02264_),
    .B(_02286_));
 sg13g2_nand2_2 _12650_ (.Y(_02288_),
    .A(_05055_),
    .B(net2412));
 sg13g2_xnor2_1 _12651_ (.Y(_02289_),
    .A(_00005_),
    .B(_02288_));
 sg13g2_xor2_1 _12652_ (.B(net2251),
    .A(net2670),
    .X(_02290_));
 sg13g2_xnor2_1 _12653_ (.Y(_02291_),
    .A(net2297),
    .B(net2202));
 sg13g2_a21oi_1 _12654_ (.A1(_00014_),
    .A2(_02290_),
    .Y(_02292_),
    .B1(_02291_));
 sg13g2_nand3_1 _12655_ (.B(_02290_),
    .C(_02291_),
    .A(_00014_),
    .Y(_02293_));
 sg13g2_nand2b_1 _12656_ (.Y(_02294_),
    .B(_02293_),
    .A_N(_02292_));
 sg13g2_xnor2_1 _12657_ (.Y(_02295_),
    .A(_02289_),
    .B(_02294_));
 sg13g2_xor2_1 _12658_ (.B(\net.in[54] ),
    .A(net2599),
    .X(_02296_));
 sg13g2_xor2_1 _12659_ (.B(\net.in[242] ),
    .A(net2703),
    .X(_02297_));
 sg13g2_xor2_1 _12660_ (.B(net2199),
    .A(net2192),
    .X(_02298_));
 sg13g2_nor2_2 _12661_ (.A(_02297_),
    .B(_02298_),
    .Y(_02299_));
 sg13g2_nor4_2 _12662_ (.A(net2308),
    .B(net2213),
    .C(_05462_),
    .Y(_02300_),
    .D(net2283));
 sg13g2_nor2b_1 _12663_ (.A(_02299_),
    .B_N(_02300_),
    .Y(_02301_));
 sg13g2_nand2b_1 _12664_ (.Y(_02302_),
    .B(_02299_),
    .A_N(_02300_));
 sg13g2_xnor2_1 _12665_ (.Y(_02303_),
    .A(_02299_),
    .B(_02300_));
 sg13g2_xnor2_1 _12666_ (.Y(_02304_),
    .A(_02296_),
    .B(_02303_));
 sg13g2_xnor2_1 _12667_ (.Y(_02305_),
    .A(net2297),
    .B(net2288));
 sg13g2_a21oi_2 _12668_ (.B1(_02305_),
    .Y(_02306_),
    .A2(_05781_),
    .A1(_05374_));
 sg13g2_xor2_1 _12669_ (.B(net2343),
    .A(net2414),
    .X(_02307_));
 sg13g2_nor2_1 _12670_ (.A(net2522),
    .B(net2427),
    .Y(_02308_));
 sg13g2_nor2_1 _12671_ (.A(net2384),
    .B(net2272),
    .Y(_02309_));
 sg13g2_xnor2_1 _12672_ (.Y(_02310_),
    .A(_02308_),
    .B(_02309_));
 sg13g2_xnor2_1 _12673_ (.Y(_02311_),
    .A(_02307_),
    .B(_02310_));
 sg13g2_xnor2_1 _12674_ (.Y(_02312_),
    .A(_02306_),
    .B(_02311_));
 sg13g2_nand2b_1 _12675_ (.Y(_02313_),
    .B(_02312_),
    .A_N(_02304_));
 sg13g2_nand2b_1 _12676_ (.Y(_02314_),
    .B(_02304_),
    .A_N(_02312_));
 sg13g2_xnor2_1 _12677_ (.Y(_02315_),
    .A(_02304_),
    .B(_02312_));
 sg13g2_xnor2_1 _12678_ (.Y(_02316_),
    .A(_02295_),
    .B(_02315_));
 sg13g2_nand2b_1 _12679_ (.Y(_02317_),
    .B(net2566),
    .A_N(net2422));
 sg13g2_xnor2_1 _12680_ (.Y(_02318_),
    .A(net2423),
    .B(net2568));
 sg13g2_xor2_1 _12681_ (.B(net2567),
    .A(\net.in[152] ),
    .X(_02319_));
 sg13g2_xor2_1 _12682_ (.B(net2379),
    .A(net2219),
    .X(_02320_));
 sg13g2_nand2_2 _12683_ (.Y(_02321_),
    .A(net2564),
    .B(_02320_));
 sg13g2_nand2b_1 _12684_ (.Y(_02322_),
    .B(net2385),
    .A_N(net2303));
 sg13g2_nand2b_1 _12685_ (.Y(_02323_),
    .B(net2303),
    .A_N(net2385));
 sg13g2_nand2b_1 _12686_ (.Y(_02324_),
    .B(net2308),
    .A_N(net2236));
 sg13g2_nand3_1 _12687_ (.B(_02323_),
    .C(_02324_),
    .A(_02322_),
    .Y(_02325_));
 sg13g2_or2_1 _12688_ (.X(_02326_),
    .B(_02325_),
    .A(_02321_));
 sg13g2_nand2_1 _12689_ (.Y(_02327_),
    .A(_02321_),
    .B(_02325_));
 sg13g2_nand2_1 _12690_ (.Y(_02328_),
    .A(_02326_),
    .B(_02327_));
 sg13g2_xnor2_1 _12691_ (.Y(_02329_),
    .A(_02318_),
    .B(_02328_));
 sg13g2_o21ai_1 _12692_ (.B1(net2628),
    .Y(_02330_),
    .A1(net2369),
    .A2(net2715));
 sg13g2_xor2_1 _12693_ (.B(net2687),
    .A(net2698),
    .X(_02331_));
 sg13g2_o21ai_1 _12694_ (.B1(_02331_),
    .Y(_02332_),
    .A1(net2785),
    .A2(_02330_));
 sg13g2_nor3_1 _12695_ (.A(net2785),
    .B(_02330_),
    .C(_02331_),
    .Y(_02333_));
 sg13g2_or3_1 _12696_ (.A(net2785),
    .B(_02330_),
    .C(_02331_),
    .X(_02334_));
 sg13g2_and2_1 _12697_ (.A(_02332_),
    .B(_02334_),
    .X(_02335_));
 sg13g2_nor2_1 _12698_ (.A(net2788),
    .B(net2240),
    .Y(_02336_));
 sg13g2_xor2_1 _12699_ (.B(net2574),
    .A(\net.in[55] ),
    .X(_02337_));
 sg13g2_xnor2_1 _12700_ (.Y(_02338_),
    .A(_02336_),
    .B(_02337_));
 sg13g2_xnor2_1 _12701_ (.Y(_02339_),
    .A(_02335_),
    .B(_02338_));
 sg13g2_xor2_1 _12702_ (.B(net2733),
    .A(net2578),
    .X(_02340_));
 sg13g2_nor2_1 _12703_ (.A(net2608),
    .B(net2496),
    .Y(_02341_));
 sg13g2_nand2_1 _12704_ (.Y(_02342_),
    .A(net2339),
    .B(net2715));
 sg13g2_xor2_1 _12705_ (.B(_02342_),
    .A(_02341_),
    .X(_02343_));
 sg13g2_nand2_1 _12706_ (.Y(_02344_),
    .A(_02340_),
    .B(_02343_));
 sg13g2_nor2_1 _12707_ (.A(_02340_),
    .B(_02343_),
    .Y(_02345_));
 sg13g2_xnor2_1 _12708_ (.Y(_02346_),
    .A(_02340_),
    .B(_02343_));
 sg13g2_xor2_1 _12709_ (.B(net2204),
    .A(net2297),
    .X(_02347_));
 sg13g2_xnor2_1 _12710_ (.Y(_02348_),
    .A(_02346_),
    .B(_02347_));
 sg13g2_nand2_1 _12711_ (.Y(_02349_),
    .A(_02339_),
    .B(_02348_));
 sg13g2_nor2_1 _12712_ (.A(_02339_),
    .B(_02348_),
    .Y(_02350_));
 sg13g2_xor2_1 _12713_ (.B(_02348_),
    .A(_02339_),
    .X(_02351_));
 sg13g2_xnor2_1 _12714_ (.Y(_02352_),
    .A(_02329_),
    .B(_02351_));
 sg13g2_nand2b_1 _12715_ (.Y(_02353_),
    .B(_02352_),
    .A_N(_02316_));
 sg13g2_nand2b_1 _12716_ (.Y(_02354_),
    .B(_02316_),
    .A_N(_02352_));
 sg13g2_xor2_1 _12717_ (.B(_02352_),
    .A(_02316_),
    .X(_02355_));
 sg13g2_xnor2_1 _12718_ (.Y(_02356_),
    .A(_02287_),
    .B(_02355_));
 sg13g2_xor2_1 _12719_ (.B(\net.in[237] ),
    .A(net2280),
    .X(_02357_));
 sg13g2_xor2_1 _12720_ (.B(net2208),
    .A(net2266),
    .X(_02358_));
 sg13g2_nor2_1 _12721_ (.A(_02357_),
    .B(_02358_),
    .Y(_02359_));
 sg13g2_nand2b_1 _12722_ (.Y(_02360_),
    .B(\net.in[204] ),
    .A_N(net2185));
 sg13g2_o21ai_1 _12723_ (.B1(_02360_),
    .Y(_02361_),
    .A1(_05286_),
    .A2(net2730));
 sg13g2_a21oi_1 _12724_ (.A1(net2185),
    .A2(_06056_),
    .Y(_02362_),
    .B1(_02361_));
 sg13g2_xor2_1 _12725_ (.B(net2791),
    .A(net2795),
    .X(_02363_));
 sg13g2_nor2b_1 _12726_ (.A(_02363_),
    .B_N(_02362_),
    .Y(_02364_));
 sg13g2_nand2b_1 _12727_ (.Y(_02365_),
    .B(_02363_),
    .A_N(_02362_));
 sg13g2_nor2b_1 _12728_ (.A(_02364_),
    .B_N(_02365_),
    .Y(_02366_));
 sg13g2_xnor2_1 _12729_ (.Y(_02367_),
    .A(_02359_),
    .B(_02366_));
 sg13g2_nor2b_1 _12730_ (.A(net2347),
    .B_N(net2479),
    .Y(_02368_));
 sg13g2_xnor2_1 _12731_ (.Y(_02369_),
    .A(net2391),
    .B(net2538));
 sg13g2_xnor2_1 _12732_ (.Y(_02370_),
    .A(_02368_),
    .B(_02369_));
 sg13g2_nor2b_1 _12733_ (.A(net2408),
    .B_N(net2433),
    .Y(_02371_));
 sg13g2_xor2_1 _12734_ (.B(net2761),
    .A(net2474),
    .X(_02372_));
 sg13g2_nor3_1 _12735_ (.A(net2314),
    .B(_02371_),
    .C(_02372_),
    .Y(_02373_));
 sg13g2_o21ai_1 _12736_ (.B1(_02371_),
    .Y(_02374_),
    .A1(net2314),
    .A2(_02372_));
 sg13g2_nand2b_1 _12737_ (.Y(_02375_),
    .B(_02374_),
    .A_N(_02373_));
 sg13g2_xnor2_1 _12738_ (.Y(_02376_),
    .A(_02370_),
    .B(_02375_));
 sg13g2_nand2b_1 _12739_ (.Y(_02377_),
    .B(net2283),
    .A_N(\net.in[81] ));
 sg13g2_and2_1 _12740_ (.A(_02296_),
    .B(_02377_),
    .X(_02378_));
 sg13g2_nor2b_1 _12741_ (.A(net2733),
    .B_N(net2400),
    .Y(_02379_));
 sg13g2_xnor2_1 _12742_ (.Y(_02380_),
    .A(net2188),
    .B(net2250));
 sg13g2_xnor2_1 _12743_ (.Y(_02381_),
    .A(_02379_),
    .B(_02380_));
 sg13g2_nor2_1 _12744_ (.A(_02229_),
    .B(_02381_),
    .Y(_02382_));
 sg13g2_nand2_1 _12745_ (.Y(_02383_),
    .A(_02229_),
    .B(_02381_));
 sg13g2_xnor2_1 _12746_ (.Y(_02384_),
    .A(_02229_),
    .B(_02381_));
 sg13g2_xnor2_1 _12747_ (.Y(_02385_),
    .A(_02378_),
    .B(_02384_));
 sg13g2_nor2_1 _12748_ (.A(_02376_),
    .B(_02385_),
    .Y(_02386_));
 sg13g2_nand2_1 _12749_ (.Y(_02387_),
    .A(_02376_),
    .B(_02385_));
 sg13g2_nor2b_1 _12750_ (.A(_02386_),
    .B_N(_02387_),
    .Y(_02388_));
 sg13g2_xnor2_1 _12751_ (.Y(_02389_),
    .A(_02367_),
    .B(_02388_));
 sg13g2_xor2_1 _12752_ (.B(net2280),
    .A(net2402),
    .X(_02390_));
 sg13g2_xnor2_1 _12753_ (.Y(_02391_),
    .A(_02016_),
    .B(_02390_));
 sg13g2_xor2_1 _12754_ (.B(net2758),
    .A(net2765),
    .X(_02392_));
 sg13g2_nor2_2 _12755_ (.A(net2313),
    .B(_02392_),
    .Y(_02393_));
 sg13g2_xnor2_1 _12756_ (.Y(_02394_),
    .A(net2474),
    .B(net2386));
 sg13g2_nand2_1 _12757_ (.Y(_02395_),
    .A(net2649),
    .B(_02394_));
 sg13g2_nand3_1 _12758_ (.B(_02393_),
    .C(_02394_),
    .A(net2649),
    .Y(_02396_));
 sg13g2_nor2b_1 _12759_ (.A(_02393_),
    .B_N(_02395_),
    .Y(_02397_));
 sg13g2_xnor2_1 _12760_ (.Y(_02398_),
    .A(_02393_),
    .B(_02395_));
 sg13g2_xnor2_1 _12761_ (.Y(_02399_),
    .A(_02391_),
    .B(_02398_));
 sg13g2_o21ai_1 _12762_ (.B1(net2617),
    .Y(_02400_),
    .A1(net2181),
    .A2(net2459));
 sg13g2_xor2_1 _12763_ (.B(net2236),
    .A(net2267),
    .X(_02401_));
 sg13g2_or3_2 _12764_ (.A(net2242),
    .B(net2213),
    .C(_02401_),
    .X(_02402_));
 sg13g2_nor2_2 _12765_ (.A(\net.in[69] ),
    .B(net2206),
    .Y(_02403_));
 sg13g2_nand2b_1 _12766_ (.Y(_02404_),
    .B(net2522),
    .A_N(net2240));
 sg13g2_xnor2_1 _12767_ (.Y(_02405_),
    .A(_02403_),
    .B(_02404_));
 sg13g2_nor2_1 _12768_ (.A(_02402_),
    .B(_02405_),
    .Y(_02406_));
 sg13g2_xor2_1 _12769_ (.B(_02405_),
    .A(_02402_),
    .X(_02407_));
 sg13g2_xnor2_1 _12770_ (.Y(_02408_),
    .A(_02400_),
    .B(_02407_));
 sg13g2_nor2_1 _12771_ (.A(net2475),
    .B(net2267),
    .Y(_02409_));
 sg13g2_xnor2_1 _12772_ (.Y(_02410_),
    .A(net2385),
    .B(net2744));
 sg13g2_xnor2_1 _12773_ (.Y(_02411_),
    .A(_02409_),
    .B(_02410_));
 sg13g2_nor2b_1 _12774_ (.A(net2250),
    .B_N(net2718),
    .Y(_02412_));
 sg13g2_xnor2_1 _12775_ (.Y(_02413_),
    .A(net2504),
    .B(_02412_));
 sg13g2_nand2b_1 _12776_ (.Y(_02414_),
    .B(net2528),
    .A_N(net2508));
 sg13g2_nor2_1 _12777_ (.A(net2653),
    .B(net2626),
    .Y(_02415_));
 sg13g2_xnor2_1 _12778_ (.Y(_02416_),
    .A(_02414_),
    .B(_02415_));
 sg13g2_nor2_1 _12779_ (.A(_02413_),
    .B(_02416_),
    .Y(_02417_));
 sg13g2_nand2_1 _12780_ (.Y(_02418_),
    .A(_02413_),
    .B(_02416_));
 sg13g2_xor2_1 _12781_ (.B(_02416_),
    .A(_02413_),
    .X(_02419_));
 sg13g2_xnor2_1 _12782_ (.Y(_02420_),
    .A(_02411_),
    .B(_02419_));
 sg13g2_nor2b_1 _12783_ (.A(_02420_),
    .B_N(_02408_),
    .Y(_02421_));
 sg13g2_nand2b_1 _12784_ (.Y(_02422_),
    .B(_02420_),
    .A_N(_02408_));
 sg13g2_xnor2_1 _12785_ (.Y(_02423_),
    .A(_02408_),
    .B(_02420_));
 sg13g2_xnor2_1 _12786_ (.Y(_02424_),
    .A(_02399_),
    .B(_02423_));
 sg13g2_xor2_1 _12787_ (.B(net2272),
    .A(net2308),
    .X(_02425_));
 sg13g2_nand3b_1 _12788_ (.B(net2644),
    .C(_02130_),
    .Y(_02426_),
    .A_N(net2788));
 sg13g2_xor2_1 _12789_ (.B(net2791),
    .A(net2692),
    .X(_02427_));
 sg13g2_xnor2_1 _12790_ (.Y(_02428_),
    .A(net2343),
    .B(net2427));
 sg13g2_nand2_2 _12791_ (.Y(_02429_),
    .A(_02427_),
    .B(_02428_));
 sg13g2_xor2_1 _12792_ (.B(_02429_),
    .A(_02426_),
    .X(_02430_));
 sg13g2_xnor2_1 _12793_ (.Y(_02431_),
    .A(_02425_),
    .B(_02430_));
 sg13g2_xnor2_1 _12794_ (.Y(_02432_),
    .A(net2303),
    .B(net2234));
 sg13g2_nor2b_2 _12795_ (.A(net2278),
    .B_N(_02432_),
    .Y(_02433_));
 sg13g2_xor2_1 _12796_ (.B(net2701),
    .A(net2767),
    .X(_02434_));
 sg13g2_nand2_1 _12797_ (.Y(_02435_),
    .A(_01995_),
    .B(_02434_));
 sg13g2_xor2_1 _12798_ (.B(net2279),
    .A(net2464),
    .X(_02436_));
 sg13g2_xor2_1 _12799_ (.B(net2378),
    .A(net2185),
    .X(_02437_));
 sg13g2_nand2_2 _12800_ (.Y(_02438_),
    .A(_02436_),
    .B(_02437_));
 sg13g2_nand2_1 _12801_ (.Y(_02439_),
    .A(_02435_),
    .B(_02438_));
 sg13g2_xor2_1 _12802_ (.B(_02438_),
    .A(_02435_),
    .X(_02440_));
 sg13g2_xnor2_1 _12803_ (.Y(_02441_),
    .A(_02433_),
    .B(_02440_));
 sg13g2_nor2b_1 _12804_ (.A(net2408),
    .B_N(net2251),
    .Y(_02442_));
 sg13g2_o21ai_1 _12805_ (.B1(_02442_),
    .Y(_02443_),
    .A1(_05396_),
    .A2(\net.in[246] ));
 sg13g2_xor2_1 _12806_ (.B(net2573),
    .A(net2474),
    .X(_02444_));
 sg13g2_xnor2_1 _12807_ (.Y(_02445_),
    .A(net2475),
    .B(net2573));
 sg13g2_nor2_1 _12808_ (.A(net2402),
    .B(\net.in[175] ),
    .Y(_02446_));
 sg13g2_xor2_1 _12809_ (.B(net2440),
    .A(net2528),
    .X(_02447_));
 sg13g2_xnor2_1 _12810_ (.Y(_02448_),
    .A(_02446_),
    .B(_02447_));
 sg13g2_nor2_1 _12811_ (.A(_02444_),
    .B(_02448_),
    .Y(_02449_));
 sg13g2_nand2_1 _12812_ (.Y(_02450_),
    .A(_02444_),
    .B(_02448_));
 sg13g2_xnor2_1 _12813_ (.Y(_02451_),
    .A(_02445_),
    .B(_02448_));
 sg13g2_xnor2_1 _12814_ (.Y(_02452_),
    .A(_02443_),
    .B(_02451_));
 sg13g2_nor2_1 _12815_ (.A(_02441_),
    .B(_02452_),
    .Y(_02453_));
 sg13g2_nand2_1 _12816_ (.Y(_02454_),
    .A(_02441_),
    .B(_02452_));
 sg13g2_xnor2_1 _12817_ (.Y(_02455_),
    .A(_02441_),
    .B(_02452_));
 sg13g2_xor2_1 _12818_ (.B(_02455_),
    .A(_02431_),
    .X(_02456_));
 sg13g2_nor2_1 _12819_ (.A(_02424_),
    .B(_02456_),
    .Y(_02457_));
 sg13g2_xor2_1 _12820_ (.B(_02456_),
    .A(_02424_),
    .X(_02458_));
 sg13g2_xnor2_1 _12821_ (.Y(_02459_),
    .A(_02389_),
    .B(_02458_));
 sg13g2_nor2_1 _12822_ (.A(_02356_),
    .B(_02459_),
    .Y(_02460_));
 sg13g2_nand2_1 _12823_ (.Y(_02461_),
    .A(_02356_),
    .B(_02459_));
 sg13g2_xnor2_1 _12824_ (.Y(_02462_),
    .A(_02356_),
    .B(_02459_));
 sg13g2_xnor2_1 _12825_ (.Y(_02463_),
    .A(_02256_),
    .B(_02462_));
 sg13g2_nand2_2 _12826_ (.Y(_02464_),
    .A(_02147_),
    .B(_02463_));
 sg13g2_or2_1 _12827_ (.X(_02465_),
    .B(_02463_),
    .A(_02147_));
 sg13g2_and2_1 _12828_ (.A(_02464_),
    .B(_02465_),
    .X(_02466_));
 sg13g2_nor2b_1 _12829_ (.A(net2733),
    .B_N(net2324),
    .Y(_02467_));
 sg13g2_xnor2_1 _12830_ (.Y(_02468_),
    .A(net2454),
    .B(net2499));
 sg13g2_xnor2_1 _12831_ (.Y(_02469_),
    .A(net2808),
    .B(net2306));
 sg13g2_nand2_1 _12832_ (.Y(_02470_),
    .A(_02468_),
    .B(_02469_));
 sg13g2_xor2_1 _12833_ (.B(net2489),
    .A(\net.in[133] ),
    .X(_02471_));
 sg13g2_nand3_1 _12834_ (.B(_05836_),
    .C(_02471_),
    .A(_05737_),
    .Y(_02472_));
 sg13g2_nand2b_1 _12835_ (.Y(_02473_),
    .B(_02470_),
    .A_N(_02472_));
 sg13g2_nand2b_1 _12836_ (.Y(_02474_),
    .B(_02472_),
    .A_N(_02470_));
 sg13g2_xor2_1 _12837_ (.B(_02472_),
    .A(_02470_),
    .X(_02475_));
 sg13g2_xnor2_1 _12838_ (.Y(_02476_),
    .A(_02467_),
    .B(_02475_));
 sg13g2_xnor2_1 _12839_ (.Y(_02477_),
    .A(net2201),
    .B(net2275));
 sg13g2_nand3_1 _12840_ (.B(_05396_),
    .C(_02477_),
    .A(net2339),
    .Y(_02478_));
 sg13g2_nor2_1 _12841_ (.A(\net.in[22] ),
    .B(net2735),
    .Y(_02479_));
 sg13g2_nor2_1 _12842_ (.A(net2228),
    .B(net2758),
    .Y(_02480_));
 sg13g2_a21oi_2 _12843_ (.B1(net2761),
    .Y(_02481_),
    .A2(net2605),
    .A1(\net.in[133] ));
 sg13g2_o21ai_1 _12844_ (.B1(_02481_),
    .Y(_02482_),
    .A1(_02479_),
    .A2(_02480_));
 sg13g2_or3_1 _12845_ (.A(_02479_),
    .B(_02480_),
    .C(_02481_),
    .X(_02483_));
 sg13g2_a21o_1 _12846_ (.A2(_02483_),
    .A1(_02482_),
    .B1(_02478_),
    .X(_02484_));
 sg13g2_nand3_1 _12847_ (.B(_02482_),
    .C(_02483_),
    .A(_02478_),
    .Y(_02485_));
 sg13g2_nor3_2 _12848_ (.A(\net.in[229] ),
    .B(net2667),
    .C(_06089_),
    .Y(_02486_));
 sg13g2_xor2_1 _12849_ (.B(net2497),
    .A(net2533),
    .X(_02487_));
 sg13g2_xnor2_1 _12850_ (.Y(_02488_),
    .A(net2227),
    .B(net2195));
 sg13g2_nor2b_1 _12851_ (.A(net2560),
    .B_N(net2256),
    .Y(_02489_));
 sg13g2_nor2b_1 _12852_ (.A(\net.in[23] ),
    .B_N(net2348),
    .Y(_02490_));
 sg13g2_and4_2 _12853_ (.A(_02487_),
    .B(_02488_),
    .C(_02489_),
    .D(_02490_),
    .X(_02491_));
 sg13g2_a22oi_1 _12854_ (.Y(_02492_),
    .B1(_02489_),
    .B2(_02490_),
    .A2(_02488_),
    .A1(_02487_));
 sg13g2_o21ai_1 _12855_ (.B1(_02486_),
    .Y(_02493_),
    .A1(_02491_),
    .A2(_02492_));
 sg13g2_or3_1 _12856_ (.A(_02486_),
    .B(_02491_),
    .C(_02492_),
    .X(_02494_));
 sg13g2_nand4_1 _12857_ (.B(_02485_),
    .C(_02493_),
    .A(_02484_),
    .Y(_02495_),
    .D(_02494_));
 sg13g2_or2_1 _12858_ (.X(_02496_),
    .B(_02495_),
    .A(_02476_));
 sg13g2_a22oi_1 _12859_ (.Y(_02497_),
    .B1(_02493_),
    .B2(_02494_),
    .A2(_02485_),
    .A1(_02484_));
 sg13g2_nand2_1 _12860_ (.Y(_02498_),
    .A(_02476_),
    .B(_02495_));
 sg13g2_o21ai_1 _12861_ (.B1(_02495_),
    .Y(_02499_),
    .A1(_02476_),
    .A2(_02497_));
 sg13g2_nand2b_1 _12862_ (.Y(_02500_),
    .B(_02498_),
    .A_N(_02497_));
 sg13g2_a22oi_1 _12863_ (.Y(_02501_),
    .B1(_02499_),
    .B2(_02496_),
    .A2(_02497_),
    .A1(_02476_));
 sg13g2_o21ai_1 _12864_ (.B1(_02489_),
    .Y(_02502_),
    .A1(net2557),
    .A2(_05660_));
 sg13g2_a21o_1 _12865_ (.A2(_05660_),
    .A1(net2557),
    .B1(_02502_),
    .X(_02503_));
 sg13g2_xor2_1 _12866_ (.B(net2627),
    .A(net2557),
    .X(_02504_));
 sg13g2_xnor2_1 _12867_ (.Y(_02505_),
    .A(net2557),
    .B(net2628));
 sg13g2_xor2_1 _12868_ (.B(net2239),
    .A(net2707),
    .X(_02506_));
 sg13g2_xor2_1 _12869_ (.B(net2678),
    .A(\net.in[43] ),
    .X(_02507_));
 sg13g2_xnor2_1 _12870_ (.Y(_02508_),
    .A(_02506_),
    .B(_02507_));
 sg13g2_nand2_1 _12871_ (.Y(_02509_),
    .A(_02505_),
    .B(_02508_));
 sg13g2_nor2_1 _12872_ (.A(_02505_),
    .B(_02508_),
    .Y(_02510_));
 sg13g2_xnor2_1 _12873_ (.Y(_02511_),
    .A(_02505_),
    .B(_02508_));
 sg13g2_xnor2_1 _12874_ (.Y(_02512_),
    .A(_02503_),
    .B(_02511_));
 sg13g2_nand2b_1 _12875_ (.Y(_02513_),
    .B(net2347),
    .A_N(net2735));
 sg13g2_nor2_1 _12876_ (.A(net2184),
    .B(net2795),
    .Y(_02514_));
 sg13g2_xnor2_1 _12877_ (.Y(_02515_),
    .A(_02513_),
    .B(_02514_));
 sg13g2_or2_1 _12878_ (.X(_02516_),
    .B(net2398),
    .A(net2392));
 sg13g2_xor2_1 _12879_ (.B(net2400),
    .A(net2391),
    .X(_02517_));
 sg13g2_o21ai_1 _12880_ (.B1(_02517_),
    .Y(_02518_),
    .A1(net2283),
    .A2(net2459));
 sg13g2_nor2_1 _12881_ (.A(net2497),
    .B(net2713),
    .Y(_02519_));
 sg13g2_nor2_1 _12882_ (.A(net2454),
    .B(net2459),
    .Y(_02520_));
 sg13g2_xor2_1 _12883_ (.B(_02520_),
    .A(_02519_),
    .X(_02521_));
 sg13g2_nand2b_1 _12884_ (.Y(_02522_),
    .B(_02521_),
    .A_N(_02518_));
 sg13g2_nor2b_1 _12885_ (.A(_02521_),
    .B_N(_02518_),
    .Y(_02523_));
 sg13g2_xor2_1 _12886_ (.B(_02521_),
    .A(_02518_),
    .X(_02524_));
 sg13g2_o21ai_1 _12887_ (.B1(_02522_),
    .Y(_02525_),
    .A1(_02515_),
    .A2(_02523_));
 sg13g2_xnor2_1 _12888_ (.Y(_02526_),
    .A(_02515_),
    .B(_02524_));
 sg13g2_or2_1 _12889_ (.X(_02527_),
    .B(_02526_),
    .A(_02512_));
 sg13g2_xor2_1 _12890_ (.B(_02526_),
    .A(_02512_),
    .X(_02528_));
 sg13g2_nor2_1 _12891_ (.A(net2258),
    .B(net2815),
    .Y(_02529_));
 sg13g2_a21o_1 _12892_ (.A2(net2815),
    .A1(net2258),
    .B1(net2180),
    .X(_02530_));
 sg13g2_nor3_1 _12893_ (.A(net2661),
    .B(_02529_),
    .C(_02530_),
    .Y(_02531_));
 sg13g2_xnor2_1 _12894_ (.Y(_02532_),
    .A(net2431),
    .B(net2497));
 sg13g2_nor4_1 _12895_ (.A(net2661),
    .B(_02529_),
    .C(_02530_),
    .D(_02532_),
    .Y(_02533_));
 sg13g2_nand2b_1 _12896_ (.Y(_02534_),
    .B(_02532_),
    .A_N(_02531_));
 sg13g2_xnor2_1 _12897_ (.Y(_02535_),
    .A(_02531_),
    .B(_02532_));
 sg13g2_nand2b_1 _12898_ (.Y(_02536_),
    .B(net2467),
    .A_N(net2218));
 sg13g2_nand2_1 _12899_ (.Y(_02537_),
    .A(net2329),
    .B(_05847_));
 sg13g2_xnor2_1 _12900_ (.Y(_02538_),
    .A(_02536_),
    .B(_02537_));
 sg13g2_xnor2_1 _12901_ (.Y(_02539_),
    .A(_02535_),
    .B(_02538_));
 sg13g2_xnor2_1 _12902_ (.Y(_02540_),
    .A(_02528_),
    .B(_02539_));
 sg13g2_nand2b_1 _12903_ (.Y(_02541_),
    .B(_02501_),
    .A_N(_02540_));
 sg13g2_nand2b_1 _12904_ (.Y(_02542_),
    .B(_02540_),
    .A_N(_02501_));
 sg13g2_xnor2_1 _12905_ (.Y(_02543_),
    .A(_02501_),
    .B(_02540_));
 sg13g2_nor2_1 _12906_ (.A(net2621),
    .B(net2546),
    .Y(_02544_));
 sg13g2_nor2b_1 _12907_ (.A(net2767),
    .B_N(net2538),
    .Y(_02545_));
 sg13g2_xnor2_1 _12908_ (.Y(_02546_),
    .A(_02544_),
    .B(_02545_));
 sg13g2_inv_1 _12909_ (.Y(_02547_),
    .A(_02546_));
 sg13g2_xnor2_1 _12910_ (.Y(_02548_),
    .A(net2673),
    .B(net2667));
 sg13g2_xnor2_1 _12911_ (.Y(_02549_),
    .A(net2678),
    .B(net2779));
 sg13g2_nand2_1 _12912_ (.Y(_02550_),
    .A(_02548_),
    .B(_02549_));
 sg13g2_xnor2_1 _12913_ (.Y(_02551_),
    .A(net2617),
    .B(net2607));
 sg13g2_xnor2_1 _12914_ (.Y(_02552_),
    .A(_00010_),
    .B(_02551_));
 sg13g2_nand2b_1 _12915_ (.Y(_02553_),
    .B(_02552_),
    .A_N(_02550_));
 sg13g2_a21oi_1 _12916_ (.A1(_02548_),
    .A2(_02549_),
    .Y(_02554_),
    .B1(_02552_));
 sg13g2_xnor2_1 _12917_ (.Y(_02555_),
    .A(_02550_),
    .B(_02552_));
 sg13g2_xnor2_1 _12918_ (.Y(_02556_),
    .A(_02546_),
    .B(_02555_));
 sg13g2_a21oi_2 _12919_ (.B1(_01233_),
    .Y(_02557_),
    .A2(_05726_),
    .A1(net2233));
 sg13g2_xor2_1 _12920_ (.B(net2442),
    .A(net2434),
    .X(_02558_));
 sg13g2_xnor2_1 _12921_ (.Y(_02559_),
    .A(net2436),
    .B(net2443));
 sg13g2_xnor2_1 _12922_ (.Y(_02560_),
    .A(net2257),
    .B(net2795));
 sg13g2_nor3_1 _12923_ (.A(net2657),
    .B(_02559_),
    .C(_02560_),
    .Y(_02561_));
 sg13g2_o21ai_1 _12924_ (.B1(_02560_),
    .Y(_02562_),
    .A1(net2657),
    .A2(_02559_));
 sg13g2_nor2b_1 _12925_ (.A(_02561_),
    .B_N(_02562_),
    .Y(_02563_));
 sg13g2_xnor2_1 _12926_ (.Y(_02564_),
    .A(_02557_),
    .B(_02563_));
 sg13g2_or2_1 _12927_ (.X(_02565_),
    .B(_02564_),
    .A(_02556_));
 sg13g2_xnor2_1 _12928_ (.Y(_02566_),
    .A(_02556_),
    .B(_02564_));
 sg13g2_nor2b_1 _12929_ (.A(net2663),
    .B_N(net2344),
    .Y(_02567_));
 sg13g2_nor2b_1 _12930_ (.A(net2192),
    .B_N(net2713),
    .Y(_02568_));
 sg13g2_nor2_1 _12931_ (.A(_05396_),
    .B(net2713),
    .Y(_02569_));
 sg13g2_nor2_1 _12932_ (.A(net2386),
    .B(net2490),
    .Y(_02570_));
 sg13g2_nor3_2 _12933_ (.A(_02568_),
    .B(_02569_),
    .C(_02570_),
    .Y(_02571_));
 sg13g2_nand2_1 _12934_ (.Y(_02572_),
    .A(net2384),
    .B(net2330));
 sg13g2_nand2_1 _12935_ (.Y(_02573_),
    .A(_05044_),
    .B(net2693));
 sg13g2_xnor2_1 _12936_ (.Y(_02574_),
    .A(_02572_),
    .B(_02573_));
 sg13g2_inv_1 _12937_ (.Y(_02575_),
    .A(_02574_));
 sg13g2_nand2_1 _12938_ (.Y(_02576_),
    .A(_02571_),
    .B(_02575_));
 sg13g2_xnor2_1 _12939_ (.Y(_02577_),
    .A(_02571_),
    .B(_02574_));
 sg13g2_xnor2_1 _12940_ (.Y(_02578_),
    .A(_02567_),
    .B(_02577_));
 sg13g2_xnor2_1 _12941_ (.Y(_02579_),
    .A(_02566_),
    .B(_02578_));
 sg13g2_xnor2_1 _12942_ (.Y(_02580_),
    .A(_02543_),
    .B(_02579_));
 sg13g2_nor2b_1 _12943_ (.A(net2229),
    .B_N(net2635),
    .Y(_02581_));
 sg13g2_nor2b_1 _12944_ (.A(net2635),
    .B_N(net2226),
    .Y(_02582_));
 sg13g2_nor2b_1 _12945_ (.A(net2335),
    .B_N(net2506),
    .Y(_02583_));
 sg13g2_nor3_2 _12946_ (.A(_02581_),
    .B(_02582_),
    .C(_02583_),
    .Y(_02584_));
 sg13g2_nor2_2 _12947_ (.A(_00439_),
    .B(_02584_),
    .Y(_02585_));
 sg13g2_xnor2_1 _12948_ (.Y(_02586_),
    .A(_00435_),
    .B(_02584_));
 sg13g2_nor2_1 _12949_ (.A(net2380),
    .B(net2489),
    .Y(_02587_));
 sg13g2_xor2_1 _12950_ (.B(\net.in[237] ),
    .A(net2195),
    .X(_02588_));
 sg13g2_xnor2_1 _12951_ (.Y(_02589_),
    .A(_02587_),
    .B(_02588_));
 sg13g2_a21oi_2 _12952_ (.B1(_02589_),
    .Y(_02590_),
    .A2(_02584_),
    .A1(_00439_));
 sg13g2_xnor2_1 _12953_ (.Y(_02591_),
    .A(_02586_),
    .B(_02589_));
 sg13g2_nor2b_2 _12954_ (.A(net2805),
    .B_N(net2681),
    .Y(_02592_));
 sg13g2_xnor2_1 _12955_ (.Y(_02593_),
    .A(net2750),
    .B(_02592_));
 sg13g2_xnor2_1 _12956_ (.Y(_02594_),
    .A(net2572),
    .B(net2675));
 sg13g2_nor2_1 _12957_ (.A(net2807),
    .B(_02594_),
    .Y(_02595_));
 sg13g2_nor2b_1 _12958_ (.A(net2793),
    .B_N(net2732),
    .Y(_02596_));
 sg13g2_nor2b_1 _12959_ (.A(net2732),
    .B_N(net2793),
    .Y(_02597_));
 sg13g2_nor2_2 _12960_ (.A(net2329),
    .B(net2321),
    .Y(_02598_));
 sg13g2_nor3_2 _12961_ (.A(_02596_),
    .B(_02597_),
    .C(_02598_),
    .Y(_02599_));
 sg13g2_nand2b_1 _12962_ (.Y(_02600_),
    .B(_02595_),
    .A_N(_02599_));
 sg13g2_nor2b_1 _12963_ (.A(_02595_),
    .B_N(_02599_),
    .Y(_02601_));
 sg13g2_xnor2_1 _12964_ (.Y(_02602_),
    .A(_02595_),
    .B(_02599_));
 sg13g2_a21oi_1 _12965_ (.A1(_02593_),
    .A2(_02600_),
    .Y(_02603_),
    .B1(_02601_));
 sg13g2_inv_1 _12966_ (.Y(_02604_),
    .A(_02603_));
 sg13g2_xnor2_1 _12967_ (.Y(_02605_),
    .A(_02593_),
    .B(_02602_));
 sg13g2_nor2_1 _12968_ (.A(_02591_),
    .B(_02605_),
    .Y(_02606_));
 sg13g2_nand2_1 _12969_ (.Y(_02607_),
    .A(_02591_),
    .B(_02605_));
 sg13g2_xor2_1 _12970_ (.B(_02605_),
    .A(_02591_),
    .X(_02608_));
 sg13g2_xor2_1 _12971_ (.B(\net.in[29] ),
    .A(\net.in[11] ),
    .X(_02609_));
 sg13g2_nand2_1 _12972_ (.Y(_02610_),
    .A(_05099_),
    .B(_02609_));
 sg13g2_o21ai_1 _12973_ (.B1(_02610_),
    .Y(_02611_),
    .A1(_05099_),
    .A2(\net.in[29] ));
 sg13g2_xnor2_1 _12974_ (.Y(_02612_),
    .A(net2499),
    .B(net2481));
 sg13g2_xnor2_1 _12975_ (.Y(_02613_),
    .A(net2652),
    .B(net2768));
 sg13g2_xor2_1 _12976_ (.B(net2202),
    .A(net2609),
    .X(_02614_));
 sg13g2_xnor2_1 _12977_ (.Y(_02615_),
    .A(_02613_),
    .B(_02614_));
 sg13g2_nor2_1 _12978_ (.A(_02612_),
    .B(_02615_),
    .Y(_02616_));
 sg13g2_nand2_1 _12979_ (.Y(_02617_),
    .A(_02612_),
    .B(_02615_));
 sg13g2_nor2b_1 _12980_ (.A(_02616_),
    .B_N(_02617_),
    .Y(_02618_));
 sg13g2_a21oi_2 _12981_ (.B1(_02616_),
    .Y(_02619_),
    .A2(_02617_),
    .A1(_02611_));
 sg13g2_xor2_1 _12982_ (.B(_02618_),
    .A(_02611_),
    .X(_02620_));
 sg13g2_xnor2_1 _12983_ (.Y(_02621_),
    .A(_02608_),
    .B(_02620_));
 sg13g2_xor2_1 _12984_ (.B(net2256),
    .A(net2292),
    .X(_02622_));
 sg13g2_nor2_1 _12985_ (.A(net2187),
    .B(net2674),
    .Y(_02623_));
 sg13g2_xor2_1 _12986_ (.B(net2271),
    .A(net2669),
    .X(_02624_));
 sg13g2_xnor2_1 _12987_ (.Y(_02625_),
    .A(_02623_),
    .B(_02624_));
 sg13g2_nor2b_1 _12988_ (.A(_02625_),
    .B_N(_02622_),
    .Y(_02626_));
 sg13g2_nor2b_1 _12989_ (.A(_02622_),
    .B_N(_02625_),
    .Y(_02627_));
 sg13g2_xnor2_1 _12990_ (.Y(_02628_),
    .A(_02622_),
    .B(_02625_));
 sg13g2_nor2_1 _12991_ (.A(net2184),
    .B(net2674),
    .Y(_02629_));
 sg13g2_nor2b_2 _12992_ (.A(net2450),
    .B_N(net2645),
    .Y(_02630_));
 sg13g2_xnor2_1 _12993_ (.Y(_02631_),
    .A(_02629_),
    .B(_02630_));
 sg13g2_xnor2_1 _12994_ (.Y(_02632_),
    .A(_02628_),
    .B(_02631_));
 sg13g2_nor2_1 _12995_ (.A(net2629),
    .B(net2669),
    .Y(_02633_));
 sg13g2_xor2_1 _12996_ (.B(\net.in[31] ),
    .A(net2662),
    .X(_02634_));
 sg13g2_xnor2_1 _12997_ (.Y(_02635_),
    .A(_02633_),
    .B(_02634_));
 sg13g2_nor2_1 _12998_ (.A(net2300),
    .B(net2355),
    .Y(_02636_));
 sg13g2_nor2_1 _12999_ (.A(net2485),
    .B(\net.in[10] ),
    .Y(_02637_));
 sg13g2_xnor2_1 _13000_ (.Y(_02638_),
    .A(net2493),
    .B(net2438));
 sg13g2_o21ai_1 _13001_ (.B1(_02638_),
    .Y(_02639_),
    .A1(_02636_),
    .A2(_02637_));
 sg13g2_or3_1 _13002_ (.A(_02636_),
    .B(_02637_),
    .C(_02638_),
    .X(_02640_));
 sg13g2_nand2_1 _13003_ (.Y(_02641_),
    .A(_02639_),
    .B(_02640_));
 sg13g2_nand2_1 _13004_ (.Y(_02642_),
    .A(_02635_),
    .B(_02640_));
 sg13g2_nand2_1 _13005_ (.Y(_02643_),
    .A(_02639_),
    .B(_02642_));
 sg13g2_inv_1 _13006_ (.Y(_02644_),
    .A(_02643_));
 sg13g2_xnor2_1 _13007_ (.Y(_02645_),
    .A(_02635_),
    .B(_02641_));
 sg13g2_xnor2_1 _13008_ (.Y(_02646_),
    .A(_02632_),
    .B(_02645_));
 sg13g2_or2_2 _13009_ (.X(_02647_),
    .B(net2435),
    .A(net2526));
 sg13g2_nand2_1 _13010_ (.Y(_02648_),
    .A(net2526),
    .B(net2435));
 sg13g2_xor2_1 _13011_ (.B(net2714),
    .A(net2190),
    .X(_02649_));
 sg13g2_a21o_1 _13012_ (.A2(_02648_),
    .A1(_02647_),
    .B1(_02649_),
    .X(_02650_));
 sg13g2_xor2_1 _13013_ (.B(net2489),
    .A(net2373),
    .X(_02651_));
 sg13g2_xnor2_1 _13014_ (.Y(_02652_),
    .A(net2742),
    .B(net2669));
 sg13g2_nand2_1 _13015_ (.Y(_02653_),
    .A(_02651_),
    .B(_02652_));
 sg13g2_nor2_1 _13016_ (.A(net2555),
    .B(net2458),
    .Y(_02654_));
 sg13g2_nor2b_1 _13017_ (.A(net2238),
    .B_N(net2711),
    .Y(_02655_));
 sg13g2_xnor2_1 _13018_ (.Y(_02656_),
    .A(_02654_),
    .B(_02655_));
 sg13g2_nand2b_1 _13019_ (.Y(_02657_),
    .B(_02656_),
    .A_N(_02653_));
 sg13g2_a21oi_1 _13020_ (.A1(_02651_),
    .A2(_02652_),
    .Y(_02658_),
    .B1(_02656_));
 sg13g2_xnor2_1 _13021_ (.Y(_02659_),
    .A(_02653_),
    .B(_02656_));
 sg13g2_xor2_1 _13022_ (.B(_02659_),
    .A(_02650_),
    .X(_02660_));
 sg13g2_xnor2_1 _13023_ (.Y(_02661_),
    .A(_02646_),
    .B(_02660_));
 sg13g2_nand2_1 _13024_ (.Y(_02662_),
    .A(_02621_),
    .B(_02661_));
 sg13g2_xor2_1 _13025_ (.B(_02661_),
    .A(_02621_),
    .X(_02663_));
 sg13g2_nand2b_1 _13026_ (.Y(_02664_),
    .B(net2275),
    .A_N(net2198));
 sg13g2_o21ai_1 _13027_ (.B1(_02664_),
    .Y(_02665_),
    .A1(net2368),
    .A2(net2362));
 sg13g2_a21oi_2 _13028_ (.B1(_02665_),
    .Y(_02666_),
    .A2(net2198),
    .A1(_05935_));
 sg13g2_o21ai_1 _13029_ (.B1(_02516_),
    .Y(_02667_),
    .A1(net2296),
    .A2(net2321));
 sg13g2_xor2_1 _13030_ (.B(net2485),
    .A(net2431),
    .X(_02668_));
 sg13g2_nand2_1 _13031_ (.Y(_02669_),
    .A(_02548_),
    .B(_02668_));
 sg13g2_nand2_1 _13032_ (.Y(_02670_),
    .A(_02667_),
    .B(_02669_));
 sg13g2_xor2_1 _13033_ (.B(_02669_),
    .A(_02667_),
    .X(_02671_));
 sg13g2_xnor2_1 _13034_ (.Y(_02672_),
    .A(_02666_),
    .B(_02671_));
 sg13g2_nand2_1 _13035_ (.Y(_02673_),
    .A(_05715_),
    .B(_05946_));
 sg13g2_o21ai_1 _13036_ (.B1(_02673_),
    .Y(_02674_),
    .A1(net2759),
    .A2(net2645));
 sg13g2_or2_1 _13037_ (.X(_02675_),
    .B(net2394),
    .A(net2340));
 sg13g2_o21ai_1 _13038_ (.B1(_02675_),
    .Y(_02676_),
    .A1(net2526),
    .A2(_05979_));
 sg13g2_and2_1 _13039_ (.A(net2742),
    .B(net2622),
    .X(_02677_));
 sg13g2_nor2_1 _13040_ (.A(net2741),
    .B(net2622),
    .Y(_02678_));
 sg13g2_nor2b_1 _13041_ (.A(net2559),
    .B_N(net2392),
    .Y(_02679_));
 sg13g2_nor3_2 _13042_ (.A(_02677_),
    .B(_02678_),
    .C(_02679_),
    .Y(_02680_));
 sg13g2_nor2_1 _13043_ (.A(_02676_),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_nand2_1 _13044_ (.Y(_02682_),
    .A(_02676_),
    .B(_02680_));
 sg13g2_xor2_1 _13045_ (.B(_02680_),
    .A(_02676_),
    .X(_02683_));
 sg13g2_xnor2_1 _13046_ (.Y(_02684_),
    .A(_02674_),
    .B(_02683_));
 sg13g2_nand2_1 _13047_ (.Y(_02685_),
    .A(_02672_),
    .B(_02684_));
 sg13g2_or2_1 _13048_ (.X(_02686_),
    .B(_02684_),
    .A(_02672_));
 sg13g2_nand2_1 _13049_ (.Y(_02687_),
    .A(_02685_),
    .B(_02686_));
 sg13g2_xnor2_1 _13050_ (.Y(_02688_),
    .A(net2435),
    .B(net2447));
 sg13g2_nor2_1 _13051_ (.A(net2660),
    .B(net2197),
    .Y(_02689_));
 sg13g2_nor2b_1 _13052_ (.A(\net.in[246] ),
    .B_N(net2344),
    .Y(_02690_));
 sg13g2_xnor2_1 _13053_ (.Y(_02691_),
    .A(\net.in[10] ),
    .B(net2774));
 sg13g2_xnor2_1 _13054_ (.Y(_02692_),
    .A(net2324),
    .B(net2217));
 sg13g2_nand2_1 _13055_ (.Y(_02693_),
    .A(_02691_),
    .B(_02692_));
 sg13g2_and3_1 _13056_ (.X(_02694_),
    .A(_02689_),
    .B(_02690_),
    .C(_02693_));
 sg13g2_a21oi_2 _13057_ (.B1(_02693_),
    .Y(_02695_),
    .A2(_02690_),
    .A1(_02689_));
 sg13g2_or2_1 _13058_ (.X(_02696_),
    .B(_02695_),
    .A(_02694_));
 sg13g2_xnor2_1 _13059_ (.Y(_02697_),
    .A(_02688_),
    .B(_02696_));
 sg13g2_xnor2_1 _13060_ (.Y(_02698_),
    .A(_02687_),
    .B(_02697_));
 sg13g2_xnor2_1 _13061_ (.Y(_02699_),
    .A(_02663_),
    .B(_02698_));
 sg13g2_o21ai_1 _13062_ (.B1(net2255),
    .Y(_02700_),
    .A1(net2300),
    .A2(net2179));
 sg13g2_nor2_2 _13063_ (.A(net2231),
    .B(_02700_),
    .Y(_02701_));
 sg13g2_xnor2_1 _13064_ (.Y(_02702_),
    .A(net2477),
    .B(net2422));
 sg13g2_xor2_1 _13065_ (.B(net2619),
    .A(net2610),
    .X(_02703_));
 sg13g2_xnor2_1 _13066_ (.Y(_02704_),
    .A(net2610),
    .B(net2620));
 sg13g2_xor2_1 _13067_ (.B(net2715),
    .A(net2630),
    .X(_02705_));
 sg13g2_nor3_1 _13068_ (.A(_02702_),
    .B(_02703_),
    .C(_02705_),
    .Y(_02706_));
 sg13g2_o21ai_1 _13069_ (.B1(_02702_),
    .Y(_02707_),
    .A1(_02703_),
    .A2(_02705_));
 sg13g2_nand2b_1 _13070_ (.Y(_02708_),
    .B(_02707_),
    .A_N(_02706_));
 sg13g2_xnor2_1 _13071_ (.Y(_02709_),
    .A(_02701_),
    .B(_02708_));
 sg13g2_nor4_2 _13072_ (.A(net2204),
    .B(net2660),
    .C(\net.in[237] ),
    .Y(_02710_),
    .D(net2274));
 sg13g2_xnor2_1 _13073_ (.Y(_02711_),
    .A(net2717),
    .B(net2776));
 sg13g2_and2_2 _13074_ (.A(_07596_),
    .B(_02711_),
    .X(_02712_));
 sg13g2_xor2_1 _13075_ (.B(net2726),
    .A(net2576),
    .X(_02713_));
 sg13g2_xor2_1 _13076_ (.B(net2714),
    .A(net2194),
    .X(_02714_));
 sg13g2_xnor2_1 _13077_ (.Y(_02715_),
    .A(_02713_),
    .B(_02714_));
 sg13g2_nor2_1 _13078_ (.A(_02712_),
    .B(_02715_),
    .Y(_02716_));
 sg13g2_xor2_1 _13079_ (.B(_02715_),
    .A(_02712_),
    .X(_02717_));
 sg13g2_xnor2_1 _13080_ (.Y(_02718_),
    .A(_02710_),
    .B(_02717_));
 sg13g2_a22oi_1 _13081_ (.Y(_02719_),
    .B1(net2323),
    .B2(net2380),
    .A2(net2805),
    .A1(net2524));
 sg13g2_o21ai_1 _13082_ (.B1(_02719_),
    .Y(_02720_),
    .A1(net2521),
    .A2(net2805));
 sg13g2_nor2_1 _13083_ (.A(net2814),
    .B(net2813),
    .Y(_02721_));
 sg13g2_nor2b_1 _13084_ (.A(net2764),
    .B_N(net2321),
    .Y(_02722_));
 sg13g2_xnor2_1 _13085_ (.Y(_02723_),
    .A(_02721_),
    .B(_02722_));
 sg13g2_nand2_1 _13086_ (.Y(_02724_),
    .A(_02720_),
    .B(_02723_));
 sg13g2_nor2_1 _13087_ (.A(_02720_),
    .B(_02723_),
    .Y(_02725_));
 sg13g2_xnor2_1 _13088_ (.Y(_02726_),
    .A(_02720_),
    .B(_02723_));
 sg13g2_nor2_1 _13089_ (.A(net2184),
    .B(net2737),
    .Y(_02727_));
 sg13g2_nor2_1 _13090_ (.A(_05231_),
    .B(net2774),
    .Y(_02728_));
 sg13g2_xnor2_1 _13091_ (.Y(_02729_),
    .A(_02727_),
    .B(_02728_));
 sg13g2_xnor2_1 _13092_ (.Y(_02730_),
    .A(_02726_),
    .B(_02729_));
 sg13g2_nand2_1 _13093_ (.Y(_02731_),
    .A(_02718_),
    .B(_02730_));
 sg13g2_nor2_1 _13094_ (.A(_02718_),
    .B(_02730_),
    .Y(_02732_));
 sg13g2_xnor2_1 _13095_ (.Y(_02733_),
    .A(_02718_),
    .B(_02730_));
 sg13g2_o21ai_1 _13096_ (.B1(_02731_),
    .Y(_02734_),
    .A1(_02709_),
    .A2(_02732_));
 sg13g2_xnor2_1 _13097_ (.Y(_02735_),
    .A(_02709_),
    .B(_02733_));
 sg13g2_xnor2_1 _13098_ (.Y(_02736_),
    .A(net2733),
    .B(net2647));
 sg13g2_o21ai_1 _13099_ (.B1(_02736_),
    .Y(_02737_),
    .A1(net2295),
    .A2(net2352));
 sg13g2_o21ai_1 _13100_ (.B1(_02704_),
    .Y(_02738_),
    .A1(_05726_),
    .A2(net2803));
 sg13g2_xnor2_1 _13101_ (.Y(_02739_),
    .A(net2630),
    .B(net2767));
 sg13g2_nand2_1 _13102_ (.Y(_02740_),
    .A(_02548_),
    .B(_02739_));
 sg13g2_or2_1 _13103_ (.X(_02741_),
    .B(_02740_),
    .A(_02738_));
 sg13g2_and2_1 _13104_ (.A(_02738_),
    .B(_02740_),
    .X(_02742_));
 sg13g2_xor2_1 _13105_ (.B(_02740_),
    .A(_02738_),
    .X(_02743_));
 sg13g2_xnor2_1 _13106_ (.Y(_02744_),
    .A(_02737_),
    .B(_02743_));
 sg13g2_nor2_1 _13107_ (.A(_05770_),
    .B(net2552),
    .Y(_02745_));
 sg13g2_nor2_2 _13108_ (.A(net2340),
    .B(net2438),
    .Y(_02746_));
 sg13g2_a21oi_1 _13109_ (.A1(_05770_),
    .A2(net2552),
    .Y(_02747_),
    .B1(_02746_));
 sg13g2_nor2b_2 _13110_ (.A(_02745_),
    .B_N(_02747_),
    .Y(_02748_));
 sg13g2_xnor2_1 _13111_ (.Y(_02749_),
    .A(net2765),
    .B(net2696));
 sg13g2_xnor2_1 _13112_ (.Y(_02750_),
    .A(net2687),
    .B(net2789));
 sg13g2_nand3_1 _13113_ (.B(_02749_),
    .C(_02750_),
    .A(_00473_),
    .Y(_02751_));
 sg13g2_a21o_1 _13114_ (.A2(_02749_),
    .A1(_00473_),
    .B1(_02750_),
    .X(_02752_));
 sg13g2_nand2_1 _13115_ (.Y(_02753_),
    .A(_02751_),
    .B(_02752_));
 sg13g2_xnor2_1 _13116_ (.Y(_02754_),
    .A(_02748_),
    .B(_02753_));
 sg13g2_nor2_1 _13117_ (.A(_02744_),
    .B(_02754_),
    .Y(_02755_));
 sg13g2_nand2_1 _13118_ (.Y(_02756_),
    .A(_02744_),
    .B(_02754_));
 sg13g2_xnor2_1 _13119_ (.Y(_02757_),
    .A(_02744_),
    .B(_02754_));
 sg13g2_a22oi_1 _13120_ (.Y(_02758_),
    .B1(net2691),
    .B2(_05990_),
    .A2(_05649_),
    .A1(net2810));
 sg13g2_o21ai_1 _13121_ (.B1(_02758_),
    .Y(_02759_),
    .A1(net2691),
    .A2(_05990_));
 sg13g2_nor2_1 _13122_ (.A(\net.in[10] ),
    .B(net2782),
    .Y(_02760_));
 sg13g2_xnor2_1 _13123_ (.Y(_02761_),
    .A(net2635),
    .B(net2666));
 sg13g2_xor2_1 _13124_ (.B(net2735),
    .A(net2681),
    .X(_02762_));
 sg13g2_xnor2_1 _13125_ (.Y(_02763_),
    .A(_02761_),
    .B(_02762_));
 sg13g2_or3_1 _13126_ (.A(_02504_),
    .B(_02760_),
    .C(_02763_),
    .X(_02764_));
 sg13g2_o21ai_1 _13127_ (.B1(_02763_),
    .Y(_02765_),
    .A1(_02504_),
    .A2(_02760_));
 sg13g2_nand2_1 _13128_ (.Y(_02766_),
    .A(_02764_),
    .B(_02765_));
 sg13g2_xor2_1 _13129_ (.B(_02766_),
    .A(_02759_),
    .X(_02767_));
 sg13g2_xnor2_1 _13130_ (.Y(_02768_),
    .A(_02757_),
    .B(_02767_));
 sg13g2_nand2b_1 _13131_ (.Y(_02769_),
    .B(net2391),
    .A_N(net2494));
 sg13g2_nand2b_1 _13132_ (.Y(_02770_),
    .B(net2494),
    .A_N(net2391));
 sg13g2_nand2b_1 _13133_ (.Y(_02771_),
    .B(net2442),
    .A_N(net2669));
 sg13g2_nand3_1 _13134_ (.B(_02770_),
    .C(_02771_),
    .A(_02769_),
    .Y(_02772_));
 sg13g2_nor2_2 _13135_ (.A(net2679),
    .B(net2672),
    .Y(_02773_));
 sg13g2_nor2b_1 _13136_ (.A(net2564),
    .B_N(net2347),
    .Y(_02774_));
 sg13g2_xnor2_1 _13137_ (.Y(_02775_),
    .A(_02773_),
    .B(_02774_));
 sg13g2_inv_1 _13138_ (.Y(_02776_),
    .A(_02775_));
 sg13g2_nand2_1 _13139_ (.Y(_02777_),
    .A(_02772_),
    .B(_02776_));
 sg13g2_xor2_1 _13140_ (.B(_02775_),
    .A(_02772_),
    .X(_02778_));
 sg13g2_nand2_1 _13141_ (.Y(_02779_),
    .A(net2485),
    .B(net2394));
 sg13g2_nor2_1 _13142_ (.A(_05407_),
    .B(net2576),
    .Y(_02780_));
 sg13g2_xnor2_1 _13143_ (.Y(_02781_),
    .A(_02779_),
    .B(_02780_));
 sg13g2_xnor2_1 _13144_ (.Y(_02782_),
    .A(_02778_),
    .B(_02781_));
 sg13g2_xnor2_1 _13145_ (.Y(_02783_),
    .A(net2446),
    .B(net2440));
 sg13g2_xor2_1 _13146_ (.B(net2673),
    .A(net2629),
    .X(_02784_));
 sg13g2_nor2_1 _13147_ (.A(net2289),
    .B(net2779),
    .Y(_02785_));
 sg13g2_o21ai_1 _13148_ (.B1(_02785_),
    .Y(_02786_),
    .A1(_02783_),
    .A2(_02784_));
 sg13g2_nor3_1 _13149_ (.A(_02783_),
    .B(_02784_),
    .C(_02785_),
    .Y(_02787_));
 sg13g2_or3_1 _13150_ (.A(_02783_),
    .B(_02784_),
    .C(_02785_),
    .X(_02788_));
 sg13g2_nand2_1 _13151_ (.Y(_02789_),
    .A(_02786_),
    .B(_02788_));
 sg13g2_xnor2_1 _13152_ (.Y(_02790_),
    .A(_02749_),
    .B(_02789_));
 sg13g2_nor2_1 _13153_ (.A(_02782_),
    .B(_02790_),
    .Y(_02791_));
 sg13g2_xnor2_1 _13154_ (.Y(_02792_),
    .A(_02782_),
    .B(_02790_));
 sg13g2_nor2_1 _13155_ (.A(net2661),
    .B(net2618),
    .Y(_02793_));
 sg13g2_nand2b_1 _13156_ (.Y(_02794_),
    .B(net2253),
    .A_N(net2190));
 sg13g2_a21oi_1 _13157_ (.A1(_05363_),
    .A2(net2754),
    .Y(_02795_),
    .B1(_02794_));
 sg13g2_nor2b_1 _13158_ (.A(net2813),
    .B_N(net2728),
    .Y(_02796_));
 sg13g2_xnor2_1 _13159_ (.Y(_02797_),
    .A(net2789),
    .B(_02796_));
 sg13g2_nand2_1 _13160_ (.Y(_02798_),
    .A(_02795_),
    .B(_02797_));
 sg13g2_or2_1 _13161_ (.X(_02799_),
    .B(_02797_),
    .A(_02795_));
 sg13g2_nand2_1 _13162_ (.Y(_02800_),
    .A(_02798_),
    .B(_02799_));
 sg13g2_xor2_1 _13163_ (.B(_02800_),
    .A(_02793_),
    .X(_02801_));
 sg13g2_xnor2_1 _13164_ (.Y(_02802_),
    .A(_02792_),
    .B(_02801_));
 sg13g2_nand2_1 _13165_ (.Y(_02803_),
    .A(_02768_),
    .B(_02802_));
 sg13g2_or2_1 _13166_ (.X(_02804_),
    .B(_02803_),
    .A(_02735_));
 sg13g2_nor2_1 _13167_ (.A(_02768_),
    .B(_02802_),
    .Y(_02805_));
 sg13g2_and2_1 _13168_ (.A(_02735_),
    .B(_02805_),
    .X(_02806_));
 sg13g2_o21ai_1 _13169_ (.B1(_02803_),
    .Y(_02807_),
    .A1(_02735_),
    .A2(_02805_));
 sg13g2_a21o_1 _13170_ (.A2(_02807_),
    .A1(_02804_),
    .B1(_02806_),
    .X(_02808_));
 sg13g2_nand2_1 _13171_ (.Y(_02809_),
    .A(_02580_),
    .B(_02699_));
 sg13g2_o21ai_1 _13172_ (.B1(_02808_),
    .Y(_02810_),
    .A1(_02580_),
    .A2(_02699_));
 sg13g2_nand2_1 _13173_ (.Y(_02811_),
    .A(_02809_),
    .B(_02810_));
 sg13g2_nor2_1 _13174_ (.A(net2260),
    .B(net2799),
    .Y(_02812_));
 sg13g2_xnor2_1 _13175_ (.Y(_02813_),
    .A(_00024_),
    .B(_02812_));
 sg13g2_xnor2_1 _13176_ (.Y(_02814_),
    .A(net2670),
    .B(net2676));
 sg13g2_nor3_2 _13177_ (.A(\net.in[4] ),
    .B(\net.in[29] ),
    .C(_02814_),
    .Y(_02815_));
 sg13g2_nand2b_1 _13178_ (.Y(_02816_),
    .B(net2582),
    .A_N(net2625));
 sg13g2_nor2_1 _13179_ (.A(net2753),
    .B(net2758),
    .Y(_02817_));
 sg13g2_xnor2_1 _13180_ (.Y(_02818_),
    .A(_02816_),
    .B(_02817_));
 sg13g2_nor2b_1 _13181_ (.A(_02818_),
    .B_N(_02815_),
    .Y(_02819_));
 sg13g2_nand2b_1 _13182_ (.Y(_02820_),
    .B(_02818_),
    .A_N(_02815_));
 sg13g2_nand2b_1 _13183_ (.Y(_02821_),
    .B(_02820_),
    .A_N(_02819_));
 sg13g2_xnor2_1 _13184_ (.Y(_02822_),
    .A(_02813_),
    .B(_02821_));
 sg13g2_nand2b_1 _13185_ (.Y(_02823_),
    .B(net2692),
    .A_N(net2589));
 sg13g2_xnor2_1 _13186_ (.Y(_02824_),
    .A(net2588),
    .B(net2691));
 sg13g2_xor2_1 _13187_ (.B(net2741),
    .A(net2661),
    .X(_02825_));
 sg13g2_xnor2_1 _13188_ (.Y(_02826_),
    .A(_02548_),
    .B(_02825_));
 sg13g2_nand3_1 _13189_ (.B(_01113_),
    .C(_02826_),
    .A(_05407_),
    .Y(_02827_));
 sg13g2_a21o_1 _13190_ (.A2(_01113_),
    .A1(_05407_),
    .B1(_02826_),
    .X(_02828_));
 sg13g2_and2_1 _13191_ (.A(_02827_),
    .B(_02828_),
    .X(_02829_));
 sg13g2_xor2_1 _13192_ (.B(_02829_),
    .A(_02824_),
    .X(_02830_));
 sg13g2_xor2_1 _13193_ (.B(net2782),
    .A(net2721),
    .X(_02831_));
 sg13g2_xor2_1 _13194_ (.B(net2213),
    .A(net2192),
    .X(_02832_));
 sg13g2_nor2_1 _13195_ (.A(_02831_),
    .B(_02832_),
    .Y(_02833_));
 sg13g2_nor2_2 _13196_ (.A(\net.in[13] ),
    .B(net2774),
    .Y(_02834_));
 sg13g2_nand2_2 _13197_ (.Y(_02835_),
    .A(net2306),
    .B(net2341));
 sg13g2_xnor2_1 _13198_ (.Y(_02836_),
    .A(net2308),
    .B(net2343));
 sg13g2_and2_2 _13199_ (.A(_02834_),
    .B(_02836_),
    .X(_02837_));
 sg13g2_xnor2_1 _13200_ (.Y(_02838_),
    .A(net2781),
    .B(_00574_));
 sg13g2_nand2_1 _13201_ (.Y(_02839_),
    .A(_02837_),
    .B(_02838_));
 sg13g2_nor2_1 _13202_ (.A(_02837_),
    .B(_02838_),
    .Y(_02840_));
 sg13g2_xnor2_1 _13203_ (.Y(_02841_),
    .A(_02837_),
    .B(_02838_));
 sg13g2_xnor2_1 _13204_ (.Y(_02842_),
    .A(_02833_),
    .B(_02841_));
 sg13g2_nand2_1 _13205_ (.Y(_02843_),
    .A(_02830_),
    .B(_02842_));
 sg13g2_nor2_1 _13206_ (.A(_02830_),
    .B(_02842_),
    .Y(_02844_));
 sg13g2_o21ai_1 _13207_ (.B1(_02843_),
    .Y(_02845_),
    .A1(_02822_),
    .A2(_02844_));
 sg13g2_xnor2_1 _13208_ (.Y(_02846_),
    .A(_02830_),
    .B(_02842_));
 sg13g2_xnor2_1 _13209_ (.Y(_02847_),
    .A(_02822_),
    .B(_02846_));
 sg13g2_nor4_2 _13210_ (.A(net2180),
    .B(net2189),
    .C(net2731),
    .Y(_02848_),
    .D(net2647));
 sg13g2_nor2_1 _13211_ (.A(net2617),
    .B(net2626),
    .Y(_02849_));
 sg13g2_xor2_1 _13212_ (.B(net2625),
    .A(net2615),
    .X(_02850_));
 sg13g2_nor2_1 _13213_ (.A(_02746_),
    .B(_02850_),
    .Y(_02851_));
 sg13g2_o21ai_1 _13214_ (.B1(_00016_),
    .Y(_02852_),
    .A1(net2300),
    .A2(net2812));
 sg13g2_a21oi_2 _13215_ (.B1(_02852_),
    .Y(_02853_),
    .A2(net2813),
    .A1(net2300));
 sg13g2_nor2_1 _13216_ (.A(_02851_),
    .B(_02853_),
    .Y(_02854_));
 sg13g2_xnor2_1 _13217_ (.Y(_02855_),
    .A(_02851_),
    .B(_02853_));
 sg13g2_xnor2_1 _13218_ (.Y(_02856_),
    .A(_02848_),
    .B(_02855_));
 sg13g2_nor2b_1 _13219_ (.A(net2730),
    .B_N(net2287),
    .Y(_02857_));
 sg13g2_xnor2_1 _13220_ (.Y(_02858_),
    .A(_00011_),
    .B(_02857_));
 sg13g2_xnor2_1 _13221_ (.Y(_02859_),
    .A(net2216),
    .B(net2711));
 sg13g2_xnor2_1 _13222_ (.Y(_02860_),
    .A(net2716),
    .B(net2635));
 sg13g2_nand2_1 _13223_ (.Y(_02861_),
    .A(_02859_),
    .B(_02860_));
 sg13g2_nand2b_1 _13224_ (.Y(_02862_),
    .B(_02858_),
    .A_N(_02861_));
 sg13g2_nor2b_1 _13225_ (.A(_02858_),
    .B_N(_02861_),
    .Y(_02863_));
 sg13g2_xor2_1 _13226_ (.B(_02861_),
    .A(_02858_),
    .X(_02864_));
 sg13g2_nand2_1 _13227_ (.Y(_02865_),
    .A(_05495_),
    .B(net2635));
 sg13g2_xnor2_1 _13228_ (.Y(_02866_),
    .A(net2661),
    .B(net2674));
 sg13g2_xnor2_1 _13229_ (.Y(_02867_),
    .A(_02865_),
    .B(_02866_));
 sg13g2_xnor2_1 _13230_ (.Y(_02868_),
    .A(_02864_),
    .B(_02867_));
 sg13g2_nor2_1 _13231_ (.A(_02856_),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_nand2_1 _13232_ (.Y(_02870_),
    .A(_02856_),
    .B(_02868_));
 sg13g2_xor2_1 _13233_ (.B(_02868_),
    .A(_02856_),
    .X(_02871_));
 sg13g2_xor2_1 _13234_ (.B(net2639),
    .A(net2721),
    .X(_02872_));
 sg13g2_xnor2_1 _13235_ (.Y(_02873_),
    .A(net2766),
    .B(net2547));
 sg13g2_nor3_2 _13236_ (.A(net2816),
    .B(net2814),
    .C(_02873_),
    .Y(_02874_));
 sg13g2_a22oi_1 _13237_ (.Y(_02875_),
    .B1(_06078_),
    .B2(net2231),
    .A2(_05847_),
    .A1(_05055_));
 sg13g2_o21ai_1 _13238_ (.B1(_02875_),
    .Y(_02876_),
    .A1(net2231),
    .A2(_06078_));
 sg13g2_nand2_1 _13239_ (.Y(_02877_),
    .A(_02874_),
    .B(_02876_));
 sg13g2_xnor2_1 _13240_ (.Y(_02878_),
    .A(_02874_),
    .B(_02876_));
 sg13g2_xnor2_1 _13241_ (.Y(_02879_),
    .A(_02872_),
    .B(_02878_));
 sg13g2_xnor2_1 _13242_ (.Y(_02880_),
    .A(_02871_),
    .B(_02879_));
 sg13g2_nor2_1 _13243_ (.A(net2452),
    .B(_05165_),
    .Y(_02881_));
 sg13g2_nand2b_1 _13244_ (.Y(_02882_),
    .B(net2777),
    .A_N(net2547));
 sg13g2_xor2_1 _13245_ (.B(net2216),
    .A(net2719),
    .X(_02883_));
 sg13g2_xnor2_1 _13246_ (.Y(_02884_),
    .A(_02882_),
    .B(_02883_));
 sg13g2_nand2_1 _13247_ (.Y(_02885_),
    .A(_02881_),
    .B(_02884_));
 sg13g2_xor2_1 _13248_ (.B(_02884_),
    .A(_02881_),
    .X(_02886_));
 sg13g2_nor2_1 _13249_ (.A(_05594_),
    .B(net2565),
    .Y(_02887_));
 sg13g2_xor2_1 _13250_ (.B(net2666),
    .A(net2674),
    .X(_02888_));
 sg13g2_xnor2_1 _13251_ (.Y(_02889_),
    .A(_02887_),
    .B(_02888_));
 sg13g2_nand2_1 _13252_ (.Y(_02890_),
    .A(_02885_),
    .B(_02889_));
 sg13g2_o21ai_1 _13253_ (.B1(_02890_),
    .Y(_02891_),
    .A1(_02881_),
    .A2(_02884_));
 sg13g2_xnor2_1 _13254_ (.Y(_02892_),
    .A(_02886_),
    .B(_02889_));
 sg13g2_nor2b_2 _13255_ (.A(net2576),
    .B_N(net2405),
    .Y(_02893_));
 sg13g2_o21ai_1 _13256_ (.B1(net2290),
    .Y(_02894_),
    .A1(net2699),
    .A2(net2425));
 sg13g2_nor3_1 _13257_ (.A(net2645),
    .B(_01203_),
    .C(_02894_),
    .Y(_02895_));
 sg13g2_o21ai_1 _13258_ (.B1(_01203_),
    .Y(_02896_),
    .A1(net2642),
    .A2(_02894_));
 sg13g2_nor2b_1 _13259_ (.A(_02895_),
    .B_N(_02896_),
    .Y(_02897_));
 sg13g2_xnor2_1 _13260_ (.Y(_02898_),
    .A(_02893_),
    .B(_02897_));
 sg13g2_nor2_1 _13261_ (.A(_02892_),
    .B(_02898_),
    .Y(_02899_));
 sg13g2_xor2_1 _13262_ (.B(_02898_),
    .A(_02892_),
    .X(_02900_));
 sg13g2_xnor2_1 _13263_ (.Y(_02901_),
    .A(net2204),
    .B(net2605));
 sg13g2_xnor2_1 _13264_ (.Y(_02902_),
    .A(net2661),
    .B(net2602));
 sg13g2_nand3_1 _13265_ (.B(_02901_),
    .C(_02902_),
    .A(_08366_),
    .Y(_02903_));
 sg13g2_a21o_1 _13266_ (.A2(_02902_),
    .A1(_02901_),
    .B1(_08366_),
    .X(_02904_));
 sg13g2_nand2_1 _13267_ (.Y(_02905_),
    .A(_02903_),
    .B(_02904_));
 sg13g2_nor2_1 _13268_ (.A(net2805),
    .B(_05792_),
    .Y(_02906_));
 sg13g2_nor2_1 _13269_ (.A(net2807),
    .B(net2187),
    .Y(_02907_));
 sg13g2_xnor2_1 _13270_ (.Y(_02908_),
    .A(_02906_),
    .B(_02907_));
 sg13g2_nand2_1 _13271_ (.Y(_02909_),
    .A(_02903_),
    .B(_02908_));
 sg13g2_xnor2_1 _13272_ (.Y(_02910_),
    .A(_02905_),
    .B(_02908_));
 sg13g2_xnor2_1 _13273_ (.Y(_02911_),
    .A(_02900_),
    .B(_02910_));
 sg13g2_nand2_1 _13274_ (.Y(_02912_),
    .A(_02880_),
    .B(_02911_));
 sg13g2_or2_1 _13275_ (.X(_02913_),
    .B(_02911_),
    .A(_02880_));
 sg13g2_inv_1 _13276_ (.Y(_02914_),
    .A(_02913_));
 sg13g2_nand2_1 _13277_ (.Y(_02915_),
    .A(_02912_),
    .B(_02913_));
 sg13g2_o21ai_1 _13278_ (.B1(_02912_),
    .Y(_02916_),
    .A1(_02847_),
    .A2(_02914_));
 sg13g2_xor2_1 _13279_ (.B(_02915_),
    .A(_02847_),
    .X(_02917_));
 sg13g2_xnor2_1 _13280_ (.Y(_02918_),
    .A(net2204),
    .B(net2197));
 sg13g2_xnor2_1 _13281_ (.Y(_02919_),
    .A(net2526),
    .B(net2635));
 sg13g2_nand2_2 _13282_ (.Y(_02920_),
    .A(_02918_),
    .B(_02919_));
 sg13g2_xnor2_1 _13283_ (.Y(_02921_),
    .A(net2498),
    .B(net2803));
 sg13g2_o21ai_1 _13284_ (.B1(_02921_),
    .Y(_02922_),
    .A1(net2678),
    .A2(_05682_));
 sg13g2_xnor2_1 _13285_ (.Y(_02923_),
    .A(net2422),
    .B(net2435));
 sg13g2_inv_1 _13286_ (.Y(_02924_),
    .A(_02923_));
 sg13g2_nor2_1 _13287_ (.A(net2187),
    .B(net2669),
    .Y(_02925_));
 sg13g2_xnor2_1 _13288_ (.Y(_02926_),
    .A(net2661),
    .B(net2221));
 sg13g2_xnor2_1 _13289_ (.Y(_02927_),
    .A(_02925_),
    .B(_02926_));
 sg13g2_nand2_1 _13290_ (.Y(_02928_),
    .A(_02924_),
    .B(_02927_));
 sg13g2_o21ai_1 _13291_ (.B1(_02922_),
    .Y(_02929_),
    .A1(_02924_),
    .A2(_02927_));
 sg13g2_nand2_2 _13292_ (.Y(_02930_),
    .A(_02928_),
    .B(_02929_));
 sg13g2_xnor2_1 _13293_ (.Y(_02931_),
    .A(_02924_),
    .B(_02927_));
 sg13g2_xnor2_1 _13294_ (.Y(_02932_),
    .A(_02922_),
    .B(_02931_));
 sg13g2_xnor2_1 _13295_ (.Y(_02933_),
    .A(net2674),
    .B(net2273));
 sg13g2_xnor2_1 _13296_ (.Y(_02934_),
    .A(net2686),
    .B(net2756));
 sg13g2_nand3_1 _13297_ (.B(_02933_),
    .C(_02934_),
    .A(net2296),
    .Y(_02935_));
 sg13g2_a21oi_1 _13298_ (.A1(net2296),
    .A2(_02933_),
    .Y(_02936_),
    .B1(_02934_));
 sg13g2_a21o_1 _13299_ (.A2(_02933_),
    .A1(net2296),
    .B1(_02934_),
    .X(_02937_));
 sg13g2_and2_1 _13300_ (.A(_02935_),
    .B(_02937_),
    .X(_02938_));
 sg13g2_xnor2_1 _13301_ (.Y(_02939_),
    .A(_02703_),
    .B(_02938_));
 sg13g2_xnor2_1 _13302_ (.Y(_02940_),
    .A(_02932_),
    .B(_02939_));
 sg13g2_nor2_2 _13303_ (.A(net2430),
    .B(net2499),
    .Y(_02941_));
 sg13g2_a22oi_1 _13304_ (.Y(_02942_),
    .B1(_06023_),
    .B2(net2378),
    .A2(_05561_),
    .A1(net2429));
 sg13g2_nor2_1 _13305_ (.A(net2400),
    .B(net2676),
    .Y(_02943_));
 sg13g2_nand2_1 _13306_ (.Y(_02944_),
    .A(net2436),
    .B(_05528_));
 sg13g2_xnor2_1 _13307_ (.Y(_02945_),
    .A(_02943_),
    .B(_02944_));
 sg13g2_nand2_1 _13308_ (.Y(_02946_),
    .A(_02942_),
    .B(_02945_));
 sg13g2_xor2_1 _13309_ (.B(_02945_),
    .A(_02942_),
    .X(_02947_));
 sg13g2_xnor2_1 _13310_ (.Y(_02948_),
    .A(_02941_),
    .B(_02947_));
 sg13g2_xnor2_1 _13311_ (.Y(_02949_),
    .A(_02940_),
    .B(_02948_));
 sg13g2_a21oi_2 _13312_ (.B1(_07552_),
    .Y(_02950_),
    .A2(net2778),
    .A1(_05814_));
 sg13g2_inv_1 _13313_ (.Y(_02951_),
    .A(_02950_));
 sg13g2_xor2_1 _13314_ (.B(net2197),
    .A(net2660),
    .X(_02952_));
 sg13g2_xor2_1 _13315_ (.B(net2572),
    .A(net2630),
    .X(_02953_));
 sg13g2_nor2_2 _13316_ (.A(_02952_),
    .B(_02953_),
    .Y(_02954_));
 sg13g2_nand2_1 _13317_ (.Y(_02955_),
    .A(net2804),
    .B(_02954_));
 sg13g2_xor2_1 _13318_ (.B(_02954_),
    .A(net2804),
    .X(_02956_));
 sg13g2_xnor2_1 _13319_ (.Y(_02957_),
    .A(_02951_),
    .B(_02956_));
 sg13g2_nand2b_1 _13320_ (.Y(_02958_),
    .B(net2781),
    .A_N(net2510));
 sg13g2_o21ai_1 _13321_ (.B1(_02958_),
    .Y(_02959_),
    .A1(net2721),
    .A2(net2754));
 sg13g2_a21oi_2 _13322_ (.B1(net2661),
    .Y(_02960_),
    .A2(_06045_),
    .A1(net2764));
 sg13g2_nand2_1 _13323_ (.Y(_02961_),
    .A(_02959_),
    .B(_02960_));
 sg13g2_xor2_1 _13324_ (.B(_02960_),
    .A(_02959_),
    .X(_02962_));
 sg13g2_nor2_1 _13325_ (.A(net2224),
    .B(\net.in[13] ),
    .Y(_02963_));
 sg13g2_nor2b_1 _13326_ (.A(net2721),
    .B_N(net2289),
    .Y(_02964_));
 sg13g2_xnor2_1 _13327_ (.Y(_02965_),
    .A(_02963_),
    .B(_02964_));
 sg13g2_xnor2_1 _13328_ (.Y(_02966_),
    .A(_02962_),
    .B(_02965_));
 sg13g2_nand2_1 _13329_ (.Y(_02967_),
    .A(_02957_),
    .B(_02966_));
 sg13g2_xor2_1 _13330_ (.B(_02966_),
    .A(_02957_),
    .X(_02968_));
 sg13g2_xnor2_1 _13331_ (.Y(_02969_),
    .A(net2348),
    .B(net2355));
 sg13g2_xor2_1 _13332_ (.B(net2276),
    .A(net2238),
    .X(_02970_));
 sg13g2_nor2_1 _13333_ (.A(_02969_),
    .B(_02970_),
    .Y(_02971_));
 sg13g2_xnor2_1 _13334_ (.Y(_02972_),
    .A(net2752),
    .B(net2557));
 sg13g2_nor3_1 _13335_ (.A(_02969_),
    .B(_02970_),
    .C(_02972_),
    .Y(_02973_));
 sg13g2_nor2b_1 _13336_ (.A(_02971_),
    .B_N(_02972_),
    .Y(_02974_));
 sg13g2_inv_1 _13337_ (.Y(_02975_),
    .A(_02974_));
 sg13g2_nor2_1 _13338_ (.A(_02973_),
    .B(_02974_),
    .Y(_02976_));
 sg13g2_xnor2_1 _13339_ (.Y(_02977_),
    .A(net2630),
    .B(_02703_));
 sg13g2_xnor2_1 _13340_ (.Y(_02978_),
    .A(_02976_),
    .B(_02977_));
 sg13g2_o21ai_1 _13341_ (.B1(_02978_),
    .Y(_02979_),
    .A1(_02957_),
    .A2(_02966_));
 sg13g2_xnor2_1 _13342_ (.Y(_02980_),
    .A(_02968_),
    .B(_02978_));
 sg13g2_nor2_1 _13343_ (.A(_02949_),
    .B(_02980_),
    .Y(_02981_));
 sg13g2_and2_1 _13344_ (.A(_02949_),
    .B(_02980_),
    .X(_02982_));
 sg13g2_nor2_1 _13345_ (.A(_02981_),
    .B(_02982_),
    .Y(_02983_));
 sg13g2_xnor2_1 _13346_ (.Y(_02984_),
    .A(_02920_),
    .B(_02983_));
 sg13g2_nand2_1 _13347_ (.Y(_02985_),
    .A(_02917_),
    .B(_02984_));
 sg13g2_xor2_1 _13348_ (.B(_02699_),
    .A(_02580_),
    .X(_02986_));
 sg13g2_xnor2_1 _13349_ (.Y(_02987_),
    .A(_02808_),
    .B(_02986_));
 sg13g2_nor2_1 _13350_ (.A(_02917_),
    .B(_02984_),
    .Y(_02988_));
 sg13g2_inv_1 _13351_ (.Y(_02989_),
    .A(_02988_));
 sg13g2_a21oi_1 _13352_ (.A1(_02985_),
    .A2(_02987_),
    .Y(_02990_),
    .B1(_02988_));
 sg13g2_and2_1 _13353_ (.A(_02811_),
    .B(_02990_),
    .X(_02991_));
 sg13g2_xor2_1 _13354_ (.B(_02990_),
    .A(_02811_),
    .X(_02992_));
 sg13g2_nand2_1 _13355_ (.Y(_02993_),
    .A(_02542_),
    .B(_02579_));
 sg13g2_o21ai_1 _13356_ (.B1(_02698_),
    .Y(_02994_),
    .A1(_02621_),
    .A2(_02661_));
 sg13g2_a22oi_1 _13357_ (.Y(_02995_),
    .B1(_02994_),
    .B2(_02662_),
    .A2(_02993_),
    .A1(_02541_));
 sg13g2_and4_1 _13358_ (.A(_02541_),
    .B(_02662_),
    .C(_02993_),
    .D(_02994_),
    .X(_02996_));
 sg13g2_nor2_1 _13359_ (.A(_02995_),
    .B(_02996_),
    .Y(_02997_));
 sg13g2_nor2_1 _13360_ (.A(_02807_),
    .B(_02995_),
    .Y(_02998_));
 sg13g2_nor2_1 _13361_ (.A(_02996_),
    .B(_02998_),
    .Y(_02999_));
 sg13g2_xnor2_1 _13362_ (.Y(_03000_),
    .A(_02807_),
    .B(_02997_));
 sg13g2_nor2_1 _13363_ (.A(_02920_),
    .B(_02981_),
    .Y(_03001_));
 sg13g2_o21ai_1 _13364_ (.B1(_02916_),
    .Y(_03002_),
    .A1(_02982_),
    .A2(_03001_));
 sg13g2_inv_1 _13365_ (.Y(_03003_),
    .A(_03002_));
 sg13g2_nor3_1 _13366_ (.A(_02916_),
    .B(_02982_),
    .C(_03001_),
    .Y(_03004_));
 sg13g2_nor2_1 _13367_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sg13g2_o21ai_1 _13368_ (.B1(_02607_),
    .Y(_03006_),
    .A1(_02606_),
    .A2(_02620_));
 sg13g2_or2_1 _13369_ (.X(_03007_),
    .B(_03006_),
    .A(_03004_));
 sg13g2_xnor2_1 _13370_ (.Y(_03008_),
    .A(_03005_),
    .B(_03006_));
 sg13g2_a21o_1 _13371_ (.A2(_03000_),
    .A1(_02992_),
    .B1(_03008_),
    .X(_03009_));
 sg13g2_o21ai_1 _13372_ (.B1(_03009_),
    .Y(_03010_),
    .A1(_02992_),
    .A2(_03000_));
 sg13g2_nand2_1 _13373_ (.Y(_03011_),
    .A(_02478_),
    .B(_02482_));
 sg13g2_and2_1 _13374_ (.A(_02483_),
    .B(_03011_),
    .X(_03012_));
 sg13g2_nor2_1 _13375_ (.A(_02688_),
    .B(_02695_),
    .Y(_03013_));
 sg13g2_nor2_1 _13376_ (.A(_02694_),
    .B(_03013_),
    .Y(_03014_));
 sg13g2_nor2_1 _13377_ (.A(_02486_),
    .B(_02491_),
    .Y(_03015_));
 sg13g2_nor2_1 _13378_ (.A(_02492_),
    .B(_03015_),
    .Y(_03016_));
 sg13g2_nor3_1 _13379_ (.A(_02694_),
    .B(_03013_),
    .C(_03016_),
    .Y(_03017_));
 sg13g2_inv_1 _13380_ (.Y(_03018_),
    .A(_03017_));
 sg13g2_nor2b_1 _13381_ (.A(_03014_),
    .B_N(_03016_),
    .Y(_03019_));
 sg13g2_a21oi_2 _13382_ (.B1(_03019_),
    .Y(_03020_),
    .A2(_03018_),
    .A1(_03012_));
 sg13g2_a21o_1 _13383_ (.A2(_03019_),
    .A1(_03012_),
    .B1(_03020_),
    .X(_03021_));
 sg13g2_o21ai_1 _13384_ (.B1(_03021_),
    .Y(_03022_),
    .A1(_03012_),
    .A2(_03018_));
 sg13g2_o21ai_1 _13385_ (.B1(_02657_),
    .Y(_03023_),
    .A1(_02650_),
    .A2(_02658_));
 sg13g2_inv_1 _13386_ (.Y(_03024_),
    .A(_03023_));
 sg13g2_a21oi_2 _13387_ (.B1(_02681_),
    .Y(_03025_),
    .A2(_02682_),
    .A1(_02674_));
 sg13g2_nand2_1 _13388_ (.Y(_03026_),
    .A(_03024_),
    .B(_03025_));
 sg13g2_nor2_1 _13389_ (.A(_03024_),
    .B(_03025_),
    .Y(_03027_));
 sg13g2_xnor2_1 _13390_ (.Y(_03028_),
    .A(_03023_),
    .B(_03025_));
 sg13g2_nand2_1 _13391_ (.Y(_03029_),
    .A(_02666_),
    .B(_02670_));
 sg13g2_o21ai_1 _13392_ (.B1(_03029_),
    .Y(_03030_),
    .A1(_02667_),
    .A2(_02669_));
 sg13g2_xnor2_1 _13393_ (.Y(_03031_),
    .A(_03028_),
    .B(_03030_));
 sg13g2_nand2_1 _13394_ (.Y(_03032_),
    .A(_03022_),
    .B(_03031_));
 sg13g2_or2_1 _13395_ (.X(_03033_),
    .B(_03031_),
    .A(_03022_));
 sg13g2_nand2_1 _13396_ (.Y(_03034_),
    .A(_03032_),
    .B(_03033_));
 sg13g2_or2_1 _13397_ (.X(_03035_),
    .B(_02510_),
    .A(_02503_));
 sg13g2_nand2_1 _13398_ (.Y(_03036_),
    .A(_02467_),
    .B(_02474_));
 sg13g2_a22oi_1 _13399_ (.Y(_03037_),
    .B1(_03036_),
    .B2(_02473_),
    .A2(_03035_),
    .A1(_02509_));
 sg13g2_nand4_1 _13400_ (.B(_02509_),
    .C(_03035_),
    .A(_02473_),
    .Y(_03038_),
    .D(_03036_));
 sg13g2_or2_1 _13401_ (.X(_03039_),
    .B(_03038_),
    .A(_02525_));
 sg13g2_a21oi_2 _13402_ (.B1(_03037_),
    .Y(_03040_),
    .A2(_03038_),
    .A1(_02525_));
 sg13g2_a22oi_1 _13403_ (.Y(_03041_),
    .B1(_03039_),
    .B2(_03040_),
    .A2(_03037_),
    .A1(_02525_));
 sg13g2_xor2_1 _13404_ (.B(_03041_),
    .A(_03034_),
    .X(_03042_));
 sg13g2_a21oi_2 _13405_ (.B1(_02561_),
    .Y(_03043_),
    .A2(_02562_),
    .A1(_02557_));
 sg13g2_a21oi_2 _13406_ (.B1(_02533_),
    .Y(_03044_),
    .A2(_02538_),
    .A1(_02534_));
 sg13g2_nand2_1 _13407_ (.Y(_03045_),
    .A(_03043_),
    .B(_03044_));
 sg13g2_nor2_1 _13408_ (.A(_03043_),
    .B(_03044_),
    .Y(_03046_));
 sg13g2_xor2_1 _13409_ (.B(_03044_),
    .A(_03043_),
    .X(_03047_));
 sg13g2_o21ai_1 _13410_ (.B1(_02553_),
    .Y(_03048_),
    .A1(_02547_),
    .A2(_02554_));
 sg13g2_xnor2_1 _13411_ (.Y(_03049_),
    .A(_03047_),
    .B(_03048_));
 sg13g2_o21ai_1 _13412_ (.B1(_02567_),
    .Y(_03050_),
    .A1(_02571_),
    .A2(_02575_));
 sg13g2_nand2_1 _13413_ (.Y(_03051_),
    .A(_02748_),
    .B(_02752_));
 sg13g2_a22oi_1 _13414_ (.Y(_03052_),
    .B1(_03051_),
    .B2(_02751_),
    .A2(_03050_),
    .A1(_02576_));
 sg13g2_nand4_1 _13415_ (.B(_02751_),
    .C(_03050_),
    .A(_02576_),
    .Y(_03053_),
    .D(_03051_));
 sg13g2_nor2b_1 _13416_ (.A(_03052_),
    .B_N(_03053_),
    .Y(_03054_));
 sg13g2_o21ai_1 _13417_ (.B1(_02741_),
    .Y(_03055_),
    .A1(_02737_),
    .A2(_02742_));
 sg13g2_xnor2_1 _13418_ (.Y(_03056_),
    .A(_03054_),
    .B(_03055_));
 sg13g2_nand2_1 _13419_ (.Y(_03057_),
    .A(_03049_),
    .B(_03056_));
 sg13g2_nor2_1 _13420_ (.A(_03049_),
    .B(_03056_),
    .Y(_03058_));
 sg13g2_xnor2_1 _13421_ (.Y(_03059_),
    .A(_03049_),
    .B(_03056_));
 sg13g2_a21o_1 _13422_ (.A2(_02786_),
    .A1(_02749_),
    .B1(_02787_),
    .X(_03060_));
 sg13g2_o21ai_1 _13423_ (.B1(_02781_),
    .Y(_03061_),
    .A1(_02772_),
    .A2(_02776_));
 sg13g2_nand2_1 _13424_ (.Y(_03062_),
    .A(_02759_),
    .B(_02765_));
 sg13g2_nand4_1 _13425_ (.B(_02777_),
    .C(_03061_),
    .A(_02764_),
    .Y(_03063_),
    .D(_03062_));
 sg13g2_a22oi_1 _13426_ (.Y(_03064_),
    .B1(_03062_),
    .B2(_02764_),
    .A2(_03061_),
    .A1(_02777_));
 sg13g2_nor2_1 _13427_ (.A(_03060_),
    .B(_03063_),
    .Y(_03065_));
 sg13g2_a21oi_2 _13428_ (.B1(_03064_),
    .Y(_03066_),
    .A2(_03063_),
    .A1(_03060_));
 sg13g2_a21oi_1 _13429_ (.A1(_03060_),
    .A2(_03064_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_nor2_2 _13430_ (.A(_03065_),
    .B(_03067_),
    .Y(_03068_));
 sg13g2_xnor2_1 _13431_ (.Y(_03069_),
    .A(_03059_),
    .B(_03068_));
 sg13g2_nand2_1 _13432_ (.Y(_03070_),
    .A(_03042_),
    .B(_03069_));
 sg13g2_or2_1 _13433_ (.X(_03071_),
    .B(_03069_),
    .A(_03042_));
 sg13g2_o21ai_1 _13434_ (.B1(_02724_),
    .Y(_03072_),
    .A1(_02725_),
    .A2(_02729_));
 sg13g2_nand2_1 _13435_ (.Y(_03073_),
    .A(_02793_),
    .B(_02799_));
 sg13g2_nand2_1 _13436_ (.Y(_03074_),
    .A(_02798_),
    .B(_03073_));
 sg13g2_a21oi_1 _13437_ (.A1(_02712_),
    .A2(_02715_),
    .Y(_03075_),
    .B1(_02710_));
 sg13g2_nor2_2 _13438_ (.A(_02716_),
    .B(_03075_),
    .Y(_03076_));
 sg13g2_xnor2_1 _13439_ (.Y(_03077_),
    .A(_03074_),
    .B(_03076_));
 sg13g2_a21o_1 _13440_ (.A2(_03076_),
    .A1(_03074_),
    .B1(_03072_),
    .X(_03078_));
 sg13g2_o21ai_1 _13441_ (.B1(_03078_),
    .Y(_03079_),
    .A1(_03074_),
    .A2(_03076_));
 sg13g2_xnor2_1 _13442_ (.Y(_03080_),
    .A(_03072_),
    .B(_03077_));
 sg13g2_nand2b_1 _13443_ (.Y(_03081_),
    .B(_02867_),
    .A_N(_02863_));
 sg13g2_a21oi_1 _13444_ (.A1(_02701_),
    .A2(_02707_),
    .Y(_03082_),
    .B1(_02706_));
 sg13g2_nand3_1 _13445_ (.B(_03081_),
    .C(_03082_),
    .A(_02862_),
    .Y(_03083_));
 sg13g2_a21o_1 _13446_ (.A2(_03081_),
    .A1(_02862_),
    .B1(_03082_),
    .X(_03084_));
 sg13g2_nand2_1 _13447_ (.Y(_03085_),
    .A(_03083_),
    .B(_03084_));
 sg13g2_a21oi_1 _13448_ (.A1(_02851_),
    .A2(_02853_),
    .Y(_03086_),
    .B1(_02848_));
 sg13g2_nor2_1 _13449_ (.A(_02854_),
    .B(_03086_),
    .Y(_03087_));
 sg13g2_nand2_1 _13450_ (.Y(_03088_),
    .A(_03083_),
    .B(_03087_));
 sg13g2_xnor2_1 _13451_ (.Y(_03089_),
    .A(_03085_),
    .B(_03087_));
 sg13g2_o21ai_1 _13452_ (.B1(_02872_),
    .Y(_03090_),
    .A1(_02874_),
    .A2(_02876_));
 sg13g2_nand2_2 _13453_ (.Y(_03091_),
    .A(_02877_),
    .B(_03090_));
 sg13g2_a21oi_2 _13454_ (.B1(_02895_),
    .Y(_03092_),
    .A2(_02896_),
    .A1(_02893_));
 sg13g2_nand2_1 _13455_ (.Y(_03093_),
    .A(_03091_),
    .B(_03092_));
 sg13g2_nor2_1 _13456_ (.A(_03091_),
    .B(_03092_),
    .Y(_03094_));
 sg13g2_xnor2_1 _13457_ (.Y(_03095_),
    .A(_03091_),
    .B(_03092_));
 sg13g2_xnor2_1 _13458_ (.Y(_03096_),
    .A(_02891_),
    .B(_03095_));
 sg13g2_a21o_1 _13459_ (.A2(_03089_),
    .A1(_03080_),
    .B1(_03096_),
    .X(_03097_));
 sg13g2_xnor2_1 _13460_ (.Y(_03098_),
    .A(_03080_),
    .B(_03089_));
 sg13g2_xnor2_1 _13461_ (.Y(_03099_),
    .A(_03096_),
    .B(_03098_));
 sg13g2_nand2_1 _13462_ (.Y(_03100_),
    .A(_03071_),
    .B(_03099_));
 sg13g2_a21oi_1 _13463_ (.A1(_03070_),
    .A2(_03100_),
    .Y(_03101_),
    .B1(_03010_));
 sg13g2_nand3_1 _13464_ (.B(_03070_),
    .C(_03100_),
    .A(_03010_),
    .Y(_03102_));
 sg13g2_nor2b_1 _13465_ (.A(_03101_),
    .B_N(_03102_),
    .Y(_03103_));
 sg13g2_a21o_1 _13466_ (.A2(_02564_),
    .A1(_02556_),
    .B1(_02578_),
    .X(_03104_));
 sg13g2_a21o_1 _13467_ (.A2(_02526_),
    .A1(_02512_),
    .B1(_02539_),
    .X(_03105_));
 sg13g2_a22oi_1 _13468_ (.Y(_03106_),
    .B1(_03105_),
    .B2(_02527_),
    .A2(_03104_),
    .A1(_02565_));
 sg13g2_and4_1 _13469_ (.A(_02527_),
    .B(_02565_),
    .C(_03104_),
    .D(_03105_),
    .X(_03107_));
 sg13g2_nor2_1 _13470_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sg13g2_o21ai_1 _13471_ (.B1(_02756_),
    .Y(_03109_),
    .A1(_02755_),
    .A2(_02767_));
 sg13g2_nor2_1 _13472_ (.A(_03106_),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_xor2_1 _13473_ (.B(_03109_),
    .A(_03108_),
    .X(_03111_));
 sg13g2_a21o_1 _13474_ (.A2(_02645_),
    .A1(_02632_),
    .B1(_02660_),
    .X(_03112_));
 sg13g2_o21ai_1 _13475_ (.B1(_03112_),
    .Y(_03113_),
    .A1(_02632_),
    .A2(_02645_));
 sg13g2_nand2_1 _13476_ (.Y(_03114_),
    .A(_02686_),
    .B(_02697_));
 sg13g2_a21oi_1 _13477_ (.A1(_02685_),
    .A2(_03114_),
    .Y(_03115_),
    .B1(_03113_));
 sg13g2_and3_1 _13478_ (.X(_03116_),
    .A(_02685_),
    .B(_03113_),
    .C(_03114_));
 sg13g2_nor2_1 _13479_ (.A(_03115_),
    .B(_03116_),
    .Y(_03117_));
 sg13g2_xnor2_1 _13480_ (.Y(_03118_),
    .A(_02500_),
    .B(_03117_));
 sg13g2_nor2b_1 _13481_ (.A(_03111_),
    .B_N(_03118_),
    .Y(_03119_));
 sg13g2_nand2b_1 _13482_ (.Y(_03120_),
    .B(_03111_),
    .A_N(_03118_));
 sg13g2_nor2_1 _13483_ (.A(_02791_),
    .B(_02801_),
    .Y(_03121_));
 sg13g2_a21oi_2 _13484_ (.B1(_03121_),
    .Y(_03122_),
    .A2(_02790_),
    .A1(_02782_));
 sg13g2_nand2_1 _13485_ (.Y(_03123_),
    .A(_02734_),
    .B(_03122_));
 sg13g2_nor2_1 _13486_ (.A(_02734_),
    .B(_03122_),
    .Y(_03124_));
 sg13g2_xor2_1 _13487_ (.B(_03122_),
    .A(_02734_),
    .X(_03125_));
 sg13g2_o21ai_1 _13488_ (.B1(_02870_),
    .Y(_03126_),
    .A1(_02869_),
    .A2(_02879_));
 sg13g2_xnor2_1 _13489_ (.Y(_03127_),
    .A(_03125_),
    .B(_03126_));
 sg13g2_o21ai_1 _13490_ (.B1(_03120_),
    .Y(_03128_),
    .A1(_03119_),
    .A2(_03127_));
 sg13g2_xnor2_1 _13491_ (.Y(_03129_),
    .A(_03103_),
    .B(_03128_));
 sg13g2_inv_1 _13492_ (.Y(_03130_),
    .A(_03129_));
 sg13g2_nor2b_1 _13493_ (.A(_03119_),
    .B_N(_03120_),
    .Y(_03131_));
 sg13g2_xnor2_1 _13494_ (.Y(_03132_),
    .A(_03127_),
    .B(_03131_));
 sg13g2_xnor2_1 _13495_ (.Y(_03133_),
    .A(_02992_),
    .B(_03000_));
 sg13g2_xnor2_1 _13496_ (.Y(_03134_),
    .A(_03008_),
    .B(_03133_));
 sg13g2_nand2_1 _13497_ (.Y(_03135_),
    .A(_03132_),
    .B(_03134_));
 sg13g2_nor2_1 _13498_ (.A(_03132_),
    .B(_03134_),
    .Y(_03136_));
 sg13g2_xnor2_1 _13499_ (.Y(_03137_),
    .A(_03132_),
    .B(_03134_));
 sg13g2_nand2_1 _13500_ (.Y(_03138_),
    .A(_02967_),
    .B(_02979_));
 sg13g2_a21oi_1 _13501_ (.A1(_02892_),
    .A2(_02898_),
    .Y(_03139_),
    .B1(_02910_));
 sg13g2_nor2_2 _13502_ (.A(_02899_),
    .B(_03139_),
    .Y(_03140_));
 sg13g2_nand2b_1 _13503_ (.Y(_03141_),
    .B(_02845_),
    .A_N(_03140_));
 sg13g2_nor2b_1 _13504_ (.A(_02845_),
    .B_N(_03140_),
    .Y(_03142_));
 sg13g2_xnor2_1 _13505_ (.Y(_03143_),
    .A(_02845_),
    .B(_03140_));
 sg13g2_xnor2_1 _13506_ (.Y(_03144_),
    .A(_03138_),
    .B(_03143_));
 sg13g2_a21o_1 _13507_ (.A2(_02939_),
    .A1(_02932_),
    .B1(_02948_),
    .X(_03145_));
 sg13g2_o21ai_1 _13508_ (.B1(_03145_),
    .Y(_03146_),
    .A1(_02932_),
    .A2(_02939_));
 sg13g2_nor3_1 _13509_ (.A(_02585_),
    .B(_02590_),
    .C(_03146_),
    .Y(_03147_));
 sg13g2_o21ai_1 _13510_ (.B1(_03146_),
    .Y(_03148_),
    .A1(_02585_),
    .A2(_02590_));
 sg13g2_nor2b_1 _13511_ (.A(_03147_),
    .B_N(_03148_),
    .Y(_03149_));
 sg13g2_xnor2_1 _13512_ (.Y(_03150_),
    .A(_02603_),
    .B(_03149_));
 sg13g2_nand2_1 _13513_ (.Y(_03151_),
    .A(_03144_),
    .B(_03150_));
 sg13g2_nor2_1 _13514_ (.A(_02626_),
    .B(_02631_),
    .Y(_03152_));
 sg13g2_nor3_1 _13515_ (.A(_02619_),
    .B(_02627_),
    .C(_03152_),
    .Y(_03153_));
 sg13g2_o21ai_1 _13516_ (.B1(_02619_),
    .Y(_03154_),
    .A1(_02627_),
    .A2(_03152_));
 sg13g2_nor2b_1 _13517_ (.A(_03153_),
    .B_N(_03154_),
    .Y(_03155_));
 sg13g2_xnor2_1 _13518_ (.Y(_03156_),
    .A(_02644_),
    .B(_03155_));
 sg13g2_nor2_1 _13519_ (.A(_03144_),
    .B(_03150_),
    .Y(_03157_));
 sg13g2_a21oi_2 _13520_ (.B1(_03157_),
    .Y(_03158_),
    .A2(_03156_),
    .A1(_03151_));
 sg13g2_a21oi_1 _13521_ (.A1(_03156_),
    .A2(_03157_),
    .Y(_03159_),
    .B1(_03158_));
 sg13g2_nor2_1 _13522_ (.A(_03151_),
    .B(_03156_),
    .Y(_03160_));
 sg13g2_nor2_2 _13523_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 sg13g2_xnor2_1 _13524_ (.Y(_03162_),
    .A(_03137_),
    .B(_03161_));
 sg13g2_nand2_1 _13525_ (.Y(_03163_),
    .A(_03070_),
    .B(_03071_));
 sg13g2_xnor2_1 _13526_ (.Y(_03164_),
    .A(_03099_),
    .B(_03163_));
 sg13g2_inv_1 _13527_ (.Y(_03165_),
    .A(_03164_));
 sg13g2_nand2_1 _13528_ (.Y(_03166_),
    .A(_03162_),
    .B(_03165_));
 sg13g2_xnor2_1 _13529_ (.Y(_03167_),
    .A(_03162_),
    .B(_03165_));
 sg13g2_nand2_1 _13530_ (.Y(_03168_),
    .A(_02813_),
    .B(_02820_));
 sg13g2_nand2b_2 _13531_ (.Y(_03169_),
    .B(_03168_),
    .A_N(_02819_));
 sg13g2_o21ai_1 _13532_ (.B1(_02951_),
    .Y(_03170_),
    .A1(net2803),
    .A2(_02954_));
 sg13g2_nand3_1 _13533_ (.B(_03169_),
    .C(_03170_),
    .A(_02955_),
    .Y(_03171_));
 sg13g2_a21o_1 _13534_ (.A2(_03170_),
    .A1(_02955_),
    .B1(_03169_),
    .X(_03172_));
 sg13g2_nand2_1 _13535_ (.Y(_03173_),
    .A(_03171_),
    .B(_03172_));
 sg13g2_o21ai_1 _13536_ (.B1(_02965_),
    .Y(_03174_),
    .A1(_02959_),
    .A2(_02960_));
 sg13g2_nand2_1 _13537_ (.Y(_03175_),
    .A(_02961_),
    .B(_03174_));
 sg13g2_xor2_1 _13538_ (.B(_03175_),
    .A(_03173_),
    .X(_03176_));
 sg13g2_nand2b_1 _13539_ (.Y(_03177_),
    .B(_02828_),
    .A_N(_02824_));
 sg13g2_a22oi_1 _13540_ (.Y(_03178_),
    .B1(_03177_),
    .B2(_02827_),
    .A2(_02909_),
    .A1(_02904_));
 sg13g2_nand4_1 _13541_ (.B(_02904_),
    .C(_02909_),
    .A(_02827_),
    .Y(_03179_),
    .D(_03177_));
 sg13g2_nand2b_1 _13542_ (.Y(_03180_),
    .B(_03179_),
    .A_N(_03178_));
 sg13g2_a21oi_2 _13543_ (.B1(_02840_),
    .Y(_03181_),
    .A2(_02839_),
    .A1(_02833_));
 sg13g2_xnor2_1 _13544_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_nand2_1 _13545_ (.Y(_03183_),
    .A(_03176_),
    .B(_03182_));
 sg13g2_xnor2_1 _13546_ (.Y(_03184_),
    .A(_03176_),
    .B(_03182_));
 sg13g2_o21ai_1 _13547_ (.B1(_02935_),
    .Y(_03185_),
    .A1(_02703_),
    .A2(_02936_));
 sg13g2_o21ai_1 _13548_ (.B1(_02975_),
    .Y(_03186_),
    .A1(_02973_),
    .A2(_02977_));
 sg13g2_nand2b_1 _13549_ (.Y(_03187_),
    .B(_03186_),
    .A_N(_03185_));
 sg13g2_nor2b_1 _13550_ (.A(_03186_),
    .B_N(_03185_),
    .Y(_03188_));
 sg13g2_xnor2_1 _13551_ (.Y(_03189_),
    .A(_03185_),
    .B(_03186_));
 sg13g2_xnor2_1 _13552_ (.Y(_03190_),
    .A(_02930_),
    .B(_03189_));
 sg13g2_xnor2_1 _13553_ (.Y(_03191_),
    .A(_03184_),
    .B(_03190_));
 sg13g2_o21ai_1 _13554_ (.B1(_03191_),
    .Y(_03192_),
    .A1(_03162_),
    .A2(_03165_));
 sg13g2_xnor2_1 _13555_ (.Y(_03193_),
    .A(_03167_),
    .B(_03191_));
 sg13g2_o21ai_1 _13556_ (.B1(_02941_),
    .Y(_03194_),
    .A1(_02942_),
    .A2(_02945_));
 sg13g2_nand2_2 _13557_ (.Y(_03195_),
    .A(_02946_),
    .B(_03194_));
 sg13g2_nand2_1 _13558_ (.Y(_03196_),
    .A(_03166_),
    .B(_03192_));
 sg13g2_nor3_1 _13559_ (.A(_03193_),
    .B(_03195_),
    .C(_03196_),
    .Y(_03197_));
 sg13g2_or3_1 _13560_ (.A(_03193_),
    .B(_03195_),
    .C(_03196_),
    .X(_03198_));
 sg13g2_o21ai_1 _13561_ (.B1(_03196_),
    .Y(_03199_),
    .A1(_03193_),
    .A2(_03195_));
 sg13g2_o21ai_1 _13562_ (.B1(_03135_),
    .Y(_03200_),
    .A1(_03136_),
    .A2(_03161_));
 sg13g2_a21o_1 _13563_ (.A2(_03199_),
    .A1(_03198_),
    .B1(_03200_),
    .X(_03201_));
 sg13g2_nand3_1 _13564_ (.B(_03199_),
    .C(_03200_),
    .A(_03198_),
    .Y(_03202_));
 sg13g2_nand3_1 _13565_ (.B(_03201_),
    .C(_03202_),
    .A(_03130_),
    .Y(_03203_));
 sg13g2_a21oi_1 _13566_ (.A1(_03201_),
    .A2(_03202_),
    .Y(_03204_),
    .B1(_03130_));
 sg13g2_a21o_1 _13567_ (.A2(_03202_),
    .A1(_03201_),
    .B1(_03130_),
    .X(_03205_));
 sg13g2_nand2_1 _13568_ (.Y(_03206_),
    .A(_03033_),
    .B(_03041_));
 sg13g2_a21oi_1 _13569_ (.A1(_03032_),
    .A2(_03206_),
    .Y(_03207_),
    .B1(_03158_));
 sg13g2_nand3_1 _13570_ (.B(_03158_),
    .C(_03206_),
    .A(_03032_),
    .Y(_03208_));
 sg13g2_nor2b_1 _13571_ (.A(_03207_),
    .B_N(_03208_),
    .Y(_03209_));
 sg13g2_a21oi_1 _13572_ (.A1(_03057_),
    .A2(_03068_),
    .Y(_03210_),
    .B1(_03058_));
 sg13g2_xnor2_1 _13573_ (.Y(_03211_),
    .A(_03209_),
    .B(_03210_));
 sg13g2_inv_1 _13574_ (.Y(_03212_),
    .A(_03211_));
 sg13g2_and3_1 _13575_ (.X(_03213_),
    .A(_03203_),
    .B(_03205_),
    .C(_03212_));
 sg13g2_a21oi_1 _13576_ (.A1(_03203_),
    .A2(_03205_),
    .Y(_03214_),
    .B1(_03212_));
 sg13g2_o21ai_1 _13577_ (.B1(_03097_),
    .Y(_03215_),
    .A1(_03080_),
    .A2(_03089_));
 sg13g2_o21ai_1 _13578_ (.B1(_03190_),
    .Y(_03216_),
    .A1(_03176_),
    .A2(_03182_));
 sg13g2_nand2_1 _13579_ (.Y(_03217_),
    .A(_03183_),
    .B(_03216_));
 sg13g2_nand2_1 _13580_ (.Y(_03218_),
    .A(_03215_),
    .B(_03217_));
 sg13g2_or2_1 _13581_ (.X(_03219_),
    .B(_03217_),
    .A(_03215_));
 sg13g2_and2_1 _13582_ (.A(_03218_),
    .B(_03219_),
    .X(_03220_));
 sg13g2_xnor2_1 _13583_ (.Y(_03221_),
    .A(_02991_),
    .B(_03220_));
 sg13g2_nor2_1 _13584_ (.A(_02500_),
    .B(_03116_),
    .Y(_03222_));
 sg13g2_nor2_2 _13585_ (.A(_03115_),
    .B(_03222_),
    .Y(_03223_));
 sg13g2_nand3_1 _13586_ (.B(_03002_),
    .C(_03007_),
    .A(_02999_),
    .Y(_03224_));
 sg13g2_a21o_1 _13587_ (.A2(_03007_),
    .A1(_03002_),
    .B1(_02999_),
    .X(_03225_));
 sg13g2_nand2_1 _13588_ (.Y(_03226_),
    .A(_03224_),
    .B(_03225_));
 sg13g2_xor2_1 _13589_ (.B(_03226_),
    .A(_03223_),
    .X(_03227_));
 sg13g2_nand2_1 _13590_ (.Y(_03228_),
    .A(_03221_),
    .B(_03227_));
 sg13g2_or2_1 _13591_ (.X(_03229_),
    .B(_03227_),
    .A(_03221_));
 sg13g2_nand2_1 _13592_ (.Y(_03230_),
    .A(_03228_),
    .B(_03229_));
 sg13g2_a21oi_2 _13593_ (.B1(_03142_),
    .Y(_03231_),
    .A2(_03141_),
    .A1(_03138_));
 sg13g2_a21oi_2 _13594_ (.B1(_03124_),
    .Y(_03232_),
    .A2(_03126_),
    .A1(_03123_));
 sg13g2_nor3_1 _13595_ (.A(_03107_),
    .B(_03110_),
    .C(_03232_),
    .Y(_03233_));
 sg13g2_o21ai_1 _13596_ (.B1(_03232_),
    .Y(_03234_),
    .A1(_03107_),
    .A2(_03110_));
 sg13g2_or2_1 _13597_ (.X(_03235_),
    .B(_03234_),
    .A(_03231_));
 sg13g2_a21oi_2 _13598_ (.B1(_03233_),
    .Y(_03236_),
    .A2(_03234_),
    .A1(_03231_));
 sg13g2_a22oi_1 _13599_ (.Y(_03237_),
    .B1(_03235_),
    .B2(_03236_),
    .A2(_03233_),
    .A1(_03231_));
 sg13g2_xor2_1 _13600_ (.B(_03237_),
    .A(_03230_),
    .X(_03238_));
 sg13g2_nor3_1 _13601_ (.A(_03213_),
    .B(_03214_),
    .C(_03238_),
    .Y(_03239_));
 sg13g2_o21ai_1 _13602_ (.B1(_03238_),
    .Y(_03240_),
    .A1(_03213_),
    .A2(_03214_));
 sg13g2_a21oi_2 _13603_ (.B1(_03027_),
    .Y(_03241_),
    .A2(_03030_),
    .A1(_03026_));
 sg13g2_a21oi_2 _13604_ (.B1(_03153_),
    .Y(_03242_),
    .A2(_03154_),
    .A1(_02644_));
 sg13g2_a21oi_1 _13605_ (.A1(_02604_),
    .A2(_03148_),
    .Y(_03243_),
    .B1(_03147_));
 sg13g2_or2_2 _13606_ (.X(_03244_),
    .B(_03243_),
    .A(_03242_));
 sg13g2_nand2_2 _13607_ (.Y(_03245_),
    .A(_03242_),
    .B(_03243_));
 sg13g2_nand2_1 _13608_ (.Y(_03246_),
    .A(_03244_),
    .B(_03245_));
 sg13g2_xor2_1 _13609_ (.B(_03246_),
    .A(_03241_),
    .X(_03247_));
 sg13g2_nand2_1 _13610_ (.Y(_03248_),
    .A(_03020_),
    .B(_03040_));
 sg13g2_xnor2_1 _13611_ (.Y(_03249_),
    .A(_03020_),
    .B(_03040_));
 sg13g2_o21ai_1 _13612_ (.B1(_03045_),
    .Y(_03250_),
    .A1(_03046_),
    .A2(_03048_));
 sg13g2_xor2_1 _13613_ (.B(_03250_),
    .A(_03249_),
    .X(_03251_));
 sg13g2_nor2_1 _13614_ (.A(_03247_),
    .B(_03251_),
    .Y(_03252_));
 sg13g2_and2_1 _13615_ (.A(_03247_),
    .B(_03251_),
    .X(_03253_));
 sg13g2_nor2_1 _13616_ (.A(_03252_),
    .B(_03253_),
    .Y(_03254_));
 sg13g2_a21oi_2 _13617_ (.B1(_03052_),
    .Y(_03255_),
    .A2(_03055_),
    .A1(_03053_));
 sg13g2_nand2_1 _13618_ (.Y(_03256_),
    .A(_03066_),
    .B(_03255_));
 sg13g2_xor2_1 _13619_ (.B(_03255_),
    .A(_03066_),
    .X(_03257_));
 sg13g2_xnor2_1 _13620_ (.Y(_03258_),
    .A(_03079_),
    .B(_03257_));
 sg13g2_xor2_1 _13621_ (.B(_03258_),
    .A(_03254_),
    .X(_03259_));
 sg13g2_inv_1 _13622_ (.Y(_03260_),
    .A(_03259_));
 sg13g2_o21ai_1 _13623_ (.B1(_03240_),
    .Y(_03261_),
    .A1(_03239_),
    .A2(_03260_));
 sg13g2_nand2b_1 _13624_ (.Y(_03262_),
    .B(_03259_),
    .A_N(_03240_));
 sg13g2_nand2_1 _13625_ (.Y(_03263_),
    .A(_03239_),
    .B(_03260_));
 sg13g2_nand2_1 _13626_ (.Y(_03264_),
    .A(_03261_),
    .B(_03262_));
 sg13g2_nand2_1 _13627_ (.Y(_03265_),
    .A(_03263_),
    .B(_03264_));
 sg13g2_a21oi_2 _13628_ (.B1(_03094_),
    .Y(_03266_),
    .A2(_03093_),
    .A1(_02891_));
 sg13g2_nand3_1 _13629_ (.B(_03088_),
    .C(_03266_),
    .A(_03084_),
    .Y(_03267_));
 sg13g2_a21o_1 _13630_ (.A2(_03088_),
    .A1(_03084_),
    .B1(_03266_),
    .X(_03268_));
 sg13g2_nand2_1 _13631_ (.Y(_03269_),
    .A(_03267_),
    .B(_03268_));
 sg13g2_o21ai_1 _13632_ (.B1(_03179_),
    .Y(_03270_),
    .A1(_03178_),
    .A2(_03181_));
 sg13g2_xor2_1 _13633_ (.B(_03270_),
    .A(_03269_),
    .X(_03271_));
 sg13g2_nand2_1 _13634_ (.Y(_03272_),
    .A(_03171_),
    .B(_03175_));
 sg13g2_nand2_1 _13635_ (.Y(_03273_),
    .A(_03172_),
    .B(_03272_));
 sg13g2_nand3_1 _13636_ (.B(_03271_),
    .C(_03272_),
    .A(_03172_),
    .Y(_03274_));
 sg13g2_nor2b_1 _13637_ (.A(_03271_),
    .B_N(_03273_),
    .Y(_03275_));
 sg13g2_xnor2_1 _13638_ (.Y(_03276_),
    .A(_03271_),
    .B(_03273_));
 sg13g2_o21ai_1 _13639_ (.B1(_03187_),
    .Y(_03277_),
    .A1(_02930_),
    .A2(_03188_));
 sg13g2_inv_1 _13640_ (.Y(_03278_),
    .A(_03277_));
 sg13g2_xnor2_1 _13641_ (.Y(_03279_),
    .A(_03276_),
    .B(_03277_));
 sg13g2_a21o_1 _13642_ (.A2(_03279_),
    .A1(_03263_),
    .B1(_03261_),
    .X(_03280_));
 sg13g2_a21oi_1 _13643_ (.A1(_03203_),
    .A2(_03212_),
    .Y(_03281_),
    .B1(_03204_));
 sg13g2_nand2_1 _13644_ (.Y(_03282_),
    .A(_03280_),
    .B(_03281_));
 sg13g2_nand2b_1 _13645_ (.Y(_03283_),
    .B(_03279_),
    .A_N(_03262_));
 sg13g2_nand2_1 _13646_ (.Y(_03284_),
    .A(_03282_),
    .B(_03283_));
 sg13g2_nand2_1 _13647_ (.Y(_03285_),
    .A(_03229_),
    .B(_03237_));
 sg13g2_nor2_1 _13648_ (.A(_03253_),
    .B(_03258_),
    .Y(_03286_));
 sg13g2_nor2_1 _13649_ (.A(_03252_),
    .B(_03286_),
    .Y(_03287_));
 sg13g2_a21oi_1 _13650_ (.A1(_03228_),
    .A2(_03285_),
    .Y(_03288_),
    .B1(_03287_));
 sg13g2_nand3_1 _13651_ (.B(_03285_),
    .C(_03287_),
    .A(_03228_),
    .Y(_03289_));
 sg13g2_a21oi_2 _13652_ (.B1(_03275_),
    .Y(_03290_),
    .A2(_03278_),
    .A1(_03274_));
 sg13g2_o21ai_1 _13653_ (.B1(_03289_),
    .Y(_03291_),
    .A1(_03288_),
    .A2(_03290_));
 sg13g2_nor2_1 _13654_ (.A(_03284_),
    .B(_03291_),
    .Y(_03292_));
 sg13g2_nand2_1 _13655_ (.Y(_03293_),
    .A(_03284_),
    .B(_03291_));
 sg13g2_a21oi_1 _13656_ (.A1(_03199_),
    .A2(_03200_),
    .Y(_03294_),
    .B1(_03197_));
 sg13g2_a21oi_1 _13657_ (.A1(_03102_),
    .A2(_03128_),
    .Y(_03295_),
    .B1(_03101_));
 sg13g2_and2_1 _13658_ (.A(_03294_),
    .B(_03295_),
    .X(_03296_));
 sg13g2_nor2_1 _13659_ (.A(_03294_),
    .B(_03295_),
    .Y(_03297_));
 sg13g2_a21o_1 _13660_ (.A2(_03210_),
    .A1(_03208_),
    .B1(_03207_),
    .X(_03298_));
 sg13g2_nor2_1 _13661_ (.A(_03296_),
    .B(_03298_),
    .Y(_03299_));
 sg13g2_nor2_1 _13662_ (.A(_03297_),
    .B(_03299_),
    .Y(_03300_));
 sg13g2_o21ai_1 _13663_ (.B1(_03293_),
    .Y(_03301_),
    .A1(_03292_),
    .A2(_03300_));
 sg13g2_nand2b_1 _13664_ (.Y(_03302_),
    .B(_03245_),
    .A_N(_03241_));
 sg13g2_o21ai_1 _13665_ (.B1(_03250_),
    .Y(_03303_),
    .A1(_03020_),
    .A2(_03040_));
 sg13g2_nand2_1 _13666_ (.Y(_03304_),
    .A(_03248_),
    .B(_03303_));
 sg13g2_nand3_1 _13667_ (.B(_03302_),
    .C(_03304_),
    .A(_03244_),
    .Y(_03305_));
 sg13g2_a21o_1 _13668_ (.A2(_03302_),
    .A1(_03244_),
    .B1(_03304_),
    .X(_03306_));
 sg13g2_o21ai_1 _13669_ (.B1(_03079_),
    .Y(_03307_),
    .A1(_03066_),
    .A2(_03255_));
 sg13g2_nand2_2 _13670_ (.Y(_03308_),
    .A(_03256_),
    .B(_03307_));
 sg13g2_nand2_1 _13671_ (.Y(_03309_),
    .A(_03306_),
    .B(_03308_));
 sg13g2_nand2_2 _13672_ (.Y(_03310_),
    .A(_03305_),
    .B(_03309_));
 sg13g2_inv_1 _13673_ (.Y(_03311_),
    .A(_03310_));
 sg13g2_nand2_1 _13674_ (.Y(_03312_),
    .A(_03223_),
    .B(_03224_));
 sg13g2_nand2_1 _13675_ (.Y(_03313_),
    .A(_02991_),
    .B(_03218_));
 sg13g2_and4_1 _13676_ (.A(_03219_),
    .B(_03225_),
    .C(_03312_),
    .D(_03313_),
    .X(_03314_));
 sg13g2_a22oi_1 _13677_ (.Y(_03315_),
    .B1(_03313_),
    .B2(_03219_),
    .A2(_03312_),
    .A1(_03225_));
 sg13g2_nor2_1 _13678_ (.A(_03236_),
    .B(_03314_),
    .Y(_03316_));
 sg13g2_nor2_2 _13679_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sg13g2_nand3_1 _13680_ (.B(_03281_),
    .C(_03283_),
    .A(_03280_),
    .Y(_03318_));
 sg13g2_a21o_1 _13681_ (.A2(_03283_),
    .A1(_03280_),
    .B1(_03281_),
    .X(_03319_));
 sg13g2_nor2b_1 _13682_ (.A(_03288_),
    .B_N(_03289_),
    .Y(_03320_));
 sg13g2_xnor2_1 _13683_ (.Y(_03321_),
    .A(_03290_),
    .B(_03320_));
 sg13g2_a21oi_1 _13684_ (.A1(_03318_),
    .A2(_03319_),
    .Y(_03322_),
    .B1(_03321_));
 sg13g2_a21o_1 _13685_ (.A2(_03319_),
    .A1(_03318_),
    .B1(_03321_),
    .X(_03323_));
 sg13g2_nand3_1 _13686_ (.B(_03319_),
    .C(_03321_),
    .A(_03318_),
    .Y(_03324_));
 sg13g2_nor2_1 _13687_ (.A(_03296_),
    .B(_03297_),
    .Y(_03325_));
 sg13g2_xor2_1 _13688_ (.B(_03325_),
    .A(_03298_),
    .X(_03326_));
 sg13g2_a21o_1 _13689_ (.A2(_03324_),
    .A1(_03323_),
    .B1(_03326_),
    .X(_03327_));
 sg13g2_nand3b_1 _13690_ (.B(_03324_),
    .C(_03326_),
    .Y(_03328_),
    .A_N(_03322_));
 sg13g2_nor2_1 _13691_ (.A(_03314_),
    .B(_03315_),
    .Y(_03329_));
 sg13g2_xnor2_1 _13692_ (.Y(_03330_),
    .A(_03236_),
    .B(_03329_));
 sg13g2_nand2_1 _13693_ (.Y(_03331_),
    .A(_03305_),
    .B(_03306_));
 sg13g2_xor2_1 _13694_ (.B(_03331_),
    .A(_03308_),
    .X(_03332_));
 sg13g2_nand2_1 _13695_ (.Y(_03333_),
    .A(_03330_),
    .B(_03332_));
 sg13g2_nor2_1 _13696_ (.A(_03330_),
    .B(_03332_),
    .Y(_03334_));
 sg13g2_xnor2_1 _13697_ (.Y(_03335_),
    .A(_03330_),
    .B(_03332_));
 sg13g2_nand2_1 _13698_ (.Y(_03336_),
    .A(_03267_),
    .B(_03270_));
 sg13g2_and2_2 _13699_ (.A(_03268_),
    .B(_03336_),
    .X(_03337_));
 sg13g2_xnor2_1 _13700_ (.Y(_03338_),
    .A(_03335_),
    .B(_03337_));
 sg13g2_a21oi_2 _13701_ (.B1(_03338_),
    .Y(_03339_),
    .A2(_03328_),
    .A1(_03327_));
 sg13g2_o21ai_1 _13702_ (.B1(_03324_),
    .Y(_03340_),
    .A1(_03322_),
    .A2(_03326_));
 sg13g2_nor3_1 _13703_ (.A(_03324_),
    .B(_03326_),
    .C(_03338_),
    .Y(_03341_));
 sg13g2_xor2_1 _13704_ (.B(_03340_),
    .A(_03339_),
    .X(_03342_));
 sg13g2_a21oi_2 _13705_ (.B1(_03334_),
    .Y(_03343_),
    .A2(_03337_),
    .A1(_03333_));
 sg13g2_o21ai_1 _13706_ (.B1(_03343_),
    .Y(_03344_),
    .A1(_03339_),
    .A2(_03340_));
 sg13g2_xnor2_1 _13707_ (.Y(_03345_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_nor2b_1 _13708_ (.A(_03292_),
    .B_N(_03293_),
    .Y(_03346_));
 sg13g2_xnor2_1 _13709_ (.Y(_03347_),
    .A(_03300_),
    .B(_03346_));
 sg13g2_inv_1 _13710_ (.Y(_03348_),
    .A(_03347_));
 sg13g2_xnor2_1 _13711_ (.Y(_03349_),
    .A(_03345_),
    .B(_03347_));
 sg13g2_a21o_1 _13712_ (.A2(_03348_),
    .A1(_03345_),
    .B1(_03317_),
    .X(_03350_));
 sg13g2_xnor2_1 _13713_ (.Y(_03351_),
    .A(_03317_),
    .B(_03349_));
 sg13g2_o21ai_1 _13714_ (.B1(_03350_),
    .Y(_03352_),
    .A1(_03345_),
    .A2(_03348_));
 sg13g2_nor4_1 _13715_ (.A(_03310_),
    .B(_03317_),
    .C(_03345_),
    .D(_03348_),
    .Y(_03353_));
 sg13g2_inv_1 _13716_ (.Y(_03354_),
    .A(_03353_));
 sg13g2_a21o_1 _13717_ (.A2(_03351_),
    .A1(_03311_),
    .B1(_03352_),
    .X(_03355_));
 sg13g2_nand2b_1 _13718_ (.Y(_03356_),
    .B(_03344_),
    .A_N(_03341_));
 sg13g2_a21o_1 _13719_ (.A2(_03355_),
    .A1(_03354_),
    .B1(_03356_),
    .X(_03357_));
 sg13g2_nand3_1 _13720_ (.B(_03355_),
    .C(_03356_),
    .A(_03354_),
    .Y(_03358_));
 sg13g2_and3_2 _13721_ (.X(_03359_),
    .A(_03301_),
    .B(_03357_),
    .C(_03358_));
 sg13g2_a21oi_1 _13722_ (.A1(_03355_),
    .A2(_03356_),
    .Y(_03360_),
    .B1(_03353_));
 sg13g2_nand2b_2 _13723_ (.Y(_03361_),
    .B(_03360_),
    .A_N(_03359_));
 sg13g2_a21oi_2 _13724_ (.B1(_02284_),
    .Y(_03362_),
    .A2(_02285_),
    .A1(_02264_));
 sg13g2_o21ai_1 _13725_ (.B1(_02349_),
    .Y(_03363_),
    .A1(_02329_),
    .A2(_02350_));
 sg13g2_a21oi_2 _13726_ (.B1(_02453_),
    .Y(_03364_),
    .A2(_02454_),
    .A1(_02431_));
 sg13g2_a21o_1 _13727_ (.A2(_03363_),
    .A1(_03362_),
    .B1(_03364_),
    .X(_03365_));
 sg13g2_o21ai_1 _13728_ (.B1(_03365_),
    .Y(_03366_),
    .A1(_03362_),
    .A2(_03363_));
 sg13g2_o21ai_1 _13729_ (.B1(_02068_),
    .Y(_03367_),
    .A1(_01994_),
    .A2(_02069_));
 sg13g2_nand2_1 _13730_ (.Y(_03368_),
    .A(_02144_),
    .B(_03367_));
 sg13g2_or2_1 _13731_ (.X(_03369_),
    .B(_03367_),
    .A(_02144_));
 sg13g2_nand2_1 _13732_ (.Y(_03370_),
    .A(_02295_),
    .B(_02313_));
 sg13g2_nand2_1 _13733_ (.Y(_03371_),
    .A(_02314_),
    .B(_03370_));
 sg13g2_nand2b_1 _13734_ (.Y(_03372_),
    .B(_03369_),
    .A_N(_03371_));
 sg13g2_nand2_1 _13735_ (.Y(_03373_),
    .A(_02287_),
    .B(_02354_));
 sg13g2_nor2_1 _13736_ (.A(_02389_),
    .B(_02457_),
    .Y(_03374_));
 sg13g2_a21oi_1 _13737_ (.A1(_02424_),
    .A2(_02456_),
    .Y(_03375_),
    .B1(_03374_));
 sg13g2_a21oi_1 _13738_ (.A1(_02353_),
    .A2(_03373_),
    .Y(_03376_),
    .B1(_03375_));
 sg13g2_and3_1 _13739_ (.X(_03377_),
    .A(_02353_),
    .B(_03373_),
    .C(_03375_));
 sg13g2_nor2_1 _13740_ (.A(_02255_),
    .B(_03376_),
    .Y(_03378_));
 sg13g2_nor2_1 _13741_ (.A(_03377_),
    .B(_03378_),
    .Y(_03379_));
 sg13g2_and3_1 _13742_ (.X(_03380_),
    .A(_03368_),
    .B(_03372_),
    .C(_03379_));
 sg13g2_inv_1 _13743_ (.Y(_03381_),
    .A(_03380_));
 sg13g2_a21oi_1 _13744_ (.A1(_03368_),
    .A2(_03372_),
    .Y(_03382_),
    .B1(_03379_));
 sg13g2_nor2_1 _13745_ (.A(_03380_),
    .B(_03382_),
    .Y(_03383_));
 sg13g2_xnor2_1 _13746_ (.Y(_03384_),
    .A(_03366_),
    .B(_03383_));
 sg13g2_a21o_1 _13747_ (.A2(_02461_),
    .A1(_02256_),
    .B1(_02460_),
    .X(_03385_));
 sg13g2_a21oi_1 _13748_ (.A1(_02147_),
    .A2(_02463_),
    .Y(_03386_),
    .B1(_03385_));
 sg13g2_nand3_1 _13749_ (.B(_02256_),
    .C(_02460_),
    .A(_02147_),
    .Y(_03387_));
 sg13g2_nand2b_1 _13750_ (.Y(_03388_),
    .B(_03387_),
    .A_N(_02146_));
 sg13g2_nor2b_1 _13751_ (.A(_03386_),
    .B_N(_03388_),
    .Y(_03389_));
 sg13g2_o21ai_1 _13752_ (.B1(_01969_),
    .Y(_03390_),
    .A1(_01963_),
    .A2(_01967_));
 sg13g2_nand2_1 _13753_ (.Y(_03391_),
    .A(_02031_),
    .B(_02035_));
 sg13g2_nand2_1 _13754_ (.Y(_03392_),
    .A(_02036_),
    .B(_03391_));
 sg13g2_nand2_1 _13755_ (.Y(_03393_),
    .A(_01974_),
    .B(_01980_));
 sg13g2_and2_2 _13756_ (.A(_01979_),
    .B(_03393_),
    .X(_03394_));
 sg13g2_xor2_1 _13757_ (.B(_03394_),
    .A(_03392_),
    .X(_03395_));
 sg13g2_a21o_1 _13758_ (.A2(_03394_),
    .A1(_03392_),
    .B1(_03390_),
    .X(_03396_));
 sg13g2_o21ai_1 _13759_ (.B1(_03396_),
    .Y(_03397_),
    .A1(_03392_),
    .A2(_03394_));
 sg13g2_xnor2_1 _13760_ (.Y(_03398_),
    .A(_03390_),
    .B(_03395_));
 sg13g2_nor2_1 _13761_ (.A(_02120_),
    .B(_02126_),
    .Y(_03399_));
 sg13g2_nor2_1 _13762_ (.A(_02125_),
    .B(_03399_),
    .Y(_03400_));
 sg13g2_nand2b_1 _13763_ (.Y(_03401_),
    .B(_01991_),
    .A_N(_01985_));
 sg13g2_nand2_1 _13764_ (.Y(_03402_),
    .A(_02129_),
    .B(_02133_));
 sg13g2_a22oi_1 _13765_ (.Y(_03403_),
    .B1(_03402_),
    .B2(_02132_),
    .A2(_03401_),
    .A1(_01990_));
 sg13g2_nand4_1 _13766_ (.B(_02132_),
    .C(_03401_),
    .A(_01990_),
    .Y(_03404_),
    .D(_03402_));
 sg13g2_nor2b_1 _13767_ (.A(_03403_),
    .B_N(_03404_),
    .Y(_03405_));
 sg13g2_xnor2_1 _13768_ (.Y(_03406_),
    .A(_03400_),
    .B(_03405_));
 sg13g2_nand2_1 _13769_ (.Y(_03407_),
    .A(_03398_),
    .B(_03406_));
 sg13g2_or2_1 _13770_ (.X(_03408_),
    .B(_03406_),
    .A(_03398_));
 sg13g2_nand2_1 _13771_ (.Y(_03409_),
    .A(_02076_),
    .B(_02080_));
 sg13g2_nand2b_2 _13772_ (.Y(_03410_),
    .B(_03409_),
    .A_N(_02079_));
 sg13g2_a21oi_2 _13773_ (.B1(_02115_),
    .Y(_03411_),
    .A2(_02114_),
    .A1(_02110_));
 sg13g2_nand2_1 _13774_ (.Y(_03412_),
    .A(_02085_),
    .B(_02089_));
 sg13g2_nand2_1 _13775_ (.Y(_03413_),
    .A(_02090_),
    .B(_03412_));
 sg13g2_nand2_1 _13776_ (.Y(_03414_),
    .A(_03411_),
    .B(_03413_));
 sg13g2_or2_1 _13777_ (.X(_03415_),
    .B(_03413_),
    .A(_03411_));
 sg13g2_inv_1 _13778_ (.Y(_03416_),
    .A(_03415_));
 sg13g2_nand2_1 _13779_ (.Y(_03417_),
    .A(_03414_),
    .B(_03415_));
 sg13g2_xor2_1 _13780_ (.B(_03417_),
    .A(_03410_),
    .X(_03418_));
 sg13g2_nand2_1 _13781_ (.Y(_03419_),
    .A(_03408_),
    .B(_03418_));
 sg13g2_nand2_1 _13782_ (.Y(_03420_),
    .A(_03407_),
    .B(_03419_));
 sg13g2_o21ai_1 _13783_ (.B1(_02022_),
    .Y(_03421_),
    .A1(_02018_),
    .A2(_02023_));
 sg13g2_o21ai_1 _13784_ (.B1(_02012_),
    .Y(_03422_),
    .A1(_02007_),
    .A2(_02013_));
 sg13g2_and2_1 _13785_ (.A(_02158_),
    .B(_03422_),
    .X(_03423_));
 sg13g2_or2_1 _13786_ (.X(_03424_),
    .B(_03422_),
    .A(_02158_));
 sg13g2_a21oi_2 _13787_ (.B1(_03423_),
    .Y(_03425_),
    .A2(_03424_),
    .A1(_03421_));
 sg13g2_inv_1 _13788_ (.Y(_03426_),
    .A(_03425_));
 sg13g2_a21o_1 _13789_ (.A2(_03423_),
    .A1(_03421_),
    .B1(_03425_),
    .X(_03427_));
 sg13g2_o21ai_1 _13790_ (.B1(_03427_),
    .Y(_03428_),
    .A1(_03421_),
    .A2(_03424_));
 sg13g2_nand2_1 _13791_ (.Y(_03429_),
    .A(_02185_),
    .B(_02191_));
 sg13g2_nand2_2 _13792_ (.Y(_03430_),
    .A(_02190_),
    .B(_03429_));
 sg13g2_nand2_1 _13793_ (.Y(_03431_),
    .A(_02168_),
    .B(_02174_));
 sg13g2_nand2_2 _13794_ (.Y(_03432_),
    .A(_02173_),
    .B(_03431_));
 sg13g2_or2_1 _13795_ (.X(_03433_),
    .B(_03432_),
    .A(_03430_));
 sg13g2_and2_1 _13796_ (.A(_03430_),
    .B(_03432_),
    .X(_03434_));
 sg13g2_xor2_1 _13797_ (.B(_03432_),
    .A(_03430_),
    .X(_03435_));
 sg13g2_a21o_1 _13798_ (.A2(_02164_),
    .A1(_02161_),
    .B1(_02160_),
    .X(_03436_));
 sg13g2_o21ai_1 _13799_ (.B1(_03436_),
    .Y(_03437_),
    .A1(_02161_),
    .A2(_02164_));
 sg13g2_xnor2_1 _13800_ (.Y(_03438_),
    .A(_03435_),
    .B(_03437_));
 sg13g2_nand2_1 _13801_ (.Y(_03439_),
    .A(_03428_),
    .B(_03438_));
 sg13g2_or2_1 _13802_ (.X(_03440_),
    .B(_03438_),
    .A(_03428_));
 sg13g2_a21oi_1 _13803_ (.A1(_02056_),
    .A2(_02059_),
    .Y(_03441_),
    .B1(_02052_));
 sg13g2_nor2_2 _13804_ (.A(_02060_),
    .B(_03441_),
    .Y(_03442_));
 sg13g2_a21oi_2 _13805_ (.B1(_02045_),
    .Y(_03443_),
    .A2(_02046_),
    .A1(_02039_));
 sg13g2_a21o_1 _13806_ (.A2(_01996_),
    .A1(_01995_),
    .B1(_02002_),
    .X(_03444_));
 sg13g2_inv_1 _13807_ (.Y(_03445_),
    .A(_03444_));
 sg13g2_o21ai_1 _13808_ (.B1(_03443_),
    .Y(_03446_),
    .A1(_02003_),
    .A2(_03445_));
 sg13g2_or3_1 _13809_ (.A(_02003_),
    .B(_03443_),
    .C(_03445_),
    .X(_03447_));
 sg13g2_nand2_1 _13810_ (.Y(_03448_),
    .A(_03446_),
    .B(_03447_));
 sg13g2_xnor2_1 _13811_ (.Y(_03449_),
    .A(_03442_),
    .B(_03448_));
 sg13g2_nand2_1 _13812_ (.Y(_03450_),
    .A(_03439_),
    .B(_03449_));
 sg13g2_nand3_1 _13813_ (.B(_03440_),
    .C(_03450_),
    .A(_03420_),
    .Y(_03451_));
 sg13g2_a21o_1 _13814_ (.A2(_03450_),
    .A1(_03440_),
    .B1(_03420_),
    .X(_03452_));
 sg13g2_and2_1 _13815_ (.A(_03451_),
    .B(_03452_),
    .X(_03453_));
 sg13g2_xnor2_1 _13816_ (.Y(_03454_),
    .A(_03389_),
    .B(_03453_));
 sg13g2_nand2_1 _13817_ (.Y(_03455_),
    .A(_03384_),
    .B(_03454_));
 sg13g2_or2_1 _13818_ (.X(_03456_),
    .B(_03454_),
    .A(_03384_));
 sg13g2_a21oi_1 _13819_ (.A1(_01971_),
    .A2(_01982_),
    .Y(_03457_),
    .B1(_01993_));
 sg13g2_nor2_1 _13820_ (.A(_01983_),
    .B(_03457_),
    .Y(_03458_));
 sg13g2_nand2_1 _13821_ (.Y(_03459_),
    .A(_02065_),
    .B(_03458_));
 sg13g2_nor2_1 _13822_ (.A(_02065_),
    .B(_03458_),
    .Y(_03460_));
 sg13g2_a21oi_2 _13823_ (.B1(_03460_),
    .Y(_03461_),
    .A2(_03459_),
    .A1(_02139_));
 sg13g2_a21o_1 _13824_ (.A2(_02422_),
    .A1(_02399_),
    .B1(_02421_),
    .X(_03462_));
 sg13g2_a21oi_2 _13825_ (.B1(_02386_),
    .Y(_03463_),
    .A2(_02387_),
    .A1(_02367_));
 sg13g2_nor2_1 _13826_ (.A(_03462_),
    .B(_03463_),
    .Y(_03464_));
 sg13g2_o21ai_1 _13827_ (.B1(_02247_),
    .Y(_03465_),
    .A1(_02226_),
    .A2(_02248_));
 sg13g2_nor2b_1 _13828_ (.A(_03464_),
    .B_N(_03465_),
    .Y(_03466_));
 sg13g2_a21oi_1 _13829_ (.A1(_03462_),
    .A2(_03463_),
    .Y(_03467_),
    .B1(_03466_));
 sg13g2_nor2_1 _13830_ (.A(_02193_),
    .B(_02213_),
    .Y(_03468_));
 sg13g2_nor3_1 _13831_ (.A(_02181_),
    .B(_02212_),
    .C(_03468_),
    .Y(_03469_));
 sg13g2_o21ai_1 _13832_ (.B1(_02181_),
    .Y(_03470_),
    .A1(_02212_),
    .A2(_03468_));
 sg13g2_a21oi_2 _13833_ (.B1(_02026_),
    .Y(_03471_),
    .A2(_02027_),
    .A1(_02005_));
 sg13g2_nand2b_1 _13834_ (.Y(_03472_),
    .B(_03471_),
    .A_N(_03469_));
 sg13g2_a21oi_2 _13835_ (.B1(_03467_),
    .Y(_03473_),
    .A2(_03472_),
    .A1(_03470_));
 sg13g2_and3_1 _13836_ (.X(_03474_),
    .A(_03467_),
    .B(_03470_),
    .C(_03472_));
 sg13g2_inv_1 _13837_ (.Y(_03475_),
    .A(_03474_));
 sg13g2_a21oi_2 _13838_ (.B1(_03473_),
    .Y(_03476_),
    .A2(_03475_),
    .A1(_03461_));
 sg13g2_nand2b_1 _13839_ (.Y(_03477_),
    .B(_03474_),
    .A_N(_03461_));
 sg13g2_a22oi_1 _13840_ (.Y(_03478_),
    .B1(_03476_),
    .B2(_03477_),
    .A2(_03473_),
    .A1(_03461_));
 sg13g2_nand2_1 _13841_ (.Y(_03479_),
    .A(_03456_),
    .B(_03478_));
 sg13g2_nand2_1 _13842_ (.Y(_03480_),
    .A(_03455_),
    .B(_03479_));
 sg13g2_o21ai_1 _13843_ (.B1(_02396_),
    .Y(_03481_),
    .A1(_02391_),
    .A2(_02397_));
 sg13g2_a21oi_1 _13844_ (.A1(_02378_),
    .A2(_02383_),
    .Y(_03482_),
    .B1(_02382_));
 sg13g2_inv_1 _13845_ (.Y(_03483_),
    .A(_03482_));
 sg13g2_nand2_1 _13846_ (.Y(_03484_),
    .A(_03481_),
    .B(_03483_));
 sg13g2_nor2_1 _13847_ (.A(_03481_),
    .B(_03483_),
    .Y(_03485_));
 sg13g2_a21oi_2 _13848_ (.B1(_02373_),
    .Y(_03486_),
    .A2(_02374_),
    .A1(_02370_));
 sg13g2_a21oi_1 _13849_ (.A1(_03484_),
    .A2(_03486_),
    .Y(_03487_),
    .B1(_03485_));
 sg13g2_inv_1 _13850_ (.Y(_03488_),
    .A(_03487_));
 sg13g2_a21oi_1 _13851_ (.A1(_02411_),
    .A2(_02418_),
    .Y(_03489_),
    .B1(_02417_));
 sg13g2_a21o_1 _13852_ (.A2(_02429_),
    .A1(_02426_),
    .B1(_02425_),
    .X(_03490_));
 sg13g2_o21ai_1 _13853_ (.B1(_03490_),
    .Y(_03491_),
    .A1(_02426_),
    .A2(_02429_));
 sg13g2_inv_1 _13854_ (.Y(_03492_),
    .A(_03491_));
 sg13g2_nand2_1 _13855_ (.Y(_03493_),
    .A(_03489_),
    .B(_03492_));
 sg13g2_nand2b_1 _13856_ (.Y(_03494_),
    .B(_03491_),
    .A_N(_03489_));
 sg13g2_a21oi_1 _13857_ (.A1(_02402_),
    .A2(_02405_),
    .Y(_03495_),
    .B1(_02400_));
 sg13g2_nor2_1 _13858_ (.A(_02406_),
    .B(_03495_),
    .Y(_03496_));
 sg13g2_nand2_1 _13859_ (.Y(_03497_),
    .A(_03494_),
    .B(_03496_));
 sg13g2_a21oi_2 _13860_ (.B1(_02261_),
    .Y(_03498_),
    .A2(_02262_),
    .A1(_02258_));
 sg13g2_nand2_1 _13861_ (.Y(_03499_),
    .A(_02433_),
    .B(_02439_));
 sg13g2_o21ai_1 _13862_ (.B1(_03499_),
    .Y(_03500_),
    .A1(_02435_),
    .A2(_02438_));
 sg13g2_or2_1 _13863_ (.X(_03501_),
    .B(_03500_),
    .A(_03498_));
 sg13g2_nand2_1 _13864_ (.Y(_03502_),
    .A(_03498_),
    .B(_03500_));
 sg13g2_a21oi_2 _13865_ (.B1(_02449_),
    .Y(_03503_),
    .A2(_02450_),
    .A1(_02443_));
 sg13g2_nand2_1 _13866_ (.Y(_03504_),
    .A(_03502_),
    .B(_03503_));
 sg13g2_a22oi_1 _13867_ (.Y(_03505_),
    .B1(_03501_),
    .B2(_03504_),
    .A2(_03497_),
    .A1(_03493_));
 sg13g2_nand4_1 _13868_ (.B(_03497_),
    .C(_03501_),
    .A(_03493_),
    .Y(_03506_),
    .D(_03504_));
 sg13g2_nor2b_1 _13869_ (.A(_03505_),
    .B_N(_03506_),
    .Y(_03507_));
 sg13g2_o21ai_1 _13870_ (.B1(_03506_),
    .Y(_03508_),
    .A1(_03488_),
    .A2(_03505_));
 sg13g2_xnor2_1 _13871_ (.Y(_03509_),
    .A(_03487_),
    .B(_03507_));
 sg13g2_o21ai_1 _13872_ (.B1(_02332_),
    .Y(_03510_),
    .A1(_02333_),
    .A2(_02338_));
 sg13g2_o21ai_1 _13873_ (.B1(_02293_),
    .Y(_03511_),
    .A1(_02289_),
    .A2(_02292_));
 sg13g2_nand2b_1 _13874_ (.Y(_03512_),
    .B(_03511_),
    .A_N(_03510_));
 sg13g2_nand2b_1 _13875_ (.Y(_03513_),
    .B(_03510_),
    .A_N(_03511_));
 sg13g2_a21oi_1 _13876_ (.A1(_02344_),
    .A2(_02347_),
    .Y(_03514_),
    .B1(_02345_));
 sg13g2_nand2_1 _13877_ (.Y(_03515_),
    .A(_03513_),
    .B(_03514_));
 sg13g2_nand2_1 _13878_ (.Y(_03516_),
    .A(_03512_),
    .B(_03515_));
 sg13g2_o21ai_1 _13879_ (.B1(_02107_),
    .Y(_03517_),
    .A1(_02082_),
    .A2(_02092_));
 sg13g2_nand2_1 _13880_ (.Y(_03518_),
    .A(_02093_),
    .B(_03517_));
 sg13g2_a21o_1 _13881_ (.A2(_02310_),
    .A1(_02307_),
    .B1(_02306_),
    .X(_03519_));
 sg13g2_o21ai_1 _13882_ (.B1(_03519_),
    .Y(_03520_),
    .A1(_02307_),
    .A2(_02310_));
 sg13g2_or2_1 _13883_ (.X(_03521_),
    .B(_03520_),
    .A(_03518_));
 sg13g2_nand2_1 _13884_ (.Y(_03522_),
    .A(_03518_),
    .B(_03520_));
 sg13g2_o21ai_1 _13885_ (.B1(_02302_),
    .Y(_03523_),
    .A1(_02296_),
    .A2(_02301_));
 sg13g2_nand2_1 _13886_ (.Y(_03524_),
    .A(_03521_),
    .B(_03523_));
 sg13g2_a21oi_1 _13887_ (.A1(_03522_),
    .A2(_03524_),
    .Y(_03525_),
    .B1(_03516_));
 sg13g2_nand3_1 _13888_ (.B(_03522_),
    .C(_03524_),
    .A(_03516_),
    .Y(_03526_));
 sg13g2_nor2b_1 _13889_ (.A(_03525_),
    .B_N(_03526_),
    .Y(_03527_));
 sg13g2_o21ai_1 _13890_ (.B1(_02274_),
    .Y(_03528_),
    .A1(_02276_),
    .A2(_02280_));
 sg13g2_nand2_1 _13891_ (.Y(_03529_),
    .A(_02318_),
    .B(_02327_));
 sg13g2_and4_1 _13892_ (.A(_02281_),
    .B(_02326_),
    .C(_03528_),
    .D(_03529_),
    .X(_03530_));
 sg13g2_a22oi_1 _13893_ (.Y(_03531_),
    .B1(_03529_),
    .B2(_02326_),
    .A2(_03528_),
    .A1(_02281_));
 sg13g2_a21oi_1 _13894_ (.A1(_02267_),
    .A2(_02270_),
    .Y(_03532_),
    .B1(_02266_));
 sg13g2_nor2_1 _13895_ (.A(_02271_),
    .B(_03532_),
    .Y(_03533_));
 sg13g2_nor2_1 _13896_ (.A(_03531_),
    .B(_03533_),
    .Y(_03534_));
 sg13g2_nor2_2 _13897_ (.A(_03530_),
    .B(_03534_),
    .Y(_03535_));
 sg13g2_inv_1 _13898_ (.Y(_03536_),
    .A(_03535_));
 sg13g2_xnor2_1 _13899_ (.Y(_03537_),
    .A(_03527_),
    .B(_03535_));
 sg13g2_nand2_1 _13900_ (.Y(_03538_),
    .A(_03509_),
    .B(_03537_));
 sg13g2_nor2_1 _13901_ (.A(_03509_),
    .B(_03537_),
    .Y(_03539_));
 sg13g2_a21oi_2 _13902_ (.B1(_02364_),
    .Y(_03540_),
    .A2(_02365_),
    .A1(_02359_));
 sg13g2_nand2_1 _13903_ (.Y(_03541_),
    .A(_02227_),
    .B(_02233_));
 sg13g2_nand3_1 _13904_ (.B(_03540_),
    .C(_03541_),
    .A(_02232_),
    .Y(_03542_));
 sg13g2_a21o_1 _13905_ (.A2(_03541_),
    .A1(_02232_),
    .B1(_03540_),
    .X(_03543_));
 sg13g2_a21oi_2 _13906_ (.B1(_02243_),
    .Y(_03544_),
    .A2(_02244_),
    .A1(_02238_));
 sg13g2_nand2_1 _13907_ (.Y(_03545_),
    .A(_03543_),
    .B(_03544_));
 sg13g2_nand2b_1 _13908_ (.Y(_03546_),
    .B(_02224_),
    .A_N(_02218_));
 sg13g2_nand2_1 _13909_ (.Y(_03547_),
    .A(_02203_),
    .B(_02209_));
 sg13g2_and4_1 _13910_ (.A(_02208_),
    .B(_02223_),
    .C(_03546_),
    .D(_03547_),
    .X(_03548_));
 sg13g2_a22oi_1 _13911_ (.Y(_03549_),
    .B1(_03547_),
    .B2(_02208_),
    .A2(_03546_),
    .A1(_02223_));
 sg13g2_inv_1 _13912_ (.Y(_03550_),
    .A(_03549_));
 sg13g2_a21o_1 _13913_ (.A2(_02200_),
    .A1(_02198_),
    .B1(_02195_),
    .X(_03551_));
 sg13g2_o21ai_1 _13914_ (.B1(_03551_),
    .Y(_03552_),
    .A1(_02198_),
    .A2(_02200_));
 sg13g2_o21ai_1 _13915_ (.B1(_03550_),
    .Y(_03553_),
    .A1(_03548_),
    .A2(_03552_));
 sg13g2_a21oi_2 _13916_ (.B1(_03553_),
    .Y(_03554_),
    .A2(_03545_),
    .A1(_03542_));
 sg13g2_nand3_1 _13917_ (.B(_03545_),
    .C(_03553_),
    .A(_03542_),
    .Y(_03555_));
 sg13g2_nor2b_1 _13918_ (.A(_03554_),
    .B_N(_03555_),
    .Y(_03556_));
 sg13g2_a21oi_1 _13919_ (.A1(_03433_),
    .A2(_03437_),
    .Y(_03557_),
    .B1(_03434_));
 sg13g2_xnor2_1 _13920_ (.Y(_03558_),
    .A(_03556_),
    .B(_03557_));
 sg13g2_a21oi_2 _13921_ (.B1(_03539_),
    .Y(_03559_),
    .A2(_03558_),
    .A1(_03538_));
 sg13g2_and2_1 _13922_ (.A(_03480_),
    .B(_03559_),
    .X(_03560_));
 sg13g2_nor2_1 _13923_ (.A(_03480_),
    .B(_03559_),
    .Y(_03561_));
 sg13g2_nor2b_1 _13924_ (.A(_03400_),
    .B_N(_03404_),
    .Y(_03562_));
 sg13g2_nor2_2 _13925_ (.A(_03403_),
    .B(_03562_),
    .Y(_03563_));
 sg13g2_nand2_1 _13926_ (.Y(_03564_),
    .A(_03442_),
    .B(_03446_));
 sg13g2_nand2_2 _13927_ (.Y(_03565_),
    .A(_03447_),
    .B(_03564_));
 sg13g2_nor2_1 _13928_ (.A(_03426_),
    .B(_03565_),
    .Y(_03566_));
 sg13g2_xnor2_1 _13929_ (.Y(_03567_),
    .A(_03425_),
    .B(_03565_));
 sg13g2_xnor2_1 _13930_ (.Y(_03568_),
    .A(_03397_),
    .B(_03567_));
 sg13g2_nor2_1 _13931_ (.A(_03563_),
    .B(_03568_),
    .Y(_03569_));
 sg13g2_and2_1 _13932_ (.A(_03563_),
    .B(_03568_),
    .X(_03570_));
 sg13g2_a21oi_2 _13933_ (.B1(_03416_),
    .Y(_03571_),
    .A2(_03414_),
    .A1(_03410_));
 sg13g2_nor2_1 _13934_ (.A(_03569_),
    .B(_03571_),
    .Y(_03572_));
 sg13g2_nor2_1 _13935_ (.A(_03570_),
    .B(_03572_),
    .Y(_03573_));
 sg13g2_nor2_1 _13936_ (.A(_03560_),
    .B(_03573_),
    .Y(_03574_));
 sg13g2_nor2_1 _13937_ (.A(_03561_),
    .B(_03574_),
    .Y(_03575_));
 sg13g2_nor2_1 _13938_ (.A(_03569_),
    .B(_03570_),
    .Y(_03576_));
 sg13g2_xnor2_1 _13939_ (.Y(_03577_),
    .A(_03571_),
    .B(_03576_));
 sg13g2_nand2_1 _13940_ (.Y(_03578_),
    .A(_03455_),
    .B(_03456_));
 sg13g2_xor2_1 _13941_ (.B(_03578_),
    .A(_03478_),
    .X(_03579_));
 sg13g2_inv_1 _13942_ (.Y(_03580_),
    .A(_03579_));
 sg13g2_nand2_1 _13943_ (.Y(_03581_),
    .A(_03521_),
    .B(_03522_));
 sg13g2_xor2_1 _13944_ (.B(_03581_),
    .A(_03523_),
    .X(_03582_));
 sg13g2_xor2_1 _13945_ (.B(_03458_),
    .A(_02065_),
    .X(_03583_));
 sg13g2_xnor2_1 _13946_ (.Y(_03584_),
    .A(_02139_),
    .B(_03583_));
 sg13g2_nand2_1 _13947_ (.Y(_03585_),
    .A(_03582_),
    .B(_03584_));
 sg13g2_or2_1 _13948_ (.X(_03586_),
    .B(_03584_),
    .A(_03582_));
 sg13g2_and2_1 _13949_ (.A(_03512_),
    .B(_03513_),
    .X(_03587_));
 sg13g2_xnor2_1 _13950_ (.Y(_03588_),
    .A(_03514_),
    .B(_03587_));
 sg13g2_nand2_1 _13951_ (.Y(_03589_),
    .A(_03585_),
    .B(_03588_));
 sg13g2_nand2_1 _13952_ (.Y(_03590_),
    .A(_03501_),
    .B(_03502_));
 sg13g2_xor2_1 _13953_ (.B(_03590_),
    .A(_03503_),
    .X(_03591_));
 sg13g2_nor2_1 _13954_ (.A(_03530_),
    .B(_03531_),
    .Y(_03592_));
 sg13g2_xnor2_1 _13955_ (.Y(_03593_),
    .A(_03533_),
    .B(_03592_));
 sg13g2_nand2b_1 _13956_ (.Y(_03594_),
    .B(_03593_),
    .A_N(_03591_));
 sg13g2_nand2b_1 _13957_ (.Y(_03595_),
    .B(_03591_),
    .A_N(_03593_));
 sg13g2_nand2_1 _13958_ (.Y(_03596_),
    .A(_03493_),
    .B(_03494_));
 sg13g2_xor2_1 _13959_ (.B(_03596_),
    .A(_03496_),
    .X(_03597_));
 sg13g2_nand2_1 _13960_ (.Y(_03598_),
    .A(_03594_),
    .B(_03597_));
 sg13g2_nand2_1 _13961_ (.Y(_03599_),
    .A(_03595_),
    .B(_03598_));
 sg13g2_a21oi_1 _13962_ (.A1(_03586_),
    .A2(_03589_),
    .Y(_03600_),
    .B1(_03599_));
 sg13g2_nand3_1 _13963_ (.B(_03589_),
    .C(_03599_),
    .A(_03586_),
    .Y(_03601_));
 sg13g2_nor2b_1 _13964_ (.A(_03600_),
    .B_N(_03601_),
    .Y(_03602_));
 sg13g2_xor2_1 _13965_ (.B(_03482_),
    .A(_03481_),
    .X(_03603_));
 sg13g2_xnor2_1 _13966_ (.Y(_03604_),
    .A(_03486_),
    .B(_03603_));
 sg13g2_nand2_1 _13967_ (.Y(_03605_),
    .A(_03542_),
    .B(_03543_));
 sg13g2_xnor2_1 _13968_ (.Y(_03606_),
    .A(_03544_),
    .B(_03605_));
 sg13g2_nand2_1 _13969_ (.Y(_03607_),
    .A(_03604_),
    .B(_03606_));
 sg13g2_nor2_1 _13970_ (.A(_03604_),
    .B(_03606_),
    .Y(_03608_));
 sg13g2_nor2_1 _13971_ (.A(_03548_),
    .B(_03549_),
    .Y(_03609_));
 sg13g2_xnor2_1 _13972_ (.Y(_03610_),
    .A(_03552_),
    .B(_03609_));
 sg13g2_a21oi_2 _13973_ (.B1(_03608_),
    .Y(_03611_),
    .A2(_03610_),
    .A1(_03607_));
 sg13g2_xnor2_1 _13974_ (.Y(_03612_),
    .A(_03602_),
    .B(_03611_));
 sg13g2_a21oi_2 _13975_ (.B1(_02103_),
    .Y(_03613_),
    .A2(_02105_),
    .A1(_02097_));
 sg13g2_inv_1 _13976_ (.Y(_03614_),
    .A(_03613_));
 sg13g2_nand2_1 _13977_ (.Y(_03615_),
    .A(_03594_),
    .B(_03595_));
 sg13g2_xor2_1 _13978_ (.B(_03615_),
    .A(_03597_),
    .X(_03616_));
 sg13g2_xor2_1 _13979_ (.B(_03606_),
    .A(_03604_),
    .X(_03617_));
 sg13g2_xnor2_1 _13980_ (.Y(_03618_),
    .A(_03610_),
    .B(_03617_));
 sg13g2_nand2_1 _13981_ (.Y(_03619_),
    .A(_03616_),
    .B(_03618_));
 sg13g2_xor2_1 _13982_ (.B(_03618_),
    .A(_03616_),
    .X(_03620_));
 sg13g2_and2_1 _13983_ (.A(_03439_),
    .B(_03440_),
    .X(_03621_));
 sg13g2_xnor2_1 _13984_ (.Y(_03622_),
    .A(_03449_),
    .B(_03621_));
 sg13g2_xnor2_1 _13985_ (.Y(_03623_),
    .A(_03620_),
    .B(_03622_));
 sg13g2_xor2_1 _13986_ (.B(_03463_),
    .A(_03462_),
    .X(_03624_));
 sg13g2_xnor2_1 _13987_ (.Y(_03625_),
    .A(_03465_),
    .B(_03624_));
 sg13g2_xnor2_1 _13988_ (.Y(_03626_),
    .A(_03362_),
    .B(_03363_));
 sg13g2_xnor2_1 _13989_ (.Y(_03627_),
    .A(_03364_),
    .B(_03626_));
 sg13g2_nand2_1 _13990_ (.Y(_03628_),
    .A(_03625_),
    .B(_03627_));
 sg13g2_nor2_1 _13991_ (.A(_03625_),
    .B(_03627_),
    .Y(_03629_));
 sg13g2_xor2_1 _13992_ (.B(_03627_),
    .A(_03625_),
    .X(_03630_));
 sg13g2_nand2b_1 _13993_ (.Y(_03631_),
    .B(_03470_),
    .A_N(_03469_));
 sg13g2_xnor2_1 _13994_ (.Y(_03632_),
    .A(_03471_),
    .B(_03631_));
 sg13g2_xnor2_1 _13995_ (.Y(_03633_),
    .A(_03630_),
    .B(_03632_));
 sg13g2_nand2b_1 _13996_ (.Y(_03634_),
    .B(_02146_),
    .A_N(_03385_));
 sg13g2_o21ai_1 _13997_ (.B1(_03634_),
    .Y(_03635_),
    .A1(_03386_),
    .A2(_03388_));
 sg13g2_nor2_1 _13998_ (.A(_03376_),
    .B(_03377_),
    .Y(_03636_));
 sg13g2_xnor2_1 _13999_ (.Y(_03637_),
    .A(_02255_),
    .B(_03636_));
 sg13g2_xor2_1 _14000_ (.B(_03637_),
    .A(_03635_),
    .X(_03638_));
 sg13g2_nand2_1 _14001_ (.Y(_03639_),
    .A(_03368_),
    .B(_03369_));
 sg13g2_xor2_1 _14002_ (.B(_03639_),
    .A(_03371_),
    .X(_03640_));
 sg13g2_xnor2_1 _14003_ (.Y(_03641_),
    .A(_03638_),
    .B(_03640_));
 sg13g2_nor2_1 _14004_ (.A(_03633_),
    .B(_03641_),
    .Y(_03642_));
 sg13g2_nand2_1 _14005_ (.Y(_03643_),
    .A(_03633_),
    .B(_03641_));
 sg13g2_xnor2_1 _14006_ (.Y(_03644_),
    .A(_03633_),
    .B(_03641_));
 sg13g2_nand2_1 _14007_ (.Y(_03645_),
    .A(_03585_),
    .B(_03586_));
 sg13g2_xor2_1 _14008_ (.B(_03645_),
    .A(_03588_),
    .X(_03646_));
 sg13g2_xnor2_1 _14009_ (.Y(_03647_),
    .A(_03644_),
    .B(_03646_));
 sg13g2_and2_1 _14010_ (.A(_03623_),
    .B(_03647_),
    .X(_03648_));
 sg13g2_or2_1 _14011_ (.X(_03649_),
    .B(_03647_),
    .A(_03623_));
 sg13g2_xor2_1 _14012_ (.B(_03647_),
    .A(_03623_),
    .X(_03650_));
 sg13g2_and2_1 _14013_ (.A(_03407_),
    .B(_03408_),
    .X(_03651_));
 sg13g2_xnor2_1 _14014_ (.Y(_03652_),
    .A(_03418_),
    .B(_03651_));
 sg13g2_xnor2_1 _14015_ (.Y(_03653_),
    .A(_03650_),
    .B(_03652_));
 sg13g2_nand2b_2 _14016_ (.Y(_03654_),
    .B(_03614_),
    .A_N(_03653_));
 sg13g2_o21ai_1 _14017_ (.B1(_03649_),
    .Y(_03655_),
    .A1(_03648_),
    .A2(_03652_));
 sg13g2_o21ai_1 _14018_ (.B1(_03655_),
    .Y(_03656_),
    .A1(_03613_),
    .A2(_03653_));
 sg13g2_and4_1 _14019_ (.A(_03614_),
    .B(_03648_),
    .C(_03649_),
    .D(_03652_),
    .X(_03657_));
 sg13g2_inv_1 _14020_ (.Y(_03658_),
    .A(_03657_));
 sg13g2_a21oi_1 _14021_ (.A1(_03643_),
    .A2(_03646_),
    .Y(_03659_),
    .B1(_03642_));
 sg13g2_nand3_1 _14022_ (.B(_03658_),
    .C(_03659_),
    .A(_03656_),
    .Y(_03660_));
 sg13g2_a21o_1 _14023_ (.A2(_03658_),
    .A1(_03656_),
    .B1(_03659_),
    .X(_03661_));
 sg13g2_a21o_1 _14024_ (.A2(_03637_),
    .A1(_03635_),
    .B1(_03640_),
    .X(_03662_));
 sg13g2_o21ai_1 _14025_ (.B1(_03662_),
    .Y(_03663_),
    .A1(_03635_),
    .A2(_03637_));
 sg13g2_o21ai_1 _14026_ (.B1(_03622_),
    .Y(_03664_),
    .A1(_03616_),
    .A2(_03618_));
 sg13g2_nand2_1 _14027_ (.Y(_03665_),
    .A(_03619_),
    .B(_03664_));
 sg13g2_nand2_1 _14028_ (.Y(_03666_),
    .A(_03663_),
    .B(_03665_));
 sg13g2_inv_1 _14029_ (.Y(_03667_),
    .A(_03666_));
 sg13g2_nor2_1 _14030_ (.A(_03663_),
    .B(_03665_),
    .Y(_03668_));
 sg13g2_nor2_1 _14031_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sg13g2_a21oi_1 _14032_ (.A1(_03628_),
    .A2(_03632_),
    .Y(_03670_),
    .B1(_03629_));
 sg13g2_xnor2_1 _14033_ (.Y(_03671_),
    .A(_03669_),
    .B(_03670_));
 sg13g2_inv_1 _14034_ (.Y(_03672_),
    .A(_03671_));
 sg13g2_a21oi_2 _14035_ (.B1(_03672_),
    .Y(_03673_),
    .A2(_03661_),
    .A1(_03660_));
 sg13g2_and3_1 _14036_ (.X(_03674_),
    .A(_03660_),
    .B(_03661_),
    .C(_03672_));
 sg13g2_nand3_1 _14037_ (.B(_03661_),
    .C(_03672_),
    .A(_03660_),
    .Y(_03675_));
 sg13g2_or3_1 _14038_ (.A(_03612_),
    .B(_03673_),
    .C(_03674_),
    .X(_03676_));
 sg13g2_o21ai_1 _14039_ (.B1(_03612_),
    .Y(_03677_),
    .A1(_03673_),
    .A2(_03674_));
 sg13g2_and3_1 _14040_ (.X(_03678_),
    .A(_03580_),
    .B(_03676_),
    .C(_03677_));
 sg13g2_a21oi_1 _14041_ (.A1(_03676_),
    .A2(_03677_),
    .Y(_03679_),
    .B1(_03580_));
 sg13g2_xor2_1 _14042_ (.B(_03537_),
    .A(_03509_),
    .X(_03680_));
 sg13g2_xnor2_1 _14043_ (.Y(_03681_),
    .A(_03558_),
    .B(_03680_));
 sg13g2_or3_1 _14044_ (.A(_03678_),
    .B(_03679_),
    .C(_03681_),
    .X(_03682_));
 sg13g2_o21ai_1 _14045_ (.B1(_03681_),
    .Y(_03683_),
    .A1(_03678_),
    .A2(_03679_));
 sg13g2_nand2_1 _14046_ (.Y(_03684_),
    .A(_03682_),
    .B(_03683_));
 sg13g2_and3_1 _14047_ (.X(_03685_),
    .A(_03577_),
    .B(_03682_),
    .C(_03683_));
 sg13g2_nor2b_1 _14048_ (.A(_03679_),
    .B_N(_03681_),
    .Y(_03686_));
 sg13g2_nor2_1 _14049_ (.A(_03678_),
    .B(_03686_),
    .Y(_03687_));
 sg13g2_nor2_1 _14050_ (.A(_03685_),
    .B(_03687_),
    .Y(_03688_));
 sg13g2_a21oi_1 _14051_ (.A1(_03612_),
    .A2(_03675_),
    .Y(_03689_),
    .B1(_03673_));
 sg13g2_a221oi_1 _14052_ (.B2(_03687_),
    .C1(_03673_),
    .B1(_03685_),
    .A1(_03612_),
    .Y(_03690_),
    .A2(_03675_));
 sg13g2_o21ai_1 _14053_ (.B1(_03575_),
    .Y(_03691_),
    .A1(_03688_),
    .A2(_03690_));
 sg13g2_nor3_1 _14054_ (.A(_03575_),
    .B(_03688_),
    .C(_03690_),
    .Y(_03692_));
 sg13g2_inv_1 _14055_ (.Y(_03693_),
    .A(_03692_));
 sg13g2_nand2_1 _14056_ (.Y(_03694_),
    .A(_03658_),
    .B(_03659_));
 sg13g2_nor2_1 _14057_ (.A(_03667_),
    .B(_03670_),
    .Y(_03695_));
 sg13g2_or2_1 _14058_ (.X(_03696_),
    .B(_03695_),
    .A(_03668_));
 sg13g2_a21o_1 _14059_ (.A2(_03694_),
    .A1(_03656_),
    .B1(_03696_),
    .X(_03697_));
 sg13g2_inv_1 _14060_ (.Y(_03698_),
    .A(_03697_));
 sg13g2_and3_1 _14061_ (.X(_03699_),
    .A(_03656_),
    .B(_03694_),
    .C(_03696_));
 sg13g2_o21ai_1 _14062_ (.B1(_03601_),
    .Y(_03700_),
    .A1(_03600_),
    .A2(_03611_));
 sg13g2_a21oi_2 _14063_ (.B1(_03699_),
    .Y(_03701_),
    .A2(_03700_),
    .A1(_03697_));
 sg13g2_inv_1 _14064_ (.Y(_03702_),
    .A(_03701_));
 sg13g2_a21oi_2 _14065_ (.B1(_03692_),
    .Y(_03703_),
    .A2(_03702_),
    .A1(_03691_));
 sg13g2_inv_1 _14066_ (.Y(_03704_),
    .A(_03703_));
 sg13g2_xnor2_1 _14067_ (.Y(_03705_),
    .A(_03685_),
    .B(_03687_));
 sg13g2_xor2_1 _14068_ (.B(_03705_),
    .A(_03689_),
    .X(_03706_));
 sg13g2_nor2_1 _14069_ (.A(_03560_),
    .B(_03561_),
    .Y(_03707_));
 sg13g2_xnor2_1 _14070_ (.Y(_03708_),
    .A(_03573_),
    .B(_03707_));
 sg13g2_nand2_1 _14071_ (.Y(_03709_),
    .A(_03706_),
    .B(_03708_));
 sg13g2_nor2_1 _14072_ (.A(_03706_),
    .B(_03708_),
    .Y(_03710_));
 sg13g2_nor2_1 _14073_ (.A(_03698_),
    .B(_03699_),
    .Y(_03711_));
 sg13g2_xnor2_1 _14074_ (.Y(_03712_),
    .A(_03700_),
    .B(_03711_));
 sg13g2_a21oi_1 _14075_ (.A1(_03709_),
    .A2(_03712_),
    .Y(_03713_),
    .B1(_03710_));
 sg13g2_nand3b_1 _14076_ (.B(_03706_),
    .C(_03708_),
    .Y(_03714_),
    .A_N(_03712_));
 sg13g2_nand2_1 _14077_ (.Y(_03715_),
    .A(_03710_),
    .B(_03712_));
 sg13g2_a22oi_1 _14078_ (.Y(_03716_),
    .B1(_03713_),
    .B2(_03714_),
    .A2(_03712_),
    .A1(_03710_));
 sg13g2_nor2_1 _14079_ (.A(_03397_),
    .B(_03566_),
    .Y(_03717_));
 sg13g2_a21o_1 _14080_ (.A2(_03565_),
    .A1(_03426_),
    .B1(_03717_),
    .X(_03718_));
 sg13g2_o21ai_1 _14081_ (.B1(_03526_),
    .Y(_03719_),
    .A1(_03525_),
    .A2(_03536_));
 sg13g2_or2_1 _14082_ (.X(_03720_),
    .B(_03719_),
    .A(_03508_));
 sg13g2_nand2_1 _14083_ (.Y(_03721_),
    .A(_03508_),
    .B(_03719_));
 sg13g2_nand2_1 _14084_ (.Y(_03722_),
    .A(_03720_),
    .B(_03721_));
 sg13g2_o21ai_1 _14085_ (.B1(_03555_),
    .Y(_03723_),
    .A1(_03554_),
    .A2(_03557_));
 sg13g2_xnor2_1 _14086_ (.Y(_03724_),
    .A(_03722_),
    .B(_03723_));
 sg13g2_nand2_1 _14087_ (.Y(_03725_),
    .A(_03389_),
    .B(_03451_));
 sg13g2_and2_1 _14088_ (.A(_03452_),
    .B(_03725_),
    .X(_03726_));
 sg13g2_a21oi_1 _14089_ (.A1(_03366_),
    .A2(_03381_),
    .Y(_03727_),
    .B1(_03382_));
 sg13g2_nor2_1 _14090_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sg13g2_and2_1 _14091_ (.A(_03726_),
    .B(_03727_),
    .X(_03729_));
 sg13g2_nor2_1 _14092_ (.A(_03476_),
    .B(_03729_),
    .Y(_03730_));
 sg13g2_nor2_1 _14093_ (.A(_03728_),
    .B(_03730_),
    .Y(_03731_));
 sg13g2_inv_1 _14094_ (.Y(_03732_),
    .A(_03731_));
 sg13g2_nand2b_1 _14095_ (.Y(_03733_),
    .B(_03728_),
    .A_N(_03476_));
 sg13g2_a22oi_1 _14096_ (.Y(_03734_),
    .B1(_03732_),
    .B2(_03733_),
    .A2(_03729_),
    .A1(_03476_));
 sg13g2_xor2_1 _14097_ (.B(_03734_),
    .A(_03724_),
    .X(_03735_));
 sg13g2_xnor2_1 _14098_ (.Y(_03736_),
    .A(_03718_),
    .B(_03735_));
 sg13g2_inv_1 _14099_ (.Y(_03737_),
    .A(_03736_));
 sg13g2_a21oi_1 _14100_ (.A1(_03715_),
    .A2(_03737_),
    .Y(_03738_),
    .B1(_03713_));
 sg13g2_a21o_1 _14101_ (.A2(_03734_),
    .A1(_03724_),
    .B1(_03718_),
    .X(_03739_));
 sg13g2_o21ai_1 _14102_ (.B1(_03739_),
    .Y(_03740_),
    .A1(_03724_),
    .A2(_03734_));
 sg13g2_nand2b_1 _14103_ (.Y(_03741_),
    .B(_03737_),
    .A_N(_03714_));
 sg13g2_nand2_1 _14104_ (.Y(_03742_),
    .A(_03740_),
    .B(_03741_));
 sg13g2_nor2b_1 _14105_ (.A(_03738_),
    .B_N(_03742_),
    .Y(_03743_));
 sg13g2_o21ai_1 _14106_ (.B1(_03703_),
    .Y(_03744_),
    .A1(_03691_),
    .A2(_03702_));
 sg13g2_o21ai_1 _14107_ (.B1(_03744_),
    .Y(_03745_),
    .A1(_03693_),
    .A2(_03701_));
 sg13g2_nand2_1 _14108_ (.Y(_03746_),
    .A(_03738_),
    .B(_03740_));
 sg13g2_or2_1 _14109_ (.X(_03747_),
    .B(_03741_),
    .A(_03740_));
 sg13g2_nand3b_1 _14110_ (.B(_03742_),
    .C(_03747_),
    .Y(_03748_),
    .A_N(_03738_));
 sg13g2_a21o_1 _14111_ (.A2(_03748_),
    .A1(_03746_),
    .B1(_03745_),
    .X(_03749_));
 sg13g2_nand3_1 _14112_ (.B(_03746_),
    .C(_03748_),
    .A(_03745_),
    .Y(_03750_));
 sg13g2_a21oi_1 _14113_ (.A1(_03749_),
    .A2(_03750_),
    .Y(_03751_),
    .B1(_03732_));
 sg13g2_and3_1 _14114_ (.X(_03752_),
    .A(_03732_),
    .B(_03749_),
    .C(_03750_));
 sg13g2_nand2_1 _14115_ (.Y(_03753_),
    .A(_03720_),
    .B(_03723_));
 sg13g2_and2_1 _14116_ (.A(_03721_),
    .B(_03753_),
    .X(_03754_));
 sg13g2_nor3_2 _14117_ (.A(_03751_),
    .B(_03752_),
    .C(_03754_),
    .Y(_03755_));
 sg13g2_inv_1 _14118_ (.Y(_03756_),
    .A(_03755_));
 sg13g2_nand2_1 _14119_ (.Y(_03757_),
    .A(_03731_),
    .B(_03750_));
 sg13g2_and2_1 _14120_ (.A(_03749_),
    .B(_03757_),
    .X(_03758_));
 sg13g2_nor2_1 _14121_ (.A(_03755_),
    .B(_03758_),
    .Y(_03759_));
 sg13g2_xnor2_1 _14122_ (.Y(_03760_),
    .A(_03755_),
    .B(_03758_));
 sg13g2_xnor2_1 _14123_ (.Y(_03761_),
    .A(_03743_),
    .B(_03760_));
 sg13g2_nor2b_1 _14124_ (.A(_03759_),
    .B_N(_03743_),
    .Y(_03762_));
 sg13g2_a221oi_1 _14125_ (.B2(_03704_),
    .C1(_03762_),
    .B1(_03761_),
    .A1(_03755_),
    .Y(_03763_),
    .A2(_03758_));
 sg13g2_nor2_1 _14126_ (.A(_03361_),
    .B(_03763_),
    .Y(_03764_));
 sg13g2_or2_1 _14127_ (.X(_03765_),
    .B(_03763_),
    .A(_03361_));
 sg13g2_xnor2_1 _14128_ (.Y(_03766_),
    .A(_03703_),
    .B(_03761_));
 sg13g2_xnor2_1 _14129_ (.Y(_03767_),
    .A(_03704_),
    .B(_03761_));
 sg13g2_a21oi_2 _14130_ (.B1(_03301_),
    .Y(_03768_),
    .A2(_03358_),
    .A1(_03357_));
 sg13g2_nor2_1 _14131_ (.A(_03359_),
    .B(_03768_),
    .Y(_03769_));
 sg13g2_nand3_1 _14132_ (.B(_03328_),
    .C(_03338_),
    .A(_03327_),
    .Y(_03770_));
 sg13g2_nor2b_2 _14133_ (.A(_03339_),
    .B_N(_03770_),
    .Y(_03771_));
 sg13g2_xor2_1 _14134_ (.B(_03195_),
    .A(_03193_),
    .X(_03772_));
 sg13g2_nand2_2 _14135_ (.Y(_03773_),
    .A(_03613_),
    .B(_03653_));
 sg13g2_nand2_2 _14136_ (.Y(_03774_),
    .A(_03654_),
    .B(_03773_));
 sg13g2_nor2_1 _14137_ (.A(_03772_),
    .B(_03774_),
    .Y(_03775_));
 sg13g2_nand2_1 _14138_ (.Y(_03776_),
    .A(_03772_),
    .B(_03774_));
 sg13g2_nand2_1 _14139_ (.Y(_03777_),
    .A(_02985_),
    .B(_02989_));
 sg13g2_xor2_1 _14140_ (.B(_03777_),
    .A(_02987_),
    .X(_03778_));
 sg13g2_nand2b_1 _14141_ (.Y(_03779_),
    .B(_03778_),
    .A_N(_02466_));
 sg13g2_a21o_1 _14142_ (.A2(_03779_),
    .A1(_03776_),
    .B1(_03775_),
    .X(_03780_));
 sg13g2_xnor2_1 _14143_ (.Y(_03781_),
    .A(_03577_),
    .B(_03684_));
 sg13g2_xor2_1 _14144_ (.B(_03279_),
    .A(_03265_),
    .X(_03782_));
 sg13g2_inv_1 _14145_ (.Y(_03783_),
    .A(_03782_));
 sg13g2_o21ai_1 _14146_ (.B1(_03782_),
    .Y(_03784_),
    .A1(_03780_),
    .A2(_03781_));
 sg13g2_inv_1 _14147_ (.Y(_03785_),
    .A(_03784_));
 sg13g2_a21oi_1 _14148_ (.A1(_03780_),
    .A2(_03781_),
    .Y(_03786_),
    .B1(_03785_));
 sg13g2_nor2_1 _14149_ (.A(_03771_),
    .B(_03786_),
    .Y(_03787_));
 sg13g2_nand2_1 _14150_ (.Y(_03788_),
    .A(_03771_),
    .B(_03786_));
 sg13g2_xnor2_1 _14151_ (.Y(_03789_),
    .A(_03716_),
    .B(_03736_));
 sg13g2_o21ai_1 _14152_ (.B1(_03788_),
    .Y(_03790_),
    .A1(_03787_),
    .A2(_03789_));
 sg13g2_xnor2_1 _14153_ (.Y(_03791_),
    .A(_03310_),
    .B(_03351_));
 sg13g2_or2_1 _14154_ (.X(_03792_),
    .B(_03791_),
    .A(_03790_));
 sg13g2_and2_1 _14155_ (.A(_03790_),
    .B(_03791_),
    .X(_03793_));
 sg13g2_o21ai_1 _14156_ (.B1(_03754_),
    .Y(_03794_),
    .A1(_03751_),
    .A2(_03752_));
 sg13g2_nand2b_1 _14157_ (.Y(_03795_),
    .B(_03794_),
    .A_N(_03755_));
 sg13g2_a21oi_1 _14158_ (.A1(_03792_),
    .A2(_03795_),
    .Y(_03796_),
    .B1(_03793_));
 sg13g2_o21ai_1 _14159_ (.B1(_03796_),
    .Y(_03797_),
    .A1(_03359_),
    .A2(_03768_));
 sg13g2_and2_1 _14160_ (.A(_03361_),
    .B(_03763_),
    .X(_03798_));
 sg13g2_nor3_1 _14161_ (.A(_03359_),
    .B(_03768_),
    .C(_03796_),
    .Y(_03799_));
 sg13g2_a21o_1 _14162_ (.A2(_03797_),
    .A1(_03767_),
    .B1(_03799_),
    .X(_03800_));
 sg13g2_a221oi_1 _14163_ (.B2(_03797_),
    .C1(_03799_),
    .B1(_03767_),
    .A1(_03361_),
    .Y(_03801_),
    .A2(_03763_));
 sg13g2_nor2_2 _14164_ (.A(net2175),
    .B(net2173),
    .Y(_03802_));
 sg13g2_nor3_2 _14165_ (.A(net2176),
    .B(_03778_),
    .C(net2174),
    .Y(_03803_));
 sg13g2_a221oi_1 _14166_ (.B2(_03800_),
    .C1(_03798_),
    .B1(_03765_),
    .A1(_02464_),
    .Y(_03804_),
    .A2(_02465_));
 sg13g2_nor2_1 _14167_ (.A(_03803_),
    .B(_03804_),
    .Y(_03805_));
 sg13g2_nand2b_1 _14168_ (.Y(_03806_),
    .B(net2609),
    .A_N(net2264));
 sg13g2_o21ai_1 _14169_ (.B1(_03806_),
    .Y(_03807_),
    .A1(net2557),
    .A2(net2535));
 sg13g2_a21oi_2 _14170_ (.B1(_03807_),
    .Y(_03808_),
    .A2(net2265),
    .A1(_05231_));
 sg13g2_nor2_1 _14171_ (.A(net2398),
    .B(net2410),
    .Y(_03809_));
 sg13g2_xor2_1 _14172_ (.B(net2658),
    .A(net2553),
    .X(_03810_));
 sg13g2_xnor2_1 _14173_ (.Y(_03811_),
    .A(_03809_),
    .B(_03810_));
 sg13g2_nor2_1 _14174_ (.A(_03808_),
    .B(_03811_),
    .Y(_03812_));
 sg13g2_nand2_1 _14175_ (.Y(_03813_),
    .A(_03808_),
    .B(_03811_));
 sg13g2_xnor2_1 _14176_ (.Y(_03814_),
    .A(net2686),
    .B(net2763));
 sg13g2_nor2_1 _14177_ (.A(net2705),
    .B(_03814_),
    .Y(_03815_));
 sg13g2_o21ai_1 _14178_ (.B1(_03813_),
    .Y(_03816_),
    .A1(_03812_),
    .A2(_03815_));
 sg13g2_inv_1 _14179_ (.Y(_03817_),
    .A(_03816_));
 sg13g2_nand2b_2 _14180_ (.Y(_03818_),
    .B(net2531),
    .A_N(net2233));
 sg13g2_nor3_2 _14181_ (.A(net2302),
    .B(net2278),
    .C(_03818_),
    .Y(_03819_));
 sg13g2_nor2b_1 _14182_ (.A(net2814),
    .B_N(net2341),
    .Y(_03820_));
 sg13g2_nor2b_1 _14183_ (.A(net2200),
    .B_N(net2425),
    .Y(_03821_));
 sg13g2_xnor2_1 _14184_ (.Y(_03822_),
    .A(_03820_),
    .B(_03821_));
 sg13g2_nand2b_1 _14185_ (.Y(_03823_),
    .B(_03822_),
    .A_N(_03819_));
 sg13g2_nor2b_1 _14186_ (.A(_03822_),
    .B_N(_03819_),
    .Y(_03824_));
 sg13g2_nor2_1 _14187_ (.A(net2720),
    .B(net2759),
    .Y(_03825_));
 sg13g2_xnor2_1 _14188_ (.Y(_03826_),
    .A(net2789),
    .B(net2497));
 sg13g2_xnor2_1 _14189_ (.Y(_03827_),
    .A(_03825_),
    .B(_03826_));
 sg13g2_a21oi_2 _14190_ (.B1(_03824_),
    .Y(_03828_),
    .A2(_03827_),
    .A1(_03823_));
 sg13g2_nand2_1 _14191_ (.Y(_03829_),
    .A(_03817_),
    .B(_03828_));
 sg13g2_nor2_1 _14192_ (.A(_03817_),
    .B(_03828_),
    .Y(_03830_));
 sg13g2_o21ai_1 _14193_ (.B1(_05297_),
    .Y(_03831_),
    .A1(net2260),
    .A2(net2728));
 sg13g2_nand2_1 _14194_ (.Y(_03832_),
    .A(net2587),
    .B(_06023_));
 sg13g2_nor2_1 _14195_ (.A(net2754),
    .B(net2734),
    .Y(_03833_));
 sg13g2_xnor2_1 _14196_ (.Y(_03834_),
    .A(_03832_),
    .B(_03833_));
 sg13g2_nor2_1 _14197_ (.A(_03831_),
    .B(_03834_),
    .Y(_03835_));
 sg13g2_a21oi_2 _14198_ (.B1(net2265),
    .Y(_03836_),
    .A2(net2738),
    .A1(_05495_));
 sg13g2_a21oi_1 _14199_ (.A1(_03831_),
    .A2(_03834_),
    .Y(_03837_),
    .B1(_03836_));
 sg13g2_nor2_2 _14200_ (.A(_03835_),
    .B(_03837_),
    .Y(_03838_));
 sg13g2_a21oi_1 _14201_ (.A1(_03829_),
    .A2(_03838_),
    .Y(_03839_),
    .B1(_03830_));
 sg13g2_inv_1 _14202_ (.Y(_03840_),
    .A(_03839_));
 sg13g2_nor2_1 _14203_ (.A(net2483),
    .B(\net.in[237] ),
    .Y(_03841_));
 sg13g2_nand2_1 _14204_ (.Y(_03842_),
    .A(net2184),
    .B(_05924_));
 sg13g2_nor2_1 _14205_ (.A(_09158_),
    .B(_03842_),
    .Y(_03843_));
 sg13g2_xnor2_1 _14206_ (.Y(_03844_),
    .A(net2762),
    .B(net2690));
 sg13g2_a21oi_1 _14207_ (.A1(_09158_),
    .A2(_03842_),
    .Y(_03845_),
    .B1(_03844_));
 sg13g2_or2_2 _14208_ (.X(_03846_),
    .B(_03845_),
    .A(_03843_));
 sg13g2_nor2_1 _14209_ (.A(net2256),
    .B(net2668),
    .Y(_03847_));
 sg13g2_nand2b_1 _14210_ (.Y(_03848_),
    .B(net2505),
    .A_N(net2716));
 sg13g2_xnor2_1 _14211_ (.Y(_03849_),
    .A(_03847_),
    .B(_03848_));
 sg13g2_and2_1 _14212_ (.A(net2567),
    .B(net2773),
    .X(_03850_));
 sg13g2_nor2_2 _14213_ (.A(net2773),
    .B(_02319_),
    .Y(_03851_));
 sg13g2_nor3_1 _14214_ (.A(_03849_),
    .B(_03850_),
    .C(_03851_),
    .Y(_03852_));
 sg13g2_o21ai_1 _14215_ (.B1(_03849_),
    .Y(_03853_),
    .A1(_03850_),
    .A2(_03851_));
 sg13g2_nand2_1 _14216_ (.Y(_03854_),
    .A(_05352_),
    .B(net2720));
 sg13g2_nand3_1 _14217_ (.B(net2728),
    .C(_03854_),
    .A(_05011_),
    .Y(_03855_));
 sg13g2_o21ai_1 _14218_ (.B1(_03853_),
    .Y(_03856_),
    .A1(_03852_),
    .A2(_03855_));
 sg13g2_inv_1 _14219_ (.Y(_03857_),
    .A(_03856_));
 sg13g2_nand2_1 _14220_ (.Y(_03858_),
    .A(_03846_),
    .B(_03857_));
 sg13g2_nor2_1 _14221_ (.A(_03846_),
    .B(_03857_),
    .Y(_03859_));
 sg13g2_nor2_1 _14222_ (.A(net2543),
    .B(net2336),
    .Y(_03860_));
 sg13g2_nor2_1 _14223_ (.A(net2787),
    .B(net2634),
    .Y(_03861_));
 sg13g2_xnor2_1 _14224_ (.Y(_03862_),
    .A(_00015_),
    .B(_03861_));
 sg13g2_nand2b_1 _14225_ (.Y(_03863_),
    .B(_03862_),
    .A_N(_03860_));
 sg13g2_nor3_1 _14226_ (.A(net2543),
    .B(net2336),
    .C(_03862_),
    .Y(_03864_));
 sg13g2_nor2_1 _14227_ (.A(net2452),
    .B(net2791),
    .Y(_03865_));
 sg13g2_xor2_1 _14228_ (.B(net2726),
    .A(net2608),
    .X(_03866_));
 sg13g2_xnor2_1 _14229_ (.Y(_03867_),
    .A(_03865_),
    .B(_03866_));
 sg13g2_o21ai_1 _14230_ (.B1(_03863_),
    .Y(_03868_),
    .A1(_03864_),
    .A2(_03867_));
 sg13g2_a21oi_2 _14231_ (.B1(_03859_),
    .Y(_03869_),
    .A2(_03868_),
    .A1(_03858_));
 sg13g2_xnor2_1 _14232_ (.Y(_03870_),
    .A(net2685),
    .B(net2790));
 sg13g2_nand2b_1 _14233_ (.Y(_03871_),
    .B(net2422),
    .A_N(net2244));
 sg13g2_nand2_1 _14234_ (.Y(_03872_),
    .A(net2349),
    .B(net2394));
 sg13g2_xnor2_1 _14235_ (.Y(_03873_),
    .A(_03871_),
    .B(_03872_));
 sg13g2_inv_1 _14236_ (.Y(_03874_),
    .A(_03873_));
 sg13g2_nor2_1 _14237_ (.A(_03870_),
    .B(_03874_),
    .Y(_03875_));
 sg13g2_xnor2_1 _14238_ (.Y(_03876_),
    .A(net2582),
    .B(net2597));
 sg13g2_nor2_1 _14239_ (.A(_03875_),
    .B(_03876_),
    .Y(_03877_));
 sg13g2_a21oi_1 _14240_ (.A1(_03870_),
    .A2(_03874_),
    .Y(_03878_),
    .B1(_03877_));
 sg13g2_nor2b_1 _14241_ (.A(net2720),
    .B_N(net2690),
    .Y(_03879_));
 sg13g2_nor3_1 _14242_ (.A(net2493),
    .B(net2705),
    .C(_03879_),
    .Y(_03880_));
 sg13g2_nand2b_1 _14243_ (.Y(_03881_),
    .B(net2576),
    .A_N(net2592));
 sg13g2_xnor2_1 _14244_ (.Y(_03882_),
    .A(net2756),
    .B(net2685));
 sg13g2_xnor2_1 _14245_ (.Y(_03883_),
    .A(_03881_),
    .B(_03882_));
 sg13g2_or4_1 _14246_ (.A(net2493),
    .B(net2705),
    .C(_03879_),
    .D(_03883_),
    .X(_03884_));
 sg13g2_nand2b_1 _14247_ (.Y(_03885_),
    .B(_03883_),
    .A_N(_03880_));
 sg13g2_xor2_1 _14248_ (.B(net2801),
    .A(net2304),
    .X(_03886_));
 sg13g2_nor2_2 _14249_ (.A(_07893_),
    .B(_03886_),
    .Y(_03887_));
 sg13g2_nand2_1 _14250_ (.Y(_03888_),
    .A(_03884_),
    .B(_03887_));
 sg13g2_nand3_1 _14251_ (.B(_03885_),
    .C(_03888_),
    .A(_03878_),
    .Y(_03889_));
 sg13g2_inv_1 _14252_ (.Y(_03890_),
    .A(_03889_));
 sg13g2_a21oi_1 _14253_ (.A1(_03885_),
    .A2(_03888_),
    .Y(_03891_),
    .B1(_03878_));
 sg13g2_nor2b_1 _14254_ (.A(net2412),
    .B_N(net2686),
    .Y(_03892_));
 sg13g2_xnor2_1 _14255_ (.Y(_03893_),
    .A(net2300),
    .B(_03892_));
 sg13g2_xnor2_1 _14256_ (.Y(_03894_),
    .A(net2245),
    .B(net2410));
 sg13g2_xnor2_1 _14257_ (.Y(_03895_),
    .A(net2716),
    .B(_03894_));
 sg13g2_inv_1 _14258_ (.Y(_03896_),
    .A(_03895_));
 sg13g2_nor2_1 _14259_ (.A(_03893_),
    .B(_03896_),
    .Y(_03897_));
 sg13g2_nand2_1 _14260_ (.Y(_03898_),
    .A(_03893_),
    .B(_03896_));
 sg13g2_nor2_1 _14261_ (.A(net2468),
    .B(net2496),
    .Y(_03899_));
 sg13g2_nand2_1 _14262_ (.Y(_03900_),
    .A(net2809),
    .B(_05616_));
 sg13g2_xnor2_1 _14263_ (.Y(_03901_),
    .A(_03899_),
    .B(_03900_));
 sg13g2_o21ai_1 _14264_ (.B1(_03898_),
    .Y(_03902_),
    .A1(_03897_),
    .A2(_03901_));
 sg13g2_a21oi_2 _14265_ (.B1(_03891_),
    .Y(_03903_),
    .A2(_03902_),
    .A1(_03889_));
 sg13g2_nand2_1 _14266_ (.Y(_03904_),
    .A(_03869_),
    .B(_03903_));
 sg13g2_nor2_1 _14267_ (.A(_03869_),
    .B(_03903_),
    .Y(_03905_));
 sg13g2_xor2_1 _14268_ (.B(_03903_),
    .A(_03869_),
    .X(_03906_));
 sg13g2_nand2_1 _14269_ (.Y(_03907_),
    .A(_05253_),
    .B(net2253));
 sg13g2_xnor2_1 _14270_ (.Y(_03908_),
    .A(net2355),
    .B(net2737));
 sg13g2_xnor2_1 _14271_ (.Y(_03909_),
    .A(_03907_),
    .B(_03908_));
 sg13g2_nor3_1 _14272_ (.A(_05495_),
    .B(net2489),
    .C(_03909_),
    .Y(_03910_));
 sg13g2_o21ai_1 _14273_ (.B1(_03909_),
    .Y(_03911_),
    .A1(_05495_),
    .A2(net2488));
 sg13g2_xor2_1 _14274_ (.B(net2761),
    .A(net2450),
    .X(_03912_));
 sg13g2_o21ai_1 _14275_ (.B1(_03911_),
    .Y(_03913_),
    .A1(_03910_),
    .A2(_03912_));
 sg13g2_nor2b_2 _14276_ (.A(net2337),
    .B_N(net2228),
    .Y(_03914_));
 sg13g2_nor3_1 _14277_ (.A(net2550),
    .B(net2817),
    .C(_03914_),
    .Y(_03915_));
 sg13g2_xor2_1 _14278_ (.B(net2614),
    .A(net2710),
    .X(_03916_));
 sg13g2_nor2b_1 _14279_ (.A(_03915_),
    .B_N(_03916_),
    .Y(_03917_));
 sg13g2_or4_1 _14280_ (.A(net2550),
    .B(net2817),
    .C(_03914_),
    .D(_03916_),
    .X(_03918_));
 sg13g2_xor2_1 _14281_ (.B(net2658),
    .A(net2418),
    .X(_03919_));
 sg13g2_xnor2_1 _14282_ (.Y(_03920_),
    .A(net2323),
    .B(net2310));
 sg13g2_nand2_1 _14283_ (.Y(_03921_),
    .A(_03919_),
    .B(_03920_));
 sg13g2_o21ai_1 _14284_ (.B1(_03918_),
    .Y(_03922_),
    .A1(_03917_),
    .A2(_03921_));
 sg13g2_nor2_1 _14285_ (.A(_03913_),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_nand2_1 _14286_ (.Y(_03924_),
    .A(_03913_),
    .B(_03922_));
 sg13g2_nand2b_2 _14287_ (.Y(_03925_),
    .B(net2376),
    .A_N(net2271));
 sg13g2_nor2_1 _14288_ (.A(_05297_),
    .B(net2463),
    .Y(_03926_));
 sg13g2_xor2_1 _14289_ (.B(net2549),
    .A(net2582),
    .X(_03927_));
 sg13g2_xnor2_1 _14290_ (.Y(_03928_),
    .A(_03926_),
    .B(_03927_));
 sg13g2_nor2_1 _14291_ (.A(_03925_),
    .B(_03928_),
    .Y(_03929_));
 sg13g2_xnor2_1 _14292_ (.Y(_03930_),
    .A(\net.in[108] ),
    .B(net2564));
 sg13g2_a21oi_1 _14293_ (.A1(_03925_),
    .A2(_03928_),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nor2_1 _14294_ (.A(_03929_),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_o21ai_1 _14295_ (.B1(_03924_),
    .Y(_03933_),
    .A1(_03923_),
    .A2(_03932_));
 sg13g2_xnor2_1 _14296_ (.Y(_03934_),
    .A(_03906_),
    .B(_03933_));
 sg13g2_xor2_1 _14297_ (.B(net2562),
    .A(net2613),
    .X(_03935_));
 sg13g2_nand2_1 _14298_ (.Y(_03936_),
    .A(_09246_),
    .B(_03935_));
 sg13g2_or2_1 _14299_ (.X(_03937_),
    .B(_03935_),
    .A(_09246_));
 sg13g2_xor2_1 _14300_ (.B(net2658),
    .A(net2306),
    .X(_03938_));
 sg13g2_a21oi_2 _14301_ (.B1(_03938_),
    .Y(_03939_),
    .A2(_05352_),
    .A1(_05165_));
 sg13g2_nand2_1 _14302_ (.Y(_03940_),
    .A(_03937_),
    .B(_03939_));
 sg13g2_xnor2_1 _14303_ (.Y(_03941_),
    .A(net2526),
    .B(net2365));
 sg13g2_xor2_1 _14304_ (.B(net2815),
    .A(net2275),
    .X(_03942_));
 sg13g2_xor2_1 _14305_ (.B(net2285),
    .A(net2218),
    .X(_03943_));
 sg13g2_o21ai_1 _14306_ (.B1(_03943_),
    .Y(_03944_),
    .A1(_03941_),
    .A2(_03942_));
 sg13g2_nor3_1 _14307_ (.A(_03941_),
    .B(_03942_),
    .C(_03943_),
    .Y(_03945_));
 sg13g2_or3_1 _14308_ (.A(_03941_),
    .B(_03942_),
    .C(_03943_),
    .X(_03946_));
 sg13g2_a21o_2 _14309_ (.A2(net2411),
    .A1(net2181),
    .B1(net2533),
    .X(_03947_));
 sg13g2_a21oi_2 _14310_ (.B1(_03945_),
    .Y(_03948_),
    .A2(_03947_),
    .A1(_03944_));
 sg13g2_nand3_1 _14311_ (.B(_03940_),
    .C(_03948_),
    .A(_03936_),
    .Y(_03949_));
 sg13g2_a21o_1 _14312_ (.A2(_03940_),
    .A1(_03936_),
    .B1(_03948_),
    .X(_03950_));
 sg13g2_xnor2_1 _14313_ (.Y(_03951_),
    .A(net2677),
    .B(net2754));
 sg13g2_a21oi_1 _14314_ (.A1(net2485),
    .A2(_05154_),
    .Y(_03952_),
    .B1(_03951_));
 sg13g2_nand3_1 _14315_ (.B(_05154_),
    .C(_03951_),
    .A(net2484),
    .Y(_03953_));
 sg13g2_xor2_1 _14316_ (.B(net2714),
    .A(net2416),
    .X(_03954_));
 sg13g2_nand2_1 _14317_ (.Y(_03955_),
    .A(net2484),
    .B(_03954_));
 sg13g2_o21ai_1 _14318_ (.B1(_03953_),
    .Y(_03956_),
    .A1(_03952_),
    .A2(_03955_));
 sg13g2_nand2_1 _14319_ (.Y(_03957_),
    .A(_03949_),
    .B(_03956_));
 sg13g2_a21oi_1 _14320_ (.A1(_03950_),
    .A2(_03957_),
    .Y(_03958_),
    .B1(_03934_));
 sg13g2_nand3_1 _14321_ (.B(_03950_),
    .C(_03957_),
    .A(_03934_),
    .Y(_03959_));
 sg13g2_a21oi_2 _14322_ (.B1(_03958_),
    .Y(_03960_),
    .A2(_03959_),
    .A1(_03840_));
 sg13g2_nor2b_1 _14323_ (.A(_03958_),
    .B_N(_03959_),
    .Y(_03961_));
 sg13g2_xnor2_1 _14324_ (.Y(_03962_),
    .A(_03839_),
    .B(_03961_));
 sg13g2_xnor2_1 _14325_ (.Y(_03963_),
    .A(net2638),
    .B(net2651));
 sg13g2_inv_1 _14326_ (.Y(_03964_),
    .A(_03963_));
 sg13g2_nor2_1 _14327_ (.A(net2682),
    .B(net2549),
    .Y(_03965_));
 sg13g2_nor2_1 _14328_ (.A(\net.in[10] ),
    .B(net2756),
    .Y(_03966_));
 sg13g2_xnor2_1 _14329_ (.Y(_03967_),
    .A(_03965_),
    .B(_03966_));
 sg13g2_nor2_1 _14330_ (.A(_03964_),
    .B(_03967_),
    .Y(_03968_));
 sg13g2_nand2_1 _14331_ (.Y(_03969_),
    .A(_03964_),
    .B(_03967_));
 sg13g2_nor2_1 _14332_ (.A(net2212),
    .B(net2774),
    .Y(_03970_));
 sg13g2_o21ai_1 _14333_ (.B1(_03969_),
    .Y(_03971_),
    .A1(_03968_),
    .A2(_03970_));
 sg13g2_nor3_2 _14334_ (.A(net2656),
    .B(net2274),
    .C(_02019_),
    .Y(_03972_));
 sg13g2_and2_1 _14335_ (.A(_09697_),
    .B(_03972_),
    .X(_03973_));
 sg13g2_nor2_1 _14336_ (.A(_09697_),
    .B(_03972_),
    .Y(_03974_));
 sg13g2_xor2_1 _14337_ (.B(net2362),
    .A(net2461),
    .X(_03975_));
 sg13g2_xnor2_1 _14338_ (.Y(_03976_),
    .A(net2624),
    .B(net2714));
 sg13g2_nand2_2 _14339_ (.Y(_03977_),
    .A(_03975_),
    .B(_03976_));
 sg13g2_nor2b_1 _14340_ (.A(_03973_),
    .B_N(_03977_),
    .Y(_03978_));
 sg13g2_nor2_1 _14341_ (.A(_00495_),
    .B(_02713_),
    .Y(_03979_));
 sg13g2_nor2b_1 _14342_ (.A(net2284),
    .B_N(net2468),
    .Y(_03980_));
 sg13g2_nor2_1 _14343_ (.A(net2520),
    .B(net2232),
    .Y(_03981_));
 sg13g2_xnor2_1 _14344_ (.Y(_03982_),
    .A(_03980_),
    .B(_03981_));
 sg13g2_nand2b_1 _14345_ (.Y(_03983_),
    .B(_03982_),
    .A_N(_03979_));
 sg13g2_nor2b_1 _14346_ (.A(_03982_),
    .B_N(_03979_),
    .Y(_03984_));
 sg13g2_nand2_1 _14347_ (.Y(_03985_),
    .A(net2438),
    .B(_05957_));
 sg13g2_nor2_1 _14348_ (.A(net2609),
    .B(net2756),
    .Y(_03986_));
 sg13g2_xnor2_1 _14349_ (.Y(_03987_),
    .A(_03985_),
    .B(_03986_));
 sg13g2_a21oi_2 _14350_ (.B1(_03984_),
    .Y(_03988_),
    .A2(_03987_),
    .A1(_03983_));
 sg13g2_nor3_1 _14351_ (.A(_03974_),
    .B(_03978_),
    .C(_03988_),
    .Y(_03989_));
 sg13g2_o21ai_1 _14352_ (.B1(_03988_),
    .Y(_03990_),
    .A1(_03974_),
    .A2(_03978_));
 sg13g2_nor2b_1 _14353_ (.A(_03989_),
    .B_N(_03990_),
    .Y(_03991_));
 sg13g2_xnor2_1 _14354_ (.Y(_03992_),
    .A(_03971_),
    .B(_03991_));
 sg13g2_xor2_1 _14355_ (.B(_03895_),
    .A(_03893_),
    .X(_03993_));
 sg13g2_xnor2_1 _14356_ (.Y(_03994_),
    .A(_03901_),
    .B(_03993_));
 sg13g2_xor2_1 _14357_ (.B(_03873_),
    .A(_03870_),
    .X(_03995_));
 sg13g2_xnor2_1 _14358_ (.Y(_03996_),
    .A(_03876_),
    .B(_03995_));
 sg13g2_nand2_1 _14359_ (.Y(_03997_),
    .A(_03994_),
    .B(_03996_));
 sg13g2_nor2_1 _14360_ (.A(_03994_),
    .B(_03996_),
    .Y(_03998_));
 sg13g2_or2_1 _14361_ (.X(_03999_),
    .B(_03921_),
    .A(_03918_));
 sg13g2_a22oi_1 _14362_ (.Y(_04000_),
    .B1(_03922_),
    .B2(_03999_),
    .A2(_03921_),
    .A1(_03917_));
 sg13g2_a21oi_2 _14363_ (.B1(_03998_),
    .Y(_04001_),
    .A2(_04000_),
    .A1(_03997_));
 sg13g2_nor2b_1 _14364_ (.A(_03910_),
    .B_N(_03911_),
    .Y(_04002_));
 sg13g2_xnor2_1 _14365_ (.Y(_04003_),
    .A(_03912_),
    .B(_04002_));
 sg13g2_xnor2_1 _14366_ (.Y(_04004_),
    .A(_03925_),
    .B(_03928_));
 sg13g2_xor2_1 _14367_ (.B(_04004_),
    .A(_03930_),
    .X(_04005_));
 sg13g2_nor2_1 _14368_ (.A(_04003_),
    .B(_04005_),
    .Y(_04006_));
 sg13g2_nand2_1 _14369_ (.Y(_04007_),
    .A(_03936_),
    .B(_03937_));
 sg13g2_xor2_1 _14370_ (.B(_04007_),
    .A(_03939_),
    .X(_04008_));
 sg13g2_nor2_1 _14371_ (.A(_04006_),
    .B(_04008_),
    .Y(_04009_));
 sg13g2_a21oi_2 _14372_ (.B1(_04009_),
    .Y(_04010_),
    .A2(_04005_),
    .A1(_04003_));
 sg13g2_nor2_1 _14373_ (.A(_04001_),
    .B(_04010_),
    .Y(_04011_));
 sg13g2_nand2_1 _14374_ (.Y(_04012_),
    .A(_04001_),
    .B(_04010_));
 sg13g2_nand2b_1 _14375_ (.Y(_04013_),
    .B(_04012_),
    .A_N(_04011_));
 sg13g2_nor2b_1 _14376_ (.A(_03952_),
    .B_N(_03953_),
    .Y(_04014_));
 sg13g2_xnor2_1 _14377_ (.Y(_04015_),
    .A(_03955_),
    .B(_04014_));
 sg13g2_nand2_1 _14378_ (.Y(_04016_),
    .A(_03944_),
    .B(_03946_));
 sg13g2_xnor2_1 _14379_ (.Y(_04017_),
    .A(_03947_),
    .B(_04016_));
 sg13g2_nor2_1 _14380_ (.A(_04015_),
    .B(_04017_),
    .Y(_04018_));
 sg13g2_nand2_1 _14381_ (.Y(_04019_),
    .A(_04015_),
    .B(_04017_));
 sg13g2_xnor2_1 _14382_ (.Y(_04020_),
    .A(_03819_),
    .B(_03822_));
 sg13g2_xnor2_1 _14383_ (.Y(_04021_),
    .A(_03827_),
    .B(_04020_));
 sg13g2_o21ai_1 _14384_ (.B1(_04019_),
    .Y(_04022_),
    .A1(_04018_),
    .A2(_04021_));
 sg13g2_xnor2_1 _14385_ (.Y(_04023_),
    .A(_04013_),
    .B(_04022_));
 sg13g2_xor2_1 _14386_ (.B(_03811_),
    .A(_03808_),
    .X(_04024_));
 sg13g2_xnor2_1 _14387_ (.Y(_04025_),
    .A(_03815_),
    .B(_04024_));
 sg13g2_xor2_1 _14388_ (.B(_03834_),
    .A(_03831_),
    .X(_04026_));
 sg13g2_xnor2_1 _14389_ (.Y(_04027_),
    .A(_03836_),
    .B(_04026_));
 sg13g2_inv_1 _14390_ (.Y(_04028_),
    .A(_04027_));
 sg13g2_nand2_1 _14391_ (.Y(_04029_),
    .A(_04025_),
    .B(_04028_));
 sg13g2_nor2_1 _14392_ (.A(_04025_),
    .B(_04028_),
    .Y(_04030_));
 sg13g2_nand2_1 _14393_ (.Y(_04031_),
    .A(net2184),
    .B(net2285));
 sg13g2_nand3b_1 _14394_ (.B(_04031_),
    .C(net2535),
    .Y(_04032_),
    .A_N(net2394));
 sg13g2_nand2_1 _14395_ (.Y(_04033_),
    .A(net2624),
    .B(net2458));
 sg13g2_nor2_1 _14396_ (.A(_05330_),
    .B(net2714),
    .Y(_04034_));
 sg13g2_xnor2_1 _14397_ (.Y(_04035_),
    .A(_04033_),
    .B(_04034_));
 sg13g2_nor2_1 _14398_ (.A(net2499),
    .B(net2365),
    .Y(_04036_));
 sg13g2_xnor2_1 _14399_ (.Y(_04037_),
    .A(_00556_),
    .B(_04036_));
 sg13g2_nor2_1 _14400_ (.A(_04035_),
    .B(_04037_),
    .Y(_04038_));
 sg13g2_nand2_1 _14401_ (.Y(_04039_),
    .A(_04035_),
    .B(_04037_));
 sg13g2_nand2b_1 _14402_ (.Y(_04040_),
    .B(_04039_),
    .A_N(_04038_));
 sg13g2_xnor2_1 _14403_ (.Y(_04041_),
    .A(_04032_),
    .B(_04040_));
 sg13g2_a21oi_1 _14404_ (.A1(_04029_),
    .A2(_04041_),
    .Y(_04042_),
    .B1(_04030_));
 sg13g2_nor2b_1 _14405_ (.A(net2809),
    .B_N(net2530),
    .Y(_04043_));
 sg13g2_xnor2_1 _14406_ (.Y(_04044_),
    .A(net2468),
    .B(_04043_));
 sg13g2_xor2_1 _14407_ (.B(net2754),
    .A(net2750),
    .X(_04045_));
 sg13g2_xnor2_1 _14408_ (.Y(_04046_),
    .A(_02835_),
    .B(_04045_));
 sg13g2_nor2_1 _14409_ (.A(_04044_),
    .B(_04046_),
    .Y(_04047_));
 sg13g2_and2_1 _14410_ (.A(_04044_),
    .B(_04046_),
    .X(_04048_));
 sg13g2_a21oi_2 _14411_ (.B1(_06122_),
    .Y(_04049_),
    .A2(net2438),
    .A1(net2382));
 sg13g2_nor2_1 _14412_ (.A(_04047_),
    .B(_04049_),
    .Y(_04050_));
 sg13g2_or3_1 _14413_ (.A(_04042_),
    .B(_04048_),
    .C(_04050_),
    .X(_04051_));
 sg13g2_o21ai_1 _14414_ (.B1(_04042_),
    .Y(_04052_),
    .A1(_04048_),
    .A2(_04050_));
 sg13g2_inv_1 _14415_ (.Y(_04053_),
    .A(_04052_));
 sg13g2_nand2_1 _14416_ (.Y(_04054_),
    .A(_04051_),
    .B(_04052_));
 sg13g2_nor2_1 _14417_ (.A(net2499),
    .B(net2425),
    .Y(_04055_));
 sg13g2_xnor2_1 _14418_ (.Y(_04056_),
    .A(net2323),
    .B(_04055_));
 sg13g2_xnor2_1 _14419_ (.Y(_04057_),
    .A(net2550),
    .B(net2249));
 sg13g2_nand2_2 _14420_ (.Y(_04058_),
    .A(_02432_),
    .B(_04057_));
 sg13g2_nand2b_1 _14421_ (.Y(_04059_),
    .B(_04056_),
    .A_N(_04058_));
 sg13g2_nor2b_1 _14422_ (.A(_04056_),
    .B_N(_04058_),
    .Y(_04060_));
 sg13g2_xor2_1 _14423_ (.B(net2230),
    .A(net2296),
    .X(_04061_));
 sg13g2_a21oi_2 _14424_ (.B1(_04060_),
    .Y(_04062_),
    .A2(_04061_),
    .A1(_04059_));
 sg13g2_xnor2_1 _14425_ (.Y(_04063_),
    .A(_04054_),
    .B(_04062_));
 sg13g2_and2_1 _14426_ (.A(_04023_),
    .B(_04063_),
    .X(_04064_));
 sg13g2_nor2_1 _14427_ (.A(_04023_),
    .B(_04063_),
    .Y(_04065_));
 sg13g2_nor2_1 _14428_ (.A(_04064_),
    .B(_04065_),
    .Y(_04066_));
 sg13g2_xnor2_1 _14429_ (.Y(_04067_),
    .A(_03992_),
    .B(_04066_));
 sg13g2_nor2b_1 _14430_ (.A(net2743),
    .B_N(net2260),
    .Y(_04068_));
 sg13g2_xnor2_1 _14431_ (.Y(_04069_),
    .A(net2721),
    .B(net2572));
 sg13g2_xnor2_1 _14432_ (.Y(_04070_),
    .A(_04068_),
    .B(_04069_));
 sg13g2_and2_1 _14433_ (.A(net2553),
    .B(net2695),
    .X(_04071_));
 sg13g2_nor2_1 _14434_ (.A(net2553),
    .B(net2695),
    .Y(_04072_));
 sg13g2_nor2b_1 _14435_ (.A(net2762),
    .B_N(net2756),
    .Y(_04073_));
 sg13g2_nor3_2 _14436_ (.A(_04071_),
    .B(_04072_),
    .C(_04073_),
    .Y(_04074_));
 sg13g2_xnor2_1 _14437_ (.Y(_04075_),
    .A(net2588),
    .B(net2602));
 sg13g2_a21o_1 _14438_ (.A2(_04075_),
    .A1(_04074_),
    .B1(_04070_),
    .X(_04076_));
 sg13g2_o21ai_1 _14439_ (.B1(_04076_),
    .Y(_04077_),
    .A1(_04074_),
    .A2(_04075_));
 sg13g2_xnor2_1 _14440_ (.Y(_04078_),
    .A(_04074_),
    .B(_04075_));
 sg13g2_xnor2_1 _14441_ (.Y(_04079_),
    .A(_04070_),
    .B(_04078_));
 sg13g2_a22oi_1 _14442_ (.Y(_04080_),
    .B1(_05748_),
    .B2(net2750),
    .A2(net2372),
    .A1(net2212));
 sg13g2_o21ai_1 _14443_ (.B1(_04080_),
    .Y(_04081_),
    .A1(net2750),
    .A2(_05748_));
 sg13g2_xor2_1 _14444_ (.B(net2762),
    .A(net2608),
    .X(_04082_));
 sg13g2_nor3_2 _14445_ (.A(net2274),
    .B(net2812),
    .C(_04082_),
    .Y(_04083_));
 sg13g2_nor2_1 _14446_ (.A(net2264),
    .B(net2281),
    .Y(_04084_));
 sg13g2_xnor2_1 _14447_ (.Y(_04085_),
    .A(net2345),
    .B(_04084_));
 sg13g2_nand2b_1 _14448_ (.Y(_04086_),
    .B(_04085_),
    .A_N(_04083_));
 sg13g2_nor2b_1 _14449_ (.A(_04085_),
    .B_N(_04083_),
    .Y(_04087_));
 sg13g2_xnor2_1 _14450_ (.Y(_04088_),
    .A(_04083_),
    .B(_04085_));
 sg13g2_xnor2_1 _14451_ (.Y(_04089_),
    .A(_04081_),
    .B(_04088_));
 sg13g2_nand2_1 _14452_ (.Y(_04090_),
    .A(_04079_),
    .B(_04089_));
 sg13g2_nor2_1 _14453_ (.A(_04079_),
    .B(_04089_),
    .Y(_04091_));
 sg13g2_xnor2_1 _14454_ (.Y(_04092_),
    .A(net2734),
    .B(net2597));
 sg13g2_xnor2_1 _14455_ (.Y(_04093_),
    .A(net2720),
    .B(_04092_));
 sg13g2_nor2b_2 _14456_ (.A(net2699),
    .B_N(net2483),
    .Y(_04094_));
 sg13g2_nor3_2 _14457_ (.A(net2535),
    .B(net2319),
    .C(_04094_),
    .Y(_04095_));
 sg13g2_nor2_1 _14458_ (.A(net2435),
    .B(net2212),
    .Y(_04096_));
 sg13g2_nor2_1 _14459_ (.A(_04095_),
    .B(_04096_),
    .Y(_04097_));
 sg13g2_xor2_1 _14460_ (.B(_04096_),
    .A(_04095_),
    .X(_04098_));
 sg13g2_xnor2_1 _14461_ (.Y(_04099_),
    .A(_04093_),
    .B(_04098_));
 sg13g2_a21oi_2 _14462_ (.B1(_04091_),
    .Y(_04100_),
    .A2(_04099_),
    .A1(_04090_));
 sg13g2_xnor2_1 _14463_ (.Y(_04101_),
    .A(_03979_),
    .B(_03982_));
 sg13g2_xnor2_1 _14464_ (.Y(_04102_),
    .A(_03987_),
    .B(_04101_));
 sg13g2_xnor2_1 _14465_ (.Y(_04103_),
    .A(_03963_),
    .B(_03967_));
 sg13g2_xnor2_1 _14466_ (.Y(_04104_),
    .A(_03970_),
    .B(_04103_));
 sg13g2_inv_1 _14467_ (.Y(_04105_),
    .A(_04104_));
 sg13g2_nand2b_1 _14468_ (.Y(_04106_),
    .B(_04104_),
    .A_N(_04102_));
 sg13g2_nand2_1 _14469_ (.Y(_04107_),
    .A(net2471),
    .B(net2505));
 sg13g2_nor2_1 _14470_ (.A(net2180),
    .B(net2271),
    .Y(_04108_));
 sg13g2_xnor2_1 _14471_ (.Y(_04109_),
    .A(_04107_),
    .B(_04108_));
 sg13g2_xnor2_1 _14472_ (.Y(_04110_),
    .A(net2652),
    .B(net2690));
 sg13g2_nor2b_1 _14473_ (.A(net2675),
    .B_N(net2738),
    .Y(_04111_));
 sg13g2_xnor2_1 _14474_ (.Y(_04112_),
    .A(net2609),
    .B(net2726));
 sg13g2_xnor2_1 _14475_ (.Y(_04113_),
    .A(_04111_),
    .B(_04112_));
 sg13g2_nand2_1 _14476_ (.Y(_04114_),
    .A(_04110_),
    .B(_04113_));
 sg13g2_or2_1 _14477_ (.X(_04115_),
    .B(_04113_),
    .A(_04110_));
 sg13g2_nand2_1 _14478_ (.Y(_04116_),
    .A(_04114_),
    .B(_04115_));
 sg13g2_nand2b_1 _14479_ (.Y(_04117_),
    .B(_04115_),
    .A_N(_04109_));
 sg13g2_xor2_1 _14480_ (.B(_04116_),
    .A(_04109_),
    .X(_04118_));
 sg13g2_a21o_1 _14481_ (.A2(_04105_),
    .A1(_04102_),
    .B1(_04118_),
    .X(_04119_));
 sg13g2_a21oi_1 _14482_ (.A1(_04106_),
    .A2(_04119_),
    .Y(_04120_),
    .B1(_04100_));
 sg13g2_nand3_1 _14483_ (.B(_04106_),
    .C(_04119_),
    .A(_04100_),
    .Y(_04121_));
 sg13g2_nor2b_1 _14484_ (.A(_04120_),
    .B_N(_04121_),
    .Y(_04122_));
 sg13g2_a22oi_1 _14485_ (.Y(_04123_),
    .B1(net2281),
    .B2(net2397),
    .A2(_05451_),
    .A1(net2720));
 sg13g2_o21ai_1 _14486_ (.B1(_04123_),
    .Y(_04124_),
    .A1(net2720),
    .A2(_05451_));
 sg13g2_o21ai_1 _14487_ (.B1(net2372),
    .Y(_04125_),
    .A1(net2539),
    .A2(net2365));
 sg13g2_xnor2_1 _14488_ (.Y(_04126_),
    .A(net2520),
    .B(net2368));
 sg13g2_nor3_1 _14489_ (.A(\net.in[112] ),
    .B(_04125_),
    .C(_04126_),
    .Y(_04127_));
 sg13g2_o21ai_1 _14490_ (.B1(_04126_),
    .Y(_04128_),
    .A1(\net.in[112] ),
    .A2(_04125_));
 sg13g2_nand2b_1 _14491_ (.Y(_04129_),
    .B(_04128_),
    .A_N(_04127_));
 sg13g2_o21ai_1 _14492_ (.B1(_04128_),
    .Y(_04130_),
    .A1(_04124_),
    .A2(_04127_));
 sg13g2_inv_1 _14493_ (.Y(_04131_),
    .A(_04130_));
 sg13g2_xnor2_1 _14494_ (.Y(_04132_),
    .A(_04124_),
    .B(_04129_));
 sg13g2_nor2b_1 _14495_ (.A(net2734),
    .B_N(net2372),
    .Y(_04133_));
 sg13g2_or3_2 _14496_ (.A(net2587),
    .B(net2774),
    .C(_04133_),
    .X(_04134_));
 sg13g2_nor2_2 _14497_ (.A(net2606),
    .B(net2362),
    .Y(_04135_));
 sg13g2_xnor2_1 _14498_ (.Y(_04136_),
    .A(net2720),
    .B(net2786));
 sg13g2_xnor2_1 _14499_ (.Y(_04137_),
    .A(_04135_),
    .B(_04136_));
 sg13g2_nand2_1 _14500_ (.Y(_04138_),
    .A(_04134_),
    .B(_04137_));
 sg13g2_xnor2_1 _14501_ (.Y(_04139_),
    .A(_04134_),
    .B(_04137_));
 sg13g2_xnor2_1 _14502_ (.Y(_04140_),
    .A(_06507_),
    .B(_04139_));
 sg13g2_nor2_1 _14503_ (.A(_04132_),
    .B(_04140_),
    .Y(_04141_));
 sg13g2_nand2_1 _14504_ (.Y(_04142_),
    .A(_04132_),
    .B(_04140_));
 sg13g2_nor2b_1 _14505_ (.A(net2431),
    .B_N(net2300),
    .Y(_04143_));
 sg13g2_xnor2_1 _14506_ (.Y(_04144_),
    .A(_00021_),
    .B(_04143_));
 sg13g2_xnor2_1 _14507_ (.Y(_04145_),
    .A(net2471),
    .B(net2572));
 sg13g2_nor2_1 _14508_ (.A(_04144_),
    .B(_04145_),
    .Y(_04146_));
 sg13g2_nand2_1 _14509_ (.Y(_04147_),
    .A(_04144_),
    .B(_04145_));
 sg13g2_nand2b_1 _14510_ (.Y(_04148_),
    .B(_04147_),
    .A_N(_04146_));
 sg13g2_nor2_2 _14511_ (.A(_05176_),
    .B(net2223),
    .Y(_04149_));
 sg13g2_nor2_1 _14512_ (.A(net2224),
    .B(net2731),
    .Y(_04150_));
 sg13g2_xnor2_1 _14513_ (.Y(_04151_),
    .A(_04149_),
    .B(_04150_));
 sg13g2_xnor2_1 _14514_ (.Y(_04152_),
    .A(_04148_),
    .B(_04151_));
 sg13g2_o21ai_1 _14515_ (.B1(_04142_),
    .Y(_04153_),
    .A1(_04141_),
    .A2(_04152_));
 sg13g2_xnor2_1 _14516_ (.Y(_04154_),
    .A(_04122_),
    .B(_04153_));
 sg13g2_nand2b_2 _14517_ (.Y(_04155_),
    .B(net2309),
    .A_N(net2320));
 sg13g2_o21ai_1 _14518_ (.B1(_04155_),
    .Y(_04156_),
    .A1(net2329),
    .A2(net2774));
 sg13g2_nor2b_1 _14519_ (.A(net2264),
    .B_N(net2332),
    .Y(_04157_));
 sg13g2_nor3_2 _14520_ (.A(net2457),
    .B(\net.in[49] ),
    .C(_04157_),
    .Y(_04158_));
 sg13g2_xnor2_1 _14521_ (.Y(_04159_),
    .A(net2380),
    .B(net2496));
 sg13g2_xor2_1 _14522_ (.B(_04159_),
    .A(_04158_),
    .X(_04160_));
 sg13g2_xnor2_1 _14523_ (.Y(_04161_),
    .A(_04156_),
    .B(_04160_));
 sg13g2_nor2_1 _14524_ (.A(net2510),
    .B(net2408),
    .Y(_04162_));
 sg13g2_xor2_1 _14525_ (.B(net2503),
    .A(net2345),
    .X(_04163_));
 sg13g2_nand2b_1 _14526_ (.Y(_04164_),
    .B(_04163_),
    .A_N(_00575_));
 sg13g2_nand2b_1 _14527_ (.Y(_04165_),
    .B(_00575_),
    .A_N(_04163_));
 sg13g2_nand2_1 _14528_ (.Y(_04166_),
    .A(_04164_),
    .B(_04165_));
 sg13g2_xor2_1 _14529_ (.B(_04166_),
    .A(_04162_),
    .X(_04167_));
 sg13g2_nor2_1 _14530_ (.A(_04161_),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_nand2_1 _14531_ (.Y(_04169_),
    .A(_04161_),
    .B(_04167_));
 sg13g2_nand2b_1 _14532_ (.Y(_04170_),
    .B(net2747),
    .A_N(net2777));
 sg13g2_a22oi_1 _14533_ (.Y(_04171_),
    .B1(_05891_),
    .B2(net2777),
    .A2(_05770_),
    .A1(net2431));
 sg13g2_nand2b_1 _14534_ (.Y(_04172_),
    .B(net2521),
    .A_N(net2695));
 sg13g2_xnor2_1 _14535_ (.Y(_04173_),
    .A(_00495_),
    .B(_04172_));
 sg13g2_a21oi_1 _14536_ (.A1(_04170_),
    .A2(_04171_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_nand3_1 _14537_ (.B(_04171_),
    .C(_04173_),
    .A(_04170_),
    .Y(_04175_));
 sg13g2_nor2b_1 _14538_ (.A(_04174_),
    .B_N(_04175_),
    .Y(_04176_));
 sg13g2_xnor2_1 _14539_ (.Y(_04177_),
    .A(net2292),
    .B(net2197));
 sg13g2_xnor2_1 _14540_ (.Y(_04178_),
    .A(_04176_),
    .B(_04177_));
 sg13g2_o21ai_1 _14541_ (.B1(_04169_),
    .Y(_04179_),
    .A1(_04168_),
    .A2(_04178_));
 sg13g2_nor3_2 _14542_ (.A(net2665),
    .B(net2232),
    .C(_06100_),
    .Y(_04180_));
 sg13g2_nor2_1 _14543_ (.A(net2493),
    .B(net2576),
    .Y(_04181_));
 sg13g2_xor2_1 _14544_ (.B(net2572),
    .A(net2300),
    .X(_04182_));
 sg13g2_xnor2_1 _14545_ (.Y(_04183_),
    .A(_04181_),
    .B(_04182_));
 sg13g2_nand2_1 _14546_ (.Y(_04184_),
    .A(_04180_),
    .B(_04183_));
 sg13g2_nor2_1 _14547_ (.A(_04180_),
    .B(_04183_),
    .Y(_04185_));
 sg13g2_xor2_1 _14548_ (.B(_04183_),
    .A(_04180_),
    .X(_04186_));
 sg13g2_nor2_2 _14549_ (.A(net2262),
    .B(_05726_),
    .Y(_04187_));
 sg13g2_xnor2_1 _14550_ (.Y(_04188_),
    .A(_00486_),
    .B(_04187_));
 sg13g2_xnor2_1 _14551_ (.Y(_04189_),
    .A(_04186_),
    .B(_04188_));
 sg13g2_nor2_1 _14552_ (.A(_05847_),
    .B(net2748),
    .Y(_04190_));
 sg13g2_o21ai_1 _14553_ (.B1(_04190_),
    .Y(_04191_),
    .A1(net2301),
    .A2(_05671_));
 sg13g2_xnor2_1 _14554_ (.Y(_04192_),
    .A(net2517),
    .B(net2700));
 sg13g2_xor2_1 _14555_ (.B(net2567),
    .A(net2558),
    .X(_04193_));
 sg13g2_nor2_1 _14556_ (.A(_04192_),
    .B(_04193_),
    .Y(_04194_));
 sg13g2_inv_1 _14557_ (.Y(_04195_),
    .A(_04194_));
 sg13g2_and2_1 _14558_ (.A(_04192_),
    .B(_04193_),
    .X(_04196_));
 sg13g2_nor2_1 _14559_ (.A(_04194_),
    .B(_04196_),
    .Y(_04197_));
 sg13g2_xor2_1 _14560_ (.B(_04197_),
    .A(_04191_),
    .X(_04198_));
 sg13g2_nor2_1 _14561_ (.A(_04189_),
    .B(_04198_),
    .Y(_04199_));
 sg13g2_nand2_1 _14562_ (.Y(_04200_),
    .A(_04189_),
    .B(_04198_));
 sg13g2_nand2_1 _14563_ (.Y(_04201_),
    .A(net2335),
    .B(net2489));
 sg13g2_xor2_1 _14564_ (.B(net2761),
    .A(net2638),
    .X(_04202_));
 sg13g2_nand3_1 _14565_ (.B(_04201_),
    .C(_04202_),
    .A(net2253),
    .Y(_04203_));
 sg13g2_inv_1 _14566_ (.Y(_04204_),
    .A(_04203_));
 sg13g2_a21oi_1 _14567_ (.A1(net2253),
    .A2(_04201_),
    .Y(_04205_),
    .B1(_04202_));
 sg13g2_nor2_1 _14568_ (.A(_04204_),
    .B(_04205_),
    .Y(_04206_));
 sg13g2_xnor2_1 _14569_ (.Y(_04207_),
    .A(net2277),
    .B(net2309));
 sg13g2_xnor2_1 _14570_ (.Y(_04208_),
    .A(_00944_),
    .B(_04207_));
 sg13g2_xnor2_1 _14571_ (.Y(_04209_),
    .A(_04206_),
    .B(_04208_));
 sg13g2_or2_1 _14572_ (.X(_04210_),
    .B(_04209_),
    .A(_04199_));
 sg13g2_nand2_1 _14573_ (.Y(_04211_),
    .A(net2415),
    .B(net2277));
 sg13g2_nor2_1 _14574_ (.A(net2415),
    .B(net2277),
    .Y(_04212_));
 sg13g2_o21ai_1 _14575_ (.B1(_04211_),
    .Y(_04213_),
    .A1(net2434),
    .A2(net2535));
 sg13g2_nor2_1 _14576_ (.A(_04212_),
    .B(_04213_),
    .Y(_04214_));
 sg13g2_xor2_1 _14577_ (.B(net2705),
    .A(net2746),
    .X(_04215_));
 sg13g2_nand2_1 _14578_ (.Y(_04216_),
    .A(_04214_),
    .B(_04215_));
 sg13g2_xnor2_1 _14579_ (.Y(_04217_),
    .A(_04214_),
    .B(_04215_));
 sg13g2_xnor2_1 _14580_ (.Y(_04218_),
    .A(_02505_),
    .B(_04217_));
 sg13g2_nor2b_1 _14581_ (.A(net2754),
    .B_N(net2629),
    .Y(_04219_));
 sg13g2_nor2b_1 _14582_ (.A(net2629),
    .B_N(net2754),
    .Y(_04220_));
 sg13g2_nor2_1 _14583_ (.A(net2510),
    .B(net2503),
    .Y(_04221_));
 sg13g2_nor3_2 _14584_ (.A(_04219_),
    .B(_04220_),
    .C(_04221_),
    .Y(_04222_));
 sg13g2_nand2b_1 _14585_ (.Y(_04223_),
    .B(net2341),
    .A_N(net2253));
 sg13g2_nand2_1 _14586_ (.Y(_04224_),
    .A(net2539),
    .B(net2492));
 sg13g2_xnor2_1 _14587_ (.Y(_04225_),
    .A(_04223_),
    .B(_04224_));
 sg13g2_nor2b_1 _14588_ (.A(_04225_),
    .B_N(_04222_),
    .Y(_04226_));
 sg13g2_nand2b_1 _14589_ (.Y(_04227_),
    .B(_04225_),
    .A_N(_04222_));
 sg13g2_nor2b_1 _14590_ (.A(_04226_),
    .B_N(_04227_),
    .Y(_04228_));
 sg13g2_xor2_1 _14591_ (.B(net2376),
    .A(net2296),
    .X(_04229_));
 sg13g2_xnor2_1 _14592_ (.Y(_04230_),
    .A(_04228_),
    .B(_04229_));
 sg13g2_nand2_1 _14593_ (.Y(_04231_),
    .A(_04218_),
    .B(_04230_));
 sg13g2_nor2_1 _14594_ (.A(_04218_),
    .B(_04230_),
    .Y(_04232_));
 sg13g2_nor2b_1 _14595_ (.A(net2638),
    .B_N(net2365),
    .Y(_04233_));
 sg13g2_xnor2_1 _14596_ (.Y(_04234_),
    .A(_00023_),
    .B(_04233_));
 sg13g2_nor2b_1 _14597_ (.A(net2609),
    .B_N(net2509),
    .Y(_04235_));
 sg13g2_nor2_1 _14598_ (.A(net2624),
    .B(net2748),
    .Y(_04236_));
 sg13g2_xnor2_1 _14599_ (.Y(_04237_),
    .A(_04235_),
    .B(_04236_));
 sg13g2_nand2_1 _14600_ (.Y(_04238_),
    .A(net2516),
    .B(net2603));
 sg13g2_xor2_1 _14601_ (.B(_04238_),
    .A(_09158_),
    .X(_04239_));
 sg13g2_nand2_1 _14602_ (.Y(_04240_),
    .A(_04237_),
    .B(_04239_));
 sg13g2_nor2_1 _14603_ (.A(_04237_),
    .B(_04239_),
    .Y(_04241_));
 sg13g2_xor2_1 _14604_ (.B(_04239_),
    .A(_04237_),
    .X(_04242_));
 sg13g2_xor2_1 _14605_ (.B(_04242_),
    .A(_04234_),
    .X(_04243_));
 sg13g2_a21oi_2 _14606_ (.B1(_04232_),
    .Y(_04244_),
    .A2(_04243_),
    .A1(_04231_));
 sg13g2_a21o_1 _14607_ (.A2(_04210_),
    .A1(_04200_),
    .B1(_04244_),
    .X(_04245_));
 sg13g2_nand3_1 _14608_ (.B(_04210_),
    .C(_04244_),
    .A(_04200_),
    .Y(_04246_));
 sg13g2_nand2_1 _14609_ (.Y(_04247_),
    .A(_04245_),
    .B(_04246_));
 sg13g2_nand2b_1 _14610_ (.Y(_04248_),
    .B(_04245_),
    .A_N(_04179_));
 sg13g2_xor2_1 _14611_ (.B(_04247_),
    .A(_04179_),
    .X(_04249_));
 sg13g2_nor2_1 _14612_ (.A(_04154_),
    .B(_04249_),
    .Y(_04250_));
 sg13g2_xor2_1 _14613_ (.B(_04249_),
    .A(_04154_),
    .X(_04251_));
 sg13g2_xnor2_1 _14614_ (.Y(_04252_),
    .A(net2816),
    .B(net2605));
 sg13g2_xnor2_1 _14615_ (.Y(_04253_),
    .A(net2404),
    .B(net2226));
 sg13g2_nand2_1 _14616_ (.Y(_04254_),
    .A(_04252_),
    .B(_04253_));
 sg13g2_nand3_1 _14617_ (.B(net2425),
    .C(net2582),
    .A(net2322),
    .Y(_04255_));
 sg13g2_a21o_1 _14618_ (.A2(net2582),
    .A1(net2425),
    .B1(net2322),
    .X(_04256_));
 sg13g2_xor2_1 _14619_ (.B(net2503),
    .A(net2336),
    .X(_04257_));
 sg13g2_nand3_1 _14620_ (.B(_04256_),
    .C(_04257_),
    .A(_04255_),
    .Y(_04258_));
 sg13g2_a21oi_1 _14621_ (.A1(_04255_),
    .A2(_04256_),
    .Y(_04259_),
    .B1(_04257_));
 sg13g2_a21o_1 _14622_ (.A2(_04256_),
    .A1(_04255_),
    .B1(_04257_),
    .X(_04260_));
 sg13g2_nand2_1 _14623_ (.Y(_04261_),
    .A(_04258_),
    .B(_04260_));
 sg13g2_o21ai_1 _14624_ (.B1(_04258_),
    .Y(_04262_),
    .A1(_04254_),
    .A2(_04259_));
 sg13g2_xnor2_1 _14625_ (.Y(_04263_),
    .A(_04254_),
    .B(_04261_));
 sg13g2_or3_1 _14626_ (.A(net2260),
    .B(net2232),
    .C(_04202_),
    .X(_04264_));
 sg13g2_nor2b_1 _14627_ (.A(net2767),
    .B_N(net2644),
    .Y(_04265_));
 sg13g2_xnor2_1 _14628_ (.Y(_04266_),
    .A(_00001_),
    .B(_04265_));
 sg13g2_nand3_1 _14629_ (.B(_05825_),
    .C(_02702_),
    .A(net2180),
    .Y(_04267_));
 sg13g2_nor2b_1 _14630_ (.A(_04266_),
    .B_N(_04267_),
    .Y(_04268_));
 sg13g2_nand2b_1 _14631_ (.Y(_04269_),
    .B(_04266_),
    .A_N(_04267_));
 sg13g2_xor2_1 _14632_ (.B(_04267_),
    .A(_04266_),
    .X(_04270_));
 sg13g2_xnor2_1 _14633_ (.Y(_04271_),
    .A(_04264_),
    .B(_04270_));
 sg13g2_nor2_1 _14634_ (.A(_04263_),
    .B(_04271_),
    .Y(_04272_));
 sg13g2_xor2_1 _14635_ (.B(\net.in[161] ),
    .A(net2432),
    .X(_04273_));
 sg13g2_xnor2_1 _14636_ (.Y(_04274_),
    .A(net2550),
    .B(\net.in[11] ));
 sg13g2_nand2_1 _14637_ (.Y(_04275_),
    .A(_04273_),
    .B(_04274_));
 sg13g2_xor2_1 _14638_ (.B(net2468),
    .A(net2357),
    .X(_04276_));
 sg13g2_nand3b_1 _14639_ (.B(_05297_),
    .C(_05242_),
    .Y(_04277_),
    .A_N(_04276_));
 sg13g2_o21ai_1 _14640_ (.B1(_04276_),
    .Y(_04278_),
    .A1(net2526),
    .A2(net2444));
 sg13g2_nand2_1 _14641_ (.Y(_04279_),
    .A(_04277_),
    .B(_04278_));
 sg13g2_xor2_1 _14642_ (.B(_04279_),
    .A(_04275_),
    .X(_04280_));
 sg13g2_nor2_1 _14643_ (.A(_04272_),
    .B(_04280_),
    .Y(_04281_));
 sg13g2_a21oi_2 _14644_ (.B1(_04281_),
    .Y(_04282_),
    .A2(_04271_),
    .A1(_04263_));
 sg13g2_nor2_1 _14645_ (.A(net2752),
    .B(_05297_),
    .Y(_04283_));
 sg13g2_xor2_1 _14646_ (.B(net2614),
    .A(net2728),
    .X(_04284_));
 sg13g2_a21oi_2 _14647_ (.B1(_04284_),
    .Y(_04285_),
    .A2(_05891_),
    .A1(net2179));
 sg13g2_xnor2_1 _14648_ (.Y(_04286_),
    .A(net2756),
    .B(net2634));
 sg13g2_xor2_1 _14649_ (.B(_04286_),
    .A(_04285_),
    .X(_04287_));
 sg13g2_xnor2_1 _14650_ (.Y(_04288_),
    .A(_04283_),
    .B(_04287_));
 sg13g2_nor2_1 _14651_ (.A(net2181),
    .B(net2758),
    .Y(_04289_));
 sg13g2_xnor2_1 _14652_ (.Y(_04290_),
    .A(_00009_),
    .B(_04289_));
 sg13g2_xnor2_1 _14653_ (.Y(_04291_),
    .A(net2406),
    .B(\net.in[215] ));
 sg13g2_and3_1 _14654_ (.X(_04292_),
    .A(net2372),
    .B(_06012_),
    .C(_04291_));
 sg13g2_nor2_1 _14655_ (.A(net2588),
    .B(net2581),
    .Y(_04293_));
 sg13g2_xnor2_1 _14656_ (.Y(_04294_),
    .A(net2421),
    .B(_04293_));
 sg13g2_nand2b_1 _14657_ (.Y(_04295_),
    .B(_04294_),
    .A_N(_04292_));
 sg13g2_nor2b_1 _14658_ (.A(_04294_),
    .B_N(_04292_),
    .Y(_04296_));
 sg13g2_xnor2_1 _14659_ (.Y(_04297_),
    .A(_04292_),
    .B(_04294_));
 sg13g2_xnor2_1 _14660_ (.Y(_04298_),
    .A(_04290_),
    .B(_04297_));
 sg13g2_nand2_1 _14661_ (.Y(_04299_),
    .A(_04288_),
    .B(_04298_));
 sg13g2_or2_1 _14662_ (.X(_04300_),
    .B(_04298_),
    .A(_04288_));
 sg13g2_nand2b_1 _14663_ (.Y(_04301_),
    .B(_03853_),
    .A_N(_03852_));
 sg13g2_xnor2_1 _14664_ (.Y(_04302_),
    .A(_03855_),
    .B(_04301_));
 sg13g2_nand2_1 _14665_ (.Y(_04303_),
    .A(_04300_),
    .B(_04302_));
 sg13g2_and3_1 _14666_ (.X(_04304_),
    .A(_04282_),
    .B(_04299_),
    .C(_04303_));
 sg13g2_inv_1 _14667_ (.Y(_04305_),
    .A(_04304_));
 sg13g2_a21oi_1 _14668_ (.A1(_04299_),
    .A2(_04303_),
    .Y(_04306_),
    .B1(_04282_));
 sg13g2_nor2_1 _14669_ (.A(_04304_),
    .B(_04306_),
    .Y(_04307_));
 sg13g2_xor2_1 _14670_ (.B(_03862_),
    .A(_03860_),
    .X(_04308_));
 sg13g2_xnor2_1 _14671_ (.Y(_04309_),
    .A(_03867_),
    .B(_04308_));
 sg13g2_xor2_1 _14672_ (.B(_03841_),
    .A(_09158_),
    .X(_04310_));
 sg13g2_xnor2_1 _14673_ (.Y(_04311_),
    .A(_03844_),
    .B(_04310_));
 sg13g2_inv_1 _14674_ (.Y(_04312_),
    .A(_04311_));
 sg13g2_nor2_1 _14675_ (.A(_04309_),
    .B(_04312_),
    .Y(_04313_));
 sg13g2_nand2_1 _14676_ (.Y(_04314_),
    .A(_04309_),
    .B(_04312_));
 sg13g2_and2_1 _14677_ (.A(_03884_),
    .B(_03885_),
    .X(_04315_));
 sg13g2_xor2_1 _14678_ (.B(_04315_),
    .A(_03887_),
    .X(_04316_));
 sg13g2_o21ai_1 _14679_ (.B1(_04314_),
    .Y(_04317_),
    .A1(_04313_),
    .A2(_04316_));
 sg13g2_xnor2_1 _14680_ (.Y(_04318_),
    .A(_04307_),
    .B(_04317_));
 sg13g2_xnor2_1 _14681_ (.Y(_04319_),
    .A(_04251_),
    .B(_04318_));
 sg13g2_xnor2_1 _14682_ (.Y(_04320_),
    .A(_03994_),
    .B(_03996_));
 sg13g2_xnor2_1 _14683_ (.Y(_04321_),
    .A(_04000_),
    .B(_04320_));
 sg13g2_xnor2_1 _14684_ (.Y(_04322_),
    .A(_04309_),
    .B(_04312_));
 sg13g2_xnor2_1 _14685_ (.Y(_04323_),
    .A(_04316_),
    .B(_04322_));
 sg13g2_nor2_1 _14686_ (.A(_04321_),
    .B(_04323_),
    .Y(_04324_));
 sg13g2_nand2_1 _14687_ (.Y(_04325_),
    .A(_04321_),
    .B(_04323_));
 sg13g2_nor2b_1 _14688_ (.A(_04324_),
    .B_N(_04325_),
    .Y(_04326_));
 sg13g2_xor2_1 _14689_ (.B(_04005_),
    .A(_04003_),
    .X(_04327_));
 sg13g2_xnor2_1 _14690_ (.Y(_04328_),
    .A(_04008_),
    .B(_04327_));
 sg13g2_inv_1 _14691_ (.Y(_04329_),
    .A(_04328_));
 sg13g2_xnor2_1 _14692_ (.Y(_04330_),
    .A(_04326_),
    .B(_04328_));
 sg13g2_xor2_1 _14693_ (.B(_04027_),
    .A(_04025_),
    .X(_04331_));
 sg13g2_xnor2_1 _14694_ (.Y(_04332_),
    .A(_04041_),
    .B(_04331_));
 sg13g2_nand2b_1 _14695_ (.Y(_04333_),
    .B(_04019_),
    .A_N(_04018_));
 sg13g2_xnor2_1 _14696_ (.Y(_04334_),
    .A(_04021_),
    .B(_04333_));
 sg13g2_nor2_1 _14697_ (.A(_04332_),
    .B(_04334_),
    .Y(_04335_));
 sg13g2_nor2_1 _14698_ (.A(net2418),
    .B(_04335_),
    .Y(_04336_));
 sg13g2_a21oi_1 _14699_ (.A1(_04332_),
    .A2(_04334_),
    .Y(_04337_),
    .B1(_04336_));
 sg13g2_xor2_1 _14700_ (.B(_04334_),
    .A(_04332_),
    .X(_04338_));
 sg13g2_xnor2_1 _14701_ (.Y(_04339_),
    .A(net2418),
    .B(_04338_));
 sg13g2_nor2_1 _14702_ (.A(_04330_),
    .B(_04339_),
    .Y(_04340_));
 sg13g2_xor2_1 _14703_ (.B(_04339_),
    .A(_04330_),
    .X(_04341_));
 sg13g2_xnor2_1 _14704_ (.Y(_04342_),
    .A(_04132_),
    .B(_04140_));
 sg13g2_xnor2_1 _14705_ (.Y(_04343_),
    .A(_04152_),
    .B(_04342_));
 sg13g2_xnor2_1 _14706_ (.Y(_04344_),
    .A(_04189_),
    .B(_04198_));
 sg13g2_xnor2_1 _14707_ (.Y(_04345_),
    .A(_04209_),
    .B(_04344_));
 sg13g2_nand2_1 _14708_ (.Y(_04346_),
    .A(_04343_),
    .B(_04345_));
 sg13g2_nor2_1 _14709_ (.A(_04343_),
    .B(_04345_),
    .Y(_04347_));
 sg13g2_xnor2_1 _14710_ (.Y(_04348_),
    .A(_04343_),
    .B(_04345_));
 sg13g2_xnor2_1 _14711_ (.Y(_04349_),
    .A(_04218_),
    .B(_04230_));
 sg13g2_xnor2_1 _14712_ (.Y(_04350_),
    .A(_04243_),
    .B(_04349_));
 sg13g2_xnor2_1 _14713_ (.Y(_04351_),
    .A(_04348_),
    .B(_04350_));
 sg13g2_or2_1 _14714_ (.X(_04352_),
    .B(_04099_),
    .A(_04090_));
 sg13g2_a22oi_1 _14715_ (.Y(_04353_),
    .B1(_04100_),
    .B2(_04352_),
    .A2(_04099_),
    .A1(_04091_));
 sg13g2_xnor2_1 _14716_ (.Y(_04354_),
    .A(_04102_),
    .B(_04104_));
 sg13g2_xnor2_1 _14717_ (.Y(_04355_),
    .A(_04118_),
    .B(_04354_));
 sg13g2_nor2_1 _14718_ (.A(_03973_),
    .B(_03974_),
    .Y(_04356_));
 sg13g2_xor2_1 _14719_ (.B(_04356_),
    .A(_03977_),
    .X(_04357_));
 sg13g2_xor2_1 _14720_ (.B(_04046_),
    .A(_04044_),
    .X(_04358_));
 sg13g2_xnor2_1 _14721_ (.Y(_04359_),
    .A(_04049_),
    .B(_04358_));
 sg13g2_xnor2_1 _14722_ (.Y(_04360_),
    .A(_04056_),
    .B(_04058_));
 sg13g2_xnor2_1 _14723_ (.Y(_04361_),
    .A(_04061_),
    .B(_04360_));
 sg13g2_nor2_1 _14724_ (.A(_04359_),
    .B(_04361_),
    .Y(_04362_));
 sg13g2_nand2_1 _14725_ (.Y(_04363_),
    .A(_04359_),
    .B(_04361_));
 sg13g2_xor2_1 _14726_ (.B(_04361_),
    .A(_04359_),
    .X(_04364_));
 sg13g2_xnor2_1 _14727_ (.Y(_04365_),
    .A(_04357_),
    .B(_04364_));
 sg13g2_nand2_1 _14728_ (.Y(_04366_),
    .A(_04355_),
    .B(_04365_));
 sg13g2_nor2_1 _14729_ (.A(_04355_),
    .B(_04365_),
    .Y(_04367_));
 sg13g2_xnor2_1 _14730_ (.Y(_04368_),
    .A(_04355_),
    .B(_04365_));
 sg13g2_xor2_1 _14731_ (.B(_04368_),
    .A(_04353_),
    .X(_04369_));
 sg13g2_nor2_1 _14732_ (.A(_04351_),
    .B(_04369_),
    .Y(_04370_));
 sg13g2_nand2_1 _14733_ (.Y(_04371_),
    .A(_04351_),
    .B(_04369_));
 sg13g2_xor2_1 _14734_ (.B(_04369_),
    .A(_04351_),
    .X(_04372_));
 sg13g2_xnor2_1 _14735_ (.Y(_04373_),
    .A(_04161_),
    .B(_04167_));
 sg13g2_xnor2_1 _14736_ (.Y(_04374_),
    .A(_04178_),
    .B(_04373_));
 sg13g2_xnor2_1 _14737_ (.Y(_04375_),
    .A(_04263_),
    .B(_04271_));
 sg13g2_xor2_1 _14738_ (.B(_04375_),
    .A(_04280_),
    .X(_04376_));
 sg13g2_nor2_1 _14739_ (.A(_04374_),
    .B(_04376_),
    .Y(_04377_));
 sg13g2_nand2_1 _14740_ (.Y(_04378_),
    .A(_04374_),
    .B(_04376_));
 sg13g2_nor2b_1 _14741_ (.A(_04377_),
    .B_N(_04378_),
    .Y(_04379_));
 sg13g2_nand2_1 _14742_ (.Y(_04380_),
    .A(_04299_),
    .B(_04300_));
 sg13g2_xor2_1 _14743_ (.B(_04380_),
    .A(_04302_),
    .X(_04381_));
 sg13g2_xnor2_1 _14744_ (.Y(_04382_),
    .A(_04379_),
    .B(_04381_));
 sg13g2_xnor2_1 _14745_ (.Y(_04383_),
    .A(_04372_),
    .B(_04382_));
 sg13g2_a21oi_2 _14746_ (.B1(_04340_),
    .Y(_04384_),
    .A2(_04383_),
    .A1(_04341_));
 sg13g2_o21ai_1 _14747_ (.B1(_04371_),
    .Y(_04385_),
    .A1(_04370_),
    .A2(_04382_));
 sg13g2_nor2b_1 _14748_ (.A(_04384_),
    .B_N(_04385_),
    .Y(_04386_));
 sg13g2_xnor2_1 _14749_ (.Y(_04387_),
    .A(_04384_),
    .B(_04385_));
 sg13g2_o21ai_1 _14750_ (.B1(_04346_),
    .Y(_04388_),
    .A1(_04347_),
    .A2(_04350_));
 sg13g2_o21ai_1 _14751_ (.B1(_04366_),
    .Y(_04389_),
    .A1(_04353_),
    .A2(_04367_));
 sg13g2_nand2b_1 _14752_ (.Y(_04390_),
    .B(_04389_),
    .A_N(_04388_));
 sg13g2_inv_1 _14753_ (.Y(_04391_),
    .A(_04390_));
 sg13g2_nor2b_1 _14754_ (.A(_04389_),
    .B_N(_04388_),
    .Y(_04392_));
 sg13g2_nor2_1 _14755_ (.A(_04391_),
    .B(_04392_),
    .Y(_04393_));
 sg13g2_a21oi_2 _14756_ (.B1(_04377_),
    .Y(_04394_),
    .A2(_04381_),
    .A1(_04378_));
 sg13g2_xnor2_1 _14757_ (.Y(_04395_),
    .A(_04393_),
    .B(_04394_));
 sg13g2_nand2_1 _14758_ (.Y(_04396_),
    .A(_04387_),
    .B(_04395_));
 sg13g2_nor2_1 _14759_ (.A(_04387_),
    .B(_04395_),
    .Y(_04397_));
 sg13g2_xnor2_1 _14760_ (.Y(_04398_),
    .A(_04387_),
    .B(_04395_));
 sg13g2_o21ai_1 _14761_ (.B1(_04363_),
    .Y(_04399_),
    .A1(_04357_),
    .A2(_04362_));
 sg13g2_o21ai_1 _14762_ (.B1(_04325_),
    .Y(_04400_),
    .A1(_04324_),
    .A2(_04329_));
 sg13g2_and2_1 _14763_ (.A(_04337_),
    .B(_04400_),
    .X(_04401_));
 sg13g2_or2_1 _14764_ (.X(_04402_),
    .B(_04400_),
    .A(_04337_));
 sg13g2_nor2b_1 _14765_ (.A(_04401_),
    .B_N(_04402_),
    .Y(_04403_));
 sg13g2_xnor2_1 _14766_ (.Y(_04404_),
    .A(_04399_),
    .B(_04403_));
 sg13g2_xnor2_1 _14767_ (.Y(_04405_),
    .A(_04398_),
    .B(_04404_));
 sg13g2_nand2_1 _14768_ (.Y(_04406_),
    .A(_04319_),
    .B(_04405_));
 sg13g2_xor2_1 _14769_ (.B(_04405_),
    .A(_04319_),
    .X(_04407_));
 sg13g2_xnor2_1 _14770_ (.Y(_04408_),
    .A(_04067_),
    .B(_04407_));
 sg13g2_a21oi_1 _14771_ (.A1(_04234_),
    .A2(_04240_),
    .Y(_04409_),
    .B1(_04241_));
 sg13g2_nand2b_1 _14772_ (.Y(_04410_),
    .B(_04165_),
    .A_N(_04162_));
 sg13g2_nand3_1 _14773_ (.B(_04409_),
    .C(_04410_),
    .A(_04164_),
    .Y(_04411_));
 sg13g2_a21o_1 _14774_ (.A2(_04410_),
    .A1(_04164_),
    .B1(_04409_),
    .X(_04412_));
 sg13g2_nand2_1 _14775_ (.Y(_04413_),
    .A(_04411_),
    .B(_04412_));
 sg13g2_a21o_1 _14776_ (.A2(_04159_),
    .A1(_04158_),
    .B1(_04156_),
    .X(_04414_));
 sg13g2_o21ai_1 _14777_ (.B1(_04414_),
    .Y(_04415_),
    .A1(_04158_),
    .A2(_04159_));
 sg13g2_nor2b_1 _14778_ (.A(_04415_),
    .B_N(_04412_),
    .Y(_04416_));
 sg13g2_inv_1 _14779_ (.Y(_04417_),
    .A(_04416_));
 sg13g2_a22oi_1 _14780_ (.Y(_04418_),
    .B1(_04416_),
    .B2(_04411_),
    .A2(_04415_),
    .A1(_04413_));
 sg13g2_o21ai_1 _14781_ (.B1(_04203_),
    .Y(_04419_),
    .A1(_04205_),
    .A2(_04208_));
 sg13g2_o21ai_1 _14782_ (.B1(_04227_),
    .Y(_04420_),
    .A1(_04226_),
    .A2(_04229_));
 sg13g2_nand2_1 _14783_ (.Y(_04421_),
    .A(_04419_),
    .B(_04420_));
 sg13g2_nor2_1 _14784_ (.A(_04419_),
    .B(_04420_),
    .Y(_04422_));
 sg13g2_xor2_1 _14785_ (.B(_04420_),
    .A(_04419_),
    .X(_04423_));
 sg13g2_o21ai_1 _14786_ (.B1(_02504_),
    .Y(_04424_),
    .A1(_04214_),
    .A2(_04215_));
 sg13g2_nand2_2 _14787_ (.Y(_04425_),
    .A(_04216_),
    .B(_04424_));
 sg13g2_xnor2_1 _14788_ (.Y(_04426_),
    .A(_04423_),
    .B(_04425_));
 sg13g2_nand2_1 _14789_ (.Y(_04427_),
    .A(_04418_),
    .B(_04426_));
 sg13g2_nor2_1 _14790_ (.A(_04418_),
    .B(_04426_),
    .Y(_04428_));
 sg13g2_xor2_1 _14791_ (.B(_04426_),
    .A(_04418_),
    .X(_04429_));
 sg13g2_o21ai_1 _14792_ (.B1(_04175_),
    .Y(_04430_),
    .A1(_04174_),
    .A2(_04177_));
 sg13g2_o21ai_1 _14793_ (.B1(_04269_),
    .Y(_04431_),
    .A1(_04264_),
    .A2(_04268_));
 sg13g2_nand2b_1 _14794_ (.Y(_04432_),
    .B(_04430_),
    .A_N(_04431_));
 sg13g2_nor2b_1 _14795_ (.A(_04430_),
    .B_N(_04431_),
    .Y(_04433_));
 sg13g2_xor2_1 _14796_ (.B(_04431_),
    .A(_04430_),
    .X(_04434_));
 sg13g2_xnor2_1 _14797_ (.Y(_04435_),
    .A(_04262_),
    .B(_04434_));
 sg13g2_xnor2_1 _14798_ (.Y(_04436_),
    .A(_04429_),
    .B(_04435_));
 sg13g2_o21ai_1 _14799_ (.B1(_06507_),
    .Y(_04437_),
    .A1(_04134_),
    .A2(_04137_));
 sg13g2_a21oi_1 _14800_ (.A1(_04095_),
    .A2(_04096_),
    .Y(_04438_),
    .B1(_04093_));
 sg13g2_nor2_1 _14801_ (.A(_04097_),
    .B(_04438_),
    .Y(_04439_));
 sg13g2_and3_1 _14802_ (.X(_04440_),
    .A(_04138_),
    .B(_04437_),
    .C(_04439_));
 sg13g2_nand3_1 _14803_ (.B(_04437_),
    .C(_04439_),
    .A(_04138_),
    .Y(_04441_));
 sg13g2_a21oi_1 _14804_ (.A1(_04138_),
    .A2(_04437_),
    .Y(_04442_),
    .B1(_04439_));
 sg13g2_o21ai_1 _14805_ (.B1(_04441_),
    .Y(_04443_),
    .A1(_04131_),
    .A2(_04442_));
 sg13g2_a21oi_1 _14806_ (.A1(_04131_),
    .A2(_04442_),
    .Y(_04444_),
    .B1(_04443_));
 sg13g2_a21oi_2 _14807_ (.B1(_04444_),
    .Y(_04445_),
    .A2(_04440_),
    .A1(_04130_));
 sg13g2_a21oi_1 _14808_ (.A1(_04114_),
    .A2(_04117_),
    .Y(_04446_),
    .B1(_04077_));
 sg13g2_nand3_1 _14809_ (.B(_04114_),
    .C(_04117_),
    .A(_04077_),
    .Y(_04447_));
 sg13g2_nand2b_1 _14810_ (.Y(_04448_),
    .B(_04447_),
    .A_N(_04446_));
 sg13g2_a21oi_1 _14811_ (.A1(_04081_),
    .A2(_04086_),
    .Y(_04449_),
    .B1(_04087_));
 sg13g2_xnor2_1 _14812_ (.Y(_04450_),
    .A(_04448_),
    .B(_04449_));
 sg13g2_nand2b_1 _14813_ (.Y(_04451_),
    .B(_04450_),
    .A_N(_04445_));
 sg13g2_nand2b_1 _14814_ (.Y(_04452_),
    .B(_04445_),
    .A_N(_04450_));
 sg13g2_nand2_1 _14815_ (.Y(_04453_),
    .A(_04451_),
    .B(_04452_));
 sg13g2_a21oi_2 _14816_ (.B1(_04185_),
    .Y(_04454_),
    .A2(_04188_),
    .A1(_04184_));
 sg13g2_o21ai_1 _14817_ (.B1(_04147_),
    .Y(_04455_),
    .A1(_04146_),
    .A2(_04151_));
 sg13g2_nand2_1 _14818_ (.Y(_04456_),
    .A(_04454_),
    .B(_04455_));
 sg13g2_xor2_1 _14819_ (.B(_04455_),
    .A(_04454_),
    .X(_04457_));
 sg13g2_o21ai_1 _14820_ (.B1(_04195_),
    .Y(_04458_),
    .A1(_04191_),
    .A2(_04196_));
 sg13g2_xnor2_1 _14821_ (.Y(_04459_),
    .A(_04457_),
    .B(_04458_));
 sg13g2_xor2_1 _14822_ (.B(_04459_),
    .A(_04453_),
    .X(_04460_));
 sg13g2_nand2_1 _14823_ (.Y(_04461_),
    .A(_04436_),
    .B(_04460_));
 sg13g2_nor2_1 _14824_ (.A(_04436_),
    .B(_04460_),
    .Y(_04462_));
 sg13g2_xnor2_1 _14825_ (.Y(_04463_),
    .A(_04436_),
    .B(_04460_));
 sg13g2_nor2_1 _14826_ (.A(_03890_),
    .B(_03891_),
    .Y(_04464_));
 sg13g2_xnor2_1 _14827_ (.Y(_04465_),
    .A(_03902_),
    .B(_04464_));
 sg13g2_xnor2_1 _14828_ (.Y(_04466_),
    .A(_03846_),
    .B(_03856_));
 sg13g2_xnor2_1 _14829_ (.Y(_04467_),
    .A(_03868_),
    .B(_04466_));
 sg13g2_inv_1 _14830_ (.Y(_04468_),
    .A(_04467_));
 sg13g2_nand2_1 _14831_ (.Y(_04469_),
    .A(_04275_),
    .B(_04278_));
 sg13g2_nand2_2 _14832_ (.Y(_04470_),
    .A(_04277_),
    .B(_04469_));
 sg13g2_a21oi_2 _14833_ (.B1(_04296_),
    .Y(_04471_),
    .A2(_04295_),
    .A1(_04290_));
 sg13g2_nand2_1 _14834_ (.Y(_04472_),
    .A(_04470_),
    .B(_04471_));
 sg13g2_xor2_1 _14835_ (.B(_04471_),
    .A(_04470_),
    .X(_04473_));
 sg13g2_a21o_1 _14836_ (.A2(_04286_),
    .A1(_04285_),
    .B1(_04283_),
    .X(_04474_));
 sg13g2_o21ai_1 _14837_ (.B1(_04474_),
    .Y(_04475_),
    .A1(_04285_),
    .A2(_04286_));
 sg13g2_xnor2_1 _14838_ (.Y(_04476_),
    .A(_04473_),
    .B(_04475_));
 sg13g2_nand2_1 _14839_ (.Y(_04477_),
    .A(_04468_),
    .B(_04476_));
 sg13g2_nor2_1 _14840_ (.A(_04468_),
    .B(_04476_),
    .Y(_04478_));
 sg13g2_o21ai_1 _14841_ (.B1(_04477_),
    .Y(_04479_),
    .A1(_04465_),
    .A2(_04478_));
 sg13g2_a21o_1 _14842_ (.A2(_04478_),
    .A1(_04465_),
    .B1(_04479_),
    .X(_04480_));
 sg13g2_o21ai_1 _14843_ (.B1(_04480_),
    .Y(_04481_),
    .A1(_04465_),
    .A2(_04477_));
 sg13g2_xnor2_1 _14844_ (.Y(_04482_),
    .A(_04463_),
    .B(_04481_));
 sg13g2_nand2b_1 _14845_ (.Y(_04483_),
    .B(_04408_),
    .A_N(_04482_));
 sg13g2_nor2b_1 _14846_ (.A(_04408_),
    .B_N(_04482_),
    .Y(_04484_));
 sg13g2_xor2_1 _14847_ (.B(_04482_),
    .A(_04408_),
    .X(_04485_));
 sg13g2_xnor2_1 _14848_ (.Y(_04486_),
    .A(_03816_),
    .B(_03828_));
 sg13g2_xnor2_1 _14849_ (.Y(_04487_),
    .A(_03838_),
    .B(_04486_));
 sg13g2_nor2b_1 _14850_ (.A(_03923_),
    .B_N(_03924_),
    .Y(_04488_));
 sg13g2_xnor2_1 _14851_ (.Y(_04489_),
    .A(_03932_),
    .B(_04488_));
 sg13g2_nand2_1 _14852_ (.Y(_04490_),
    .A(_03949_),
    .B(_03950_));
 sg13g2_xor2_1 _14853_ (.B(_04490_),
    .A(_03956_),
    .X(_04491_));
 sg13g2_nand2b_1 _14854_ (.Y(_04492_),
    .B(_04489_),
    .A_N(_04491_));
 sg13g2_nor2b_1 _14855_ (.A(_04489_),
    .B_N(_04491_),
    .Y(_04493_));
 sg13g2_xnor2_1 _14856_ (.Y(_04494_),
    .A(_04489_),
    .B(_04491_));
 sg13g2_xnor2_1 _14857_ (.Y(_04495_),
    .A(_04487_),
    .B(_04494_));
 sg13g2_xnor2_1 _14858_ (.Y(_04496_),
    .A(_04485_),
    .B(_04495_));
 sg13g2_o21ai_1 _14859_ (.B1(_04039_),
    .Y(_04497_),
    .A1(_04032_),
    .A2(_04038_));
 sg13g2_a21o_1 _14860_ (.A2(_04495_),
    .A1(_04483_),
    .B1(_04484_),
    .X(_04498_));
 sg13g2_a21oi_1 _14861_ (.A1(_04483_),
    .A2(_04495_),
    .Y(_04499_),
    .B1(_04484_));
 sg13g2_a21o_1 _14862_ (.A2(_04497_),
    .A1(_04496_),
    .B1(_04498_),
    .X(_04500_));
 sg13g2_nand3b_1 _14863_ (.B(_04496_),
    .C(_04497_),
    .Y(_04501_),
    .A_N(_04499_));
 sg13g2_nand2_1 _14864_ (.Y(_04502_),
    .A(_04067_),
    .B(_04406_));
 sg13g2_o21ai_1 _14865_ (.B1(_04502_),
    .Y(_04503_),
    .A1(_04319_),
    .A2(_04405_));
 sg13g2_and3_1 _14866_ (.X(_04504_),
    .A(_04500_),
    .B(_04501_),
    .C(_04503_));
 sg13g2_a21oi_1 _14867_ (.A1(_04500_),
    .A2(_04501_),
    .Y(_04505_),
    .B1(_04503_));
 sg13g2_or2_1 _14868_ (.X(_04506_),
    .B(_04404_),
    .A(_04397_));
 sg13g2_a21oi_1 _14869_ (.A1(_04461_),
    .A2(_04481_),
    .Y(_04507_),
    .B1(_04462_));
 sg13g2_a21o_1 _14870_ (.A2(_04506_),
    .A1(_04396_),
    .B1(_04507_),
    .X(_04508_));
 sg13g2_nand3_1 _14871_ (.B(_04506_),
    .C(_04507_),
    .A(_04396_),
    .Y(_04509_));
 sg13g2_nand2_1 _14872_ (.Y(_04510_),
    .A(_04508_),
    .B(_04509_));
 sg13g2_nor2_1 _14873_ (.A(_04250_),
    .B(_04318_),
    .Y(_04511_));
 sg13g2_a21oi_2 _14874_ (.B1(_04511_),
    .Y(_04512_),
    .A2(_04249_),
    .A1(_04154_));
 sg13g2_xnor2_1 _14875_ (.Y(_04513_),
    .A(_04510_),
    .B(_04512_));
 sg13g2_inv_1 _14876_ (.Y(_04514_),
    .A(_04513_));
 sg13g2_o21ai_1 _14877_ (.B1(_04514_),
    .Y(_04515_),
    .A1(_04504_),
    .A2(_04505_));
 sg13g2_inv_1 _14878_ (.Y(_04516_),
    .A(_04515_));
 sg13g2_or3_1 _14879_ (.A(_04504_),
    .B(_04505_),
    .C(_04514_),
    .X(_04517_));
 sg13g2_nor2_1 _14880_ (.A(_03992_),
    .B(_04065_),
    .Y(_04518_));
 sg13g2_nand2_1 _14881_ (.Y(_04519_),
    .A(_04451_),
    .B(_04459_));
 sg13g2_nand2_1 _14882_ (.Y(_04520_),
    .A(_04452_),
    .B(_04519_));
 sg13g2_o21ai_1 _14883_ (.B1(_04520_),
    .Y(_04521_),
    .A1(_04064_),
    .A2(_04518_));
 sg13g2_or3_1 _14884_ (.A(_04064_),
    .B(_04518_),
    .C(_04520_),
    .X(_04522_));
 sg13g2_and2_1 _14885_ (.A(_04521_),
    .B(_04522_),
    .X(_04523_));
 sg13g2_a21oi_2 _14886_ (.B1(_04428_),
    .Y(_04524_),
    .A2(_04435_),
    .A1(_04427_));
 sg13g2_xor2_1 _14887_ (.B(_04524_),
    .A(_04523_),
    .X(_04525_));
 sg13g2_a21o_1 _14888_ (.A2(_04517_),
    .A1(_04515_),
    .B1(_04525_),
    .X(_04526_));
 sg13g2_nand3_1 _14889_ (.B(_04517_),
    .C(_04525_),
    .A(_04515_),
    .Y(_04527_));
 sg13g2_a21oi_1 _14890_ (.A1(_04399_),
    .A2(_04402_),
    .Y(_04528_),
    .B1(_04401_));
 sg13g2_and2_1 _14891_ (.A(_04390_),
    .B(_04394_),
    .X(_04529_));
 sg13g2_o21ai_1 _14892_ (.B1(_04528_),
    .Y(_04530_),
    .A1(_04392_),
    .A2(_04529_));
 sg13g2_nor3_1 _14893_ (.A(_04392_),
    .B(_04528_),
    .C(_04529_),
    .Y(_04531_));
 sg13g2_inv_1 _14894_ (.Y(_04532_),
    .A(_04531_));
 sg13g2_nand2_1 _14895_ (.Y(_04533_),
    .A(_04530_),
    .B(_04532_));
 sg13g2_a21oi_2 _14896_ (.B1(_04120_),
    .Y(_04534_),
    .A2(_04153_),
    .A1(_04121_));
 sg13g2_xnor2_1 _14897_ (.Y(_04535_),
    .A(_04533_),
    .B(_04534_));
 sg13g2_o21ai_1 _14898_ (.B1(_04492_),
    .Y(_04536_),
    .A1(_04487_),
    .A2(_04493_));
 sg13g2_or2_1 _14899_ (.X(_04537_),
    .B(_04536_),
    .A(_04479_));
 sg13g2_inv_1 _14900_ (.Y(_04538_),
    .A(_04537_));
 sg13g2_and2_1 _14901_ (.A(_04479_),
    .B(_04536_),
    .X(_04539_));
 sg13g2_nor2_1 _14902_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sg13g2_xnor2_1 _14903_ (.Y(_04541_),
    .A(_04386_),
    .B(_04540_));
 sg13g2_nand2_1 _14904_ (.Y(_04542_),
    .A(_04535_),
    .B(_04541_));
 sg13g2_xnor2_1 _14905_ (.Y(_04543_),
    .A(_04535_),
    .B(_04541_));
 sg13g2_o21ai_1 _14906_ (.B1(_04305_),
    .Y(_04544_),
    .A1(_04306_),
    .A2(_04317_));
 sg13g2_a21oi_1 _14907_ (.A1(_04246_),
    .A2(_04248_),
    .Y(_04545_),
    .B1(_04544_));
 sg13g2_and3_1 _14908_ (.X(_04546_),
    .A(_04246_),
    .B(_04248_),
    .C(_04544_));
 sg13g2_inv_1 _14909_ (.Y(_04547_),
    .A(_04546_));
 sg13g2_nor2_1 _14910_ (.A(_04545_),
    .B(_04546_),
    .Y(_04548_));
 sg13g2_a21oi_2 _14911_ (.B1(_04011_),
    .Y(_04549_),
    .A2(_04022_),
    .A1(_04012_));
 sg13g2_xor2_1 _14912_ (.B(_04549_),
    .A(_04548_),
    .X(_04550_));
 sg13g2_xnor2_1 _14913_ (.Y(_04551_),
    .A(_04543_),
    .B(_04550_));
 sg13g2_and3_1 _14914_ (.X(_04552_),
    .A(_04526_),
    .B(_04527_),
    .C(_04551_));
 sg13g2_a21oi_1 _14915_ (.A1(_04526_),
    .A2(_04527_),
    .Y(_04553_),
    .B1(_04551_));
 sg13g2_a21o_1 _14916_ (.A2(_04527_),
    .A1(_04526_),
    .B1(_04551_),
    .X(_04554_));
 sg13g2_a21oi_1 _14917_ (.A1(_04262_),
    .A2(_04432_),
    .Y(_04555_),
    .B1(_04433_));
 sg13g2_inv_1 _14918_ (.Y(_04556_),
    .A(_04555_));
 sg13g2_a21oi_1 _14919_ (.A1(_04411_),
    .A2(_04417_),
    .Y(_04557_),
    .B1(_04556_));
 sg13g2_and3_1 _14920_ (.X(_04558_),
    .A(_04411_),
    .B(_04417_),
    .C(_04556_));
 sg13g2_nor2_1 _14921_ (.A(_04557_),
    .B(_04558_),
    .Y(_04559_));
 sg13g2_o21ai_1 _14922_ (.B1(_04475_),
    .Y(_04560_),
    .A1(_04470_),
    .A2(_04471_));
 sg13g2_and2_1 _14923_ (.A(_04472_),
    .B(_04560_),
    .X(_04561_));
 sg13g2_xnor2_1 _14924_ (.Y(_04562_),
    .A(_04559_),
    .B(_04561_));
 sg13g2_nand2_1 _14925_ (.Y(_04563_),
    .A(_04456_),
    .B(_04458_));
 sg13g2_o21ai_1 _14926_ (.B1(_04563_),
    .Y(_04564_),
    .A1(_04454_),
    .A2(_04455_));
 sg13g2_nor2_1 _14927_ (.A(_04443_),
    .B(_04564_),
    .Y(_04565_));
 sg13g2_nand2_1 _14928_ (.Y(_04566_),
    .A(_04443_),
    .B(_04564_));
 sg13g2_nor2b_1 _14929_ (.A(_04565_),
    .B_N(_04566_),
    .Y(_04567_));
 sg13g2_a21oi_1 _14930_ (.A1(_04421_),
    .A2(_04425_),
    .Y(_04568_),
    .B1(_04422_));
 sg13g2_inv_1 _14931_ (.Y(_04569_),
    .A(_04568_));
 sg13g2_xnor2_1 _14932_ (.Y(_04570_),
    .A(_04567_),
    .B(_04569_));
 sg13g2_o21ai_1 _14933_ (.B1(_04447_),
    .Y(_04571_),
    .A1(_04446_),
    .A2(_04449_));
 sg13g2_a21oi_2 _14934_ (.B1(_03989_),
    .Y(_04572_),
    .A2(_03990_),
    .A1(_03971_));
 sg13g2_a21oi_1 _14935_ (.A1(_04051_),
    .A2(_04062_),
    .Y(_04573_),
    .B1(_04053_));
 sg13g2_or2_1 _14936_ (.X(_04574_),
    .B(_04573_),
    .A(_04572_));
 sg13g2_nand2_1 _14937_ (.Y(_04575_),
    .A(_04572_),
    .B(_04573_));
 sg13g2_nand2_1 _14938_ (.Y(_04576_),
    .A(_04574_),
    .B(_04575_));
 sg13g2_xor2_1 _14939_ (.B(_04576_),
    .A(_04571_),
    .X(_04577_));
 sg13g2_nor2_1 _14940_ (.A(_04570_),
    .B(_04577_),
    .Y(_04578_));
 sg13g2_nor3_1 _14941_ (.A(_04562_),
    .B(_04570_),
    .C(_04577_),
    .Y(_04579_));
 sg13g2_a21oi_1 _14942_ (.A1(_04570_),
    .A2(_04577_),
    .Y(_04580_),
    .B1(_04562_));
 sg13g2_nor2_2 _14943_ (.A(_04578_),
    .B(_04580_),
    .Y(_04581_));
 sg13g2_nand3_1 _14944_ (.B(_04570_),
    .C(_04577_),
    .A(_04562_),
    .Y(_04582_));
 sg13g2_a21oi_2 _14945_ (.B1(_04579_),
    .Y(_04583_),
    .A2(_04582_),
    .A1(_04581_));
 sg13g2_o21ai_1 _14946_ (.B1(_04583_),
    .Y(_04584_),
    .A1(_04552_),
    .A2(_04553_));
 sg13g2_or3_1 _14947_ (.A(_04552_),
    .B(_04553_),
    .C(_04583_),
    .X(_04585_));
 sg13g2_and2_1 _14948_ (.A(_04584_),
    .B(_04585_),
    .X(_04586_));
 sg13g2_nand3_1 _14949_ (.B(_04584_),
    .C(_04585_),
    .A(_03962_),
    .Y(_04587_));
 sg13g2_o21ai_1 _14950_ (.B1(_04554_),
    .Y(_04588_),
    .A1(_04552_),
    .A2(_04583_));
 sg13g2_a21oi_1 _14951_ (.A1(_03962_),
    .A2(_04586_),
    .Y(_04589_),
    .B1(_04588_));
 sg13g2_nor2b_1 _14952_ (.A(_04587_),
    .B_N(_04588_),
    .Y(_04590_));
 sg13g2_a21oi_1 _14953_ (.A1(_04517_),
    .A2(_04525_),
    .Y(_04591_),
    .B1(_04516_));
 sg13g2_nor2_1 _14954_ (.A(_04590_),
    .B(_04591_),
    .Y(_04592_));
 sg13g2_o21ai_1 _14955_ (.B1(_04550_),
    .Y(_04593_),
    .A1(_04535_),
    .A2(_04541_));
 sg13g2_nand2_1 _14956_ (.Y(_04594_),
    .A(_04542_),
    .B(_04593_));
 sg13g2_nand2_1 _14957_ (.Y(_04595_),
    .A(_04581_),
    .B(_04594_));
 sg13g2_o21ai_1 _14958_ (.B1(_03960_),
    .Y(_04596_),
    .A1(_04581_),
    .A2(_04594_));
 sg13g2_nand2_1 _14959_ (.Y(_04597_),
    .A(_04595_),
    .B(_04596_));
 sg13g2_o21ai_1 _14960_ (.B1(_04597_),
    .Y(_04598_),
    .A1(_04589_),
    .A2(_04592_));
 sg13g2_nor3_1 _14961_ (.A(_04589_),
    .B(_04592_),
    .C(_04597_),
    .Y(_04599_));
 sg13g2_nand2_1 _14962_ (.Y(_04600_),
    .A(_04500_),
    .B(_04503_));
 sg13g2_and2_1 _14963_ (.A(_04501_),
    .B(_04600_),
    .X(_04601_));
 sg13g2_nand2_1 _14964_ (.Y(_04602_),
    .A(_04509_),
    .B(_04512_));
 sg13g2_nand2_1 _14965_ (.Y(_04603_),
    .A(_04508_),
    .B(_04602_));
 sg13g2_nand2b_1 _14966_ (.Y(_04604_),
    .B(_04601_),
    .A_N(_04603_));
 sg13g2_nor2b_1 _14967_ (.A(_04601_),
    .B_N(_04603_),
    .Y(_04605_));
 sg13g2_nand2_1 _14968_ (.Y(_04606_),
    .A(_04521_),
    .B(_04524_));
 sg13g2_and2_1 _14969_ (.A(_04522_),
    .B(_04606_),
    .X(_04607_));
 sg13g2_a21o_1 _14970_ (.A2(_04607_),
    .A1(_04604_),
    .B1(_04605_),
    .X(_04608_));
 sg13g2_a21oi_2 _14971_ (.B1(_04599_),
    .Y(_04609_),
    .A2(_04608_),
    .A1(_04598_));
 sg13g2_inv_2 _14972_ (.Y(_04610_),
    .A(_04609_));
 sg13g2_nor2_1 _14973_ (.A(_04558_),
    .B(_04561_),
    .Y(_04611_));
 sg13g2_nor2_2 _14974_ (.A(_04557_),
    .B(_04611_),
    .Y(_04612_));
 sg13g2_nand2_1 _14975_ (.Y(_04613_),
    .A(_04571_),
    .B(_04575_));
 sg13g2_o21ai_1 _14976_ (.B1(_04566_),
    .Y(_04614_),
    .A1(_04565_),
    .A2(_04569_));
 sg13g2_nand3_1 _14977_ (.B(_04613_),
    .C(_04614_),
    .A(_04574_),
    .Y(_04615_));
 sg13g2_inv_1 _14978_ (.Y(_04616_),
    .A(_04615_));
 sg13g2_a21oi_1 _14979_ (.A1(_04574_),
    .A2(_04613_),
    .Y(_04617_),
    .B1(_04614_));
 sg13g2_nor2_1 _14980_ (.A(_04616_),
    .B(_04617_),
    .Y(_04618_));
 sg13g2_xor2_1 _14981_ (.B(_04618_),
    .A(_04612_),
    .X(_04619_));
 sg13g2_or2_1 _14982_ (.X(_04620_),
    .B(_04539_),
    .A(_04386_));
 sg13g2_nand2_1 _14983_ (.Y(_04621_),
    .A(_04532_),
    .B(_04534_));
 sg13g2_a22oi_1 _14984_ (.Y(_04622_),
    .B1(_04621_),
    .B2(_04530_),
    .A2(_04620_),
    .A1(_04537_));
 sg13g2_inv_1 _14985_ (.Y(_04623_),
    .A(_04622_));
 sg13g2_and4_1 _14986_ (.A(_04530_),
    .B(_04537_),
    .C(_04620_),
    .D(_04621_),
    .X(_04624_));
 sg13g2_nor2_1 _14987_ (.A(_04622_),
    .B(_04624_),
    .Y(_04625_));
 sg13g2_a21oi_2 _14988_ (.B1(_04545_),
    .Y(_04626_),
    .A2(_04549_),
    .A1(_04547_));
 sg13g2_xor2_1 _14989_ (.B(_04626_),
    .A(_04625_),
    .X(_04627_));
 sg13g2_nor2_1 _14990_ (.A(_04619_),
    .B(_04627_),
    .Y(_04628_));
 sg13g2_xor2_1 _14991_ (.B(_04627_),
    .A(_04619_),
    .X(_04629_));
 sg13g2_a21oi_2 _14992_ (.B1(_03905_),
    .Y(_04630_),
    .A2(_03933_),
    .A1(_03904_));
 sg13g2_xnor2_1 _14993_ (.Y(_04631_),
    .A(_04629_),
    .B(_04630_));
 sg13g2_xor2_1 _14994_ (.B(_04594_),
    .A(_04581_),
    .X(_04632_));
 sg13g2_xnor2_1 _14995_ (.Y(_04633_),
    .A(_03960_),
    .B(_04632_));
 sg13g2_xnor2_1 _14996_ (.Y(_04634_),
    .A(_04587_),
    .B(_04588_));
 sg13g2_xor2_1 _14997_ (.B(_04634_),
    .A(_04591_),
    .X(_04635_));
 sg13g2_nand2_1 _14998_ (.Y(_04636_),
    .A(_04633_),
    .B(_04635_));
 sg13g2_xnor2_1 _14999_ (.Y(_04637_),
    .A(_04601_),
    .B(_04603_));
 sg13g2_xnor2_1 _15000_ (.Y(_04638_),
    .A(_04607_),
    .B(_04637_));
 sg13g2_nor2_1 _15001_ (.A(_04636_),
    .B(_04638_),
    .Y(_04639_));
 sg13g2_nor2_1 _15002_ (.A(_04633_),
    .B(_04635_),
    .Y(_04640_));
 sg13g2_o21ai_1 _15003_ (.B1(_04636_),
    .Y(_04641_),
    .A1(_04638_),
    .A2(_04640_));
 sg13g2_xor2_1 _15004_ (.B(_04635_),
    .A(_04633_),
    .X(_04642_));
 sg13g2_xnor2_1 _15005_ (.Y(_04643_),
    .A(_04638_),
    .B(_04642_));
 sg13g2_and2_1 _15006_ (.A(_04631_),
    .B(_04639_),
    .X(_04644_));
 sg13g2_nand2_1 _15007_ (.Y(_04645_),
    .A(_04631_),
    .B(_04639_));
 sg13g2_a21oi_2 _15008_ (.B1(_04641_),
    .Y(_04646_),
    .A2(_04643_),
    .A1(_04631_));
 sg13g2_nor2_1 _15009_ (.A(_04628_),
    .B(_04630_),
    .Y(_04647_));
 sg13g2_a21oi_2 _15010_ (.B1(_04647_),
    .Y(_04648_),
    .A2(_04627_),
    .A1(_04619_));
 sg13g2_a21oi_2 _15011_ (.B1(_04646_),
    .Y(_04649_),
    .A2(_04648_),
    .A1(_04645_));
 sg13g2_nor2_1 _15012_ (.A(_04598_),
    .B(_04608_),
    .Y(_04650_));
 sg13g2_nand2_1 _15013_ (.Y(_04651_),
    .A(_04599_),
    .B(_04608_));
 sg13g2_o21ai_1 _15014_ (.B1(_04651_),
    .Y(_04652_),
    .A1(_04610_),
    .A2(_04650_));
 sg13g2_o21ai_1 _15015_ (.B1(_04648_),
    .Y(_04653_),
    .A1(_04644_),
    .A2(_04646_));
 sg13g2_or3_1 _15016_ (.A(_04644_),
    .B(_04646_),
    .C(_04648_),
    .X(_04654_));
 sg13g2_a21oi_1 _15017_ (.A1(_04653_),
    .A2(_04654_),
    .Y(_04655_),
    .B1(_04652_));
 sg13g2_and3_1 _15018_ (.X(_04656_),
    .A(_04652_),
    .B(_04653_),
    .C(_04654_));
 sg13g2_nand3_1 _15019_ (.B(_04653_),
    .C(_04654_),
    .A(_04652_),
    .Y(_04657_));
 sg13g2_a21oi_2 _15020_ (.B1(_04624_),
    .Y(_04658_),
    .A2(_04626_),
    .A1(_04623_));
 sg13g2_nor2_1 _15021_ (.A(_04655_),
    .B(_04658_),
    .Y(_04659_));
 sg13g2_nor2_1 _15022_ (.A(_04656_),
    .B(_04659_),
    .Y(_04660_));
 sg13g2_o21ai_1 _15023_ (.B1(_04658_),
    .Y(_04661_),
    .A1(_04655_),
    .A2(_04656_));
 sg13g2_or3_1 _15024_ (.A(_04655_),
    .B(_04656_),
    .C(_04658_),
    .X(_04662_));
 sg13g2_and2_1 _15025_ (.A(_04661_),
    .B(_04662_),
    .X(_04663_));
 sg13g2_a21oi_1 _15026_ (.A1(_04612_),
    .A2(_04615_),
    .Y(_04664_),
    .B1(_04617_));
 sg13g2_inv_1 _15027_ (.Y(_04665_),
    .A(_04664_));
 sg13g2_nand3_1 _15028_ (.B(_04662_),
    .C(_04665_),
    .A(_04661_),
    .Y(_04666_));
 sg13g2_nor3_1 _15029_ (.A(_04657_),
    .B(_04658_),
    .C(_04664_),
    .Y(_04667_));
 sg13g2_xor2_1 _15030_ (.B(_04666_),
    .A(_04660_),
    .X(_04668_));
 sg13g2_xnor2_1 _15031_ (.Y(_04669_),
    .A(_04649_),
    .B(_04668_));
 sg13g2_xor2_1 _15032_ (.B(_04668_),
    .A(_04649_),
    .X(_04670_));
 sg13g2_xnor2_1 _15033_ (.Y(_04671_),
    .A(_04610_),
    .B(_04669_));
 sg13g2_xnor2_1 _15034_ (.Y(_04672_),
    .A(_04609_),
    .B(_04669_));
 sg13g2_nor2_1 _15035_ (.A(_04649_),
    .B(_04667_),
    .Y(_04673_));
 sg13g2_a21oi_1 _15036_ (.A1(_04660_),
    .A2(_04666_),
    .Y(_04674_),
    .B1(_04673_));
 sg13g2_a21oi_2 _15037_ (.B1(_04674_),
    .Y(_04675_),
    .A2(_04670_),
    .A1(_04610_));
 sg13g2_a21o_2 _15038_ (.A2(_04670_),
    .A1(_04610_),
    .B1(_04674_),
    .X(_04676_));
 sg13g2_nor2_1 _15039_ (.A(net2261),
    .B(net2536),
    .Y(_04677_));
 sg13g2_nor2_2 _15040_ (.A(_08421_),
    .B(_04677_),
    .Y(_04678_));
 sg13g2_nor2b_1 _15041_ (.A(net2358),
    .B_N(net2352),
    .Y(_04679_));
 sg13g2_xnor2_1 _15042_ (.Y(_04680_),
    .A(net2358),
    .B(net2350));
 sg13g2_nand2b_1 _15043_ (.Y(_04681_),
    .B(net2424),
    .A_N(net2604));
 sg13g2_o21ai_1 _15044_ (.B1(_04680_),
    .Y(_04682_),
    .A1(net2745),
    .A2(_04681_));
 sg13g2_or3_1 _15045_ (.A(net2745),
    .B(_04680_),
    .C(_04681_),
    .X(_04683_));
 sg13g2_nand2_1 _15046_ (.Y(_04684_),
    .A(_04682_),
    .B(_04683_));
 sg13g2_xor2_1 _15047_ (.B(_04684_),
    .A(_04678_),
    .X(_04685_));
 sg13g2_nor2b_1 _15048_ (.A(net2620),
    .B_N(net2529),
    .Y(_04686_));
 sg13g2_xnor2_1 _15049_ (.Y(_04687_),
    .A(_00001_),
    .B(_04686_));
 sg13g2_xor2_1 _15050_ (.B(net2395),
    .A(net2445),
    .X(_04688_));
 sg13g2_a21o_2 _15051_ (.A2(net2511),
    .A1(_05066_),
    .B1(_04688_),
    .X(_04689_));
 sg13g2_nand2b_1 _15052_ (.Y(_04690_),
    .B(_04687_),
    .A_N(_04689_));
 sg13g2_nor2b_1 _15053_ (.A(_04687_),
    .B_N(_04689_),
    .Y(_04691_));
 sg13g2_xnor2_1 _15054_ (.Y(_04692_),
    .A(_04687_),
    .B(_04689_));
 sg13g2_xnor2_1 _15055_ (.Y(_04693_),
    .A(_02704_),
    .B(_04692_));
 sg13g2_nor2_1 _15056_ (.A(_04685_),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_nand2_1 _15057_ (.Y(_04695_),
    .A(_04685_),
    .B(_04693_));
 sg13g2_nor2_1 _15058_ (.A(net2486),
    .B(net2670),
    .Y(_04696_));
 sg13g2_xnor2_1 _15059_ (.Y(_04697_),
    .A(net2261),
    .B(_04696_));
 sg13g2_xor2_1 _15060_ (.B(net2715),
    .A(net2619),
    .X(_04698_));
 sg13g2_xnor2_1 _15061_ (.Y(_04699_),
    .A(net2419),
    .B(net2401));
 sg13g2_and3_1 _15062_ (.X(_04700_),
    .A(_04697_),
    .B(_04698_),
    .C(_04699_));
 sg13g2_inv_1 _15063_ (.Y(_04701_),
    .A(_04700_));
 sg13g2_xnor2_1 _15064_ (.Y(_04702_),
    .A(net2755),
    .B(net2672));
 sg13g2_a21oi_1 _15065_ (.A1(_04698_),
    .A2(_04699_),
    .Y(_04703_),
    .B1(_04697_));
 sg13g2_a21oi_2 _15066_ (.B1(_04703_),
    .Y(_04704_),
    .A2(_04702_),
    .A1(_04701_));
 sg13g2_nor2_1 _15067_ (.A(_04700_),
    .B(_04703_),
    .Y(_04705_));
 sg13g2_xnor2_1 _15068_ (.Y(_04706_),
    .A(_04702_),
    .B(_04705_));
 sg13g2_o21ai_1 _15069_ (.B1(_04695_),
    .Y(_04707_),
    .A1(_04694_),
    .A2(_04706_));
 sg13g2_xnor2_1 _15070_ (.Y(_04708_),
    .A(net2507),
    .B(net2470));
 sg13g2_xnor2_1 _15071_ (.Y(_04709_),
    .A(net2527),
    .B(net2739));
 sg13g2_nor2_1 _15072_ (.A(_04708_),
    .B(_04709_),
    .Y(_04710_));
 sg13g2_nor2_1 _15073_ (.A(net2428),
    .B(net2223),
    .Y(_04711_));
 sg13g2_nor2_1 _15074_ (.A(_05187_),
    .B(net2250),
    .Y(_04712_));
 sg13g2_xnor2_1 _15075_ (.Y(_04713_),
    .A(_04711_),
    .B(_04712_));
 sg13g2_nand2_1 _15076_ (.Y(_04714_),
    .A(_04708_),
    .B(_04709_));
 sg13g2_nor2b_1 _15077_ (.A(_04710_),
    .B_N(_04714_),
    .Y(_04715_));
 sg13g2_xnor2_1 _15078_ (.Y(_04716_),
    .A(_04713_),
    .B(_04715_));
 sg13g2_a22oi_1 _15079_ (.Y(_04717_),
    .B1(net2619),
    .B2(net2554),
    .A2(net2636),
    .A1(net2631));
 sg13g2_o21ai_1 _15080_ (.B1(_04717_),
    .Y(_04718_),
    .A1(net2554),
    .A2(net2619));
 sg13g2_xor2_1 _15081_ (.B(net2775),
    .A(net2276),
    .X(_04719_));
 sg13g2_xor2_1 _15082_ (.B(net2198),
    .A(net2308),
    .X(_04720_));
 sg13g2_nor2_2 _15083_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sg13g2_nor2_1 _15084_ (.A(net2663),
    .B(net2446),
    .Y(_04722_));
 sg13g2_xnor2_1 _15085_ (.Y(_04723_),
    .A(_02504_),
    .B(_04722_));
 sg13g2_nand2_1 _15086_ (.Y(_04724_),
    .A(_04721_),
    .B(_04723_));
 sg13g2_nor2_1 _15087_ (.A(_04721_),
    .B(_04723_),
    .Y(_04725_));
 sg13g2_inv_1 _15088_ (.Y(_04726_),
    .A(_04725_));
 sg13g2_nand2_1 _15089_ (.Y(_04727_),
    .A(_04724_),
    .B(_04726_));
 sg13g2_xor2_1 _15090_ (.B(_04727_),
    .A(_04718_),
    .X(_04728_));
 sg13g2_nor2_1 _15091_ (.A(_04716_),
    .B(_04728_),
    .Y(_04729_));
 sg13g2_nand2_1 _15092_ (.Y(_04730_),
    .A(_04716_),
    .B(_04728_));
 sg13g2_xor2_1 _15093_ (.B(net2330),
    .A(net2697),
    .X(_04731_));
 sg13g2_nor2_1 _15094_ (.A(net2486),
    .B(net2607),
    .Y(_04732_));
 sg13g2_xnor2_1 _15095_ (.Y(_04733_),
    .A(net2428),
    .B(_04732_));
 sg13g2_nand2b_1 _15096_ (.Y(_04734_),
    .B(net2470),
    .A_N(net2736));
 sg13g2_nor2_1 _15097_ (.A(net2563),
    .B(net2648),
    .Y(_04735_));
 sg13g2_xnor2_1 _15098_ (.Y(_04736_),
    .A(_04734_),
    .B(_04735_));
 sg13g2_nand2_1 _15099_ (.Y(_04737_),
    .A(_04733_),
    .B(_04736_));
 sg13g2_nor2_1 _15100_ (.A(_04733_),
    .B(_04736_),
    .Y(_04738_));
 sg13g2_inv_1 _15101_ (.Y(_04739_),
    .A(_04738_));
 sg13g2_nand2_1 _15102_ (.Y(_04740_),
    .A(_04737_),
    .B(_04739_));
 sg13g2_xnor2_1 _15103_ (.Y(_04741_),
    .A(_04731_),
    .B(_04740_));
 sg13g2_o21ai_1 _15104_ (.B1(_04730_),
    .Y(_04742_),
    .A1(_04729_),
    .A2(_04741_));
 sg13g2_or2_1 _15105_ (.X(_04743_),
    .B(_04742_),
    .A(_04707_));
 sg13g2_inv_1 _15106_ (.Y(_04744_),
    .A(_04743_));
 sg13g2_and2_1 _15107_ (.A(_04707_),
    .B(_04742_),
    .X(_04745_));
 sg13g2_xor2_1 _15108_ (.B(net2504),
    .A(net2563),
    .X(_04746_));
 sg13g2_nor3_2 _15109_ (.A(net2455),
    .B(\net.in[19] ),
    .C(_04746_),
    .Y(_04747_));
 sg13g2_or2_1 _15110_ (.X(_04748_),
    .B(net2648),
    .A(net2257));
 sg13g2_o21ai_1 _15111_ (.B1(_04748_),
    .Y(_04749_),
    .A1(_05561_),
    .A2(net2580));
 sg13g2_xor2_1 _15112_ (.B(net2667),
    .A(net2679),
    .X(_04750_));
 sg13g2_xnor2_1 _15113_ (.Y(_04751_),
    .A(net2616),
    .B(net2749));
 sg13g2_nand2_2 _15114_ (.Y(_04752_),
    .A(_04750_),
    .B(_04751_));
 sg13g2_nand2b_1 _15115_ (.Y(_04753_),
    .B(_04749_),
    .A_N(_04752_));
 sg13g2_nor2b_1 _15116_ (.A(_04749_),
    .B_N(_04752_),
    .Y(_04754_));
 sg13g2_xor2_1 _15117_ (.B(_04752_),
    .A(_04749_),
    .X(_04755_));
 sg13g2_xnor2_1 _15118_ (.Y(_04756_),
    .A(_04747_),
    .B(_04755_));
 sg13g2_xor2_1 _15119_ (.B(net2632),
    .A(net2561),
    .X(_04757_));
 sg13g2_o21ai_1 _15120_ (.B1(_00472_),
    .Y(_04758_),
    .A1(net2670),
    .A2(_04757_));
 sg13g2_xor2_1 _15121_ (.B(\net.in[75] ),
    .A(net2563),
    .X(_04759_));
 sg13g2_or2_1 _15122_ (.X(_04760_),
    .B(_04759_),
    .A(_04758_));
 sg13g2_nand2_1 _15123_ (.Y(_04761_),
    .A(_04758_),
    .B(_04759_));
 sg13g2_xor2_1 _15124_ (.B(_04759_),
    .A(_04758_),
    .X(_04762_));
 sg13g2_xnor2_1 _15125_ (.Y(_04763_),
    .A(_04757_),
    .B(_04762_));
 sg13g2_nor2_1 _15126_ (.A(_04756_),
    .B(_04763_),
    .Y(_04764_));
 sg13g2_nand2_1 _15127_ (.Y(_04765_),
    .A(_04756_),
    .B(_04763_));
 sg13g2_xor2_1 _15128_ (.B(net2396),
    .A(net2401),
    .X(_04766_));
 sg13g2_a21oi_1 _15129_ (.A1(_05605_),
    .A2(_05847_),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_xnor2_1 _15130_ (.Y(_04768_),
    .A(\net.in[108] ),
    .B(\net.in[110] ));
 sg13g2_xnor2_1 _15131_ (.Y(_04769_),
    .A(_02703_),
    .B(_04768_));
 sg13g2_xnor2_1 _15132_ (.Y(_04770_),
    .A(_04767_),
    .B(_04769_));
 sg13g2_o21ai_1 _15133_ (.B1(_04765_),
    .Y(_04771_),
    .A1(_04764_),
    .A2(_04770_));
 sg13g2_nand2b_1 _15134_ (.Y(_04772_),
    .B(_04771_),
    .A_N(_04745_));
 sg13g2_a22oi_1 _15135_ (.Y(_04773_),
    .B1(net2627),
    .B2(net2439),
    .A2(net2225),
    .A1(_05121_));
 sg13g2_nor2_1 _15136_ (.A(net2783),
    .B(net2604),
    .Y(_04774_));
 sg13g2_xnor2_1 _15137_ (.Y(_04775_),
    .A(_00008_),
    .B(_04774_));
 sg13g2_o21ai_1 _15138_ (.B1(_02551_),
    .Y(_04776_),
    .A1(_05363_),
    .A2(net2666));
 sg13g2_nand2_1 _15139_ (.Y(_04777_),
    .A(_04775_),
    .B(_04776_));
 sg13g2_xor2_1 _15140_ (.B(_04776_),
    .A(_04775_),
    .X(_04778_));
 sg13g2_xnor2_1 _15141_ (.Y(_04779_),
    .A(_04773_),
    .B(_04778_));
 sg13g2_xnor2_1 _15142_ (.Y(_04780_),
    .A(net2507),
    .B(net2619));
 sg13g2_nor2b_1 _15143_ (.A(net2313),
    .B_N(net2676),
    .Y(_04781_));
 sg13g2_xnor2_1 _15144_ (.Y(_04782_),
    .A(net2443),
    .B(_04781_));
 sg13g2_nand3b_1 _15145_ (.B(_05253_),
    .C(_02703_),
    .Y(_04783_),
    .A_N(_04782_));
 sg13g2_o21ai_1 _15146_ (.B1(_04782_),
    .Y(_04784_),
    .A1(net2186),
    .A2(_02704_));
 sg13g2_and2_1 _15147_ (.A(_04783_),
    .B(_04784_),
    .X(_04785_));
 sg13g2_xnor2_1 _15148_ (.Y(_04786_),
    .A(_04780_),
    .B(_04785_));
 sg13g2_nand2_1 _15149_ (.Y(_04787_),
    .A(_04779_),
    .B(_04786_));
 sg13g2_xor2_1 _15150_ (.B(net2670),
    .A(net2664),
    .X(_04788_));
 sg13g2_xor2_1 _15151_ (.B(\net.in[161] ),
    .A(net2806),
    .X(_04789_));
 sg13g2_nor2_1 _15152_ (.A(_03930_),
    .B(_04789_),
    .Y(_04790_));
 sg13g2_xnor2_1 _15153_ (.Y(_04791_),
    .A(net2610),
    .B(net2604));
 sg13g2_nor2b_1 _15154_ (.A(_04790_),
    .B_N(_04791_),
    .Y(_04792_));
 sg13g2_nor3_1 _15155_ (.A(_03930_),
    .B(_04789_),
    .C(_04791_),
    .Y(_04793_));
 sg13g2_nor2_1 _15156_ (.A(_04792_),
    .B(_04793_),
    .Y(_04794_));
 sg13g2_nor2_1 _15157_ (.A(_04788_),
    .B(_04793_),
    .Y(_04795_));
 sg13g2_xor2_1 _15158_ (.B(_04794_),
    .A(_04788_),
    .X(_04796_));
 sg13g2_nor2_1 _15159_ (.A(_04779_),
    .B(_04786_),
    .Y(_04797_));
 sg13g2_a21oi_2 _15160_ (.B1(_04797_),
    .Y(_04798_),
    .A2(_04796_),
    .A1(_04787_));
 sg13g2_nor2_1 _15161_ (.A(\net.in[5] ),
    .B(\net.in[34] ),
    .Y(_04799_));
 sg13g2_xnor2_1 _15162_ (.Y(_04800_),
    .A(net2561),
    .B(\net.in[110] ));
 sg13g2_xnor2_1 _15163_ (.Y(_04801_),
    .A(_04799_),
    .B(_04800_));
 sg13g2_nand2b_1 _15164_ (.Y(_04802_),
    .B(net2579),
    .A_N(net2771));
 sg13g2_nand2b_1 _15165_ (.Y(_04803_),
    .B(net2771),
    .A_N(net2578));
 sg13g2_nand2b_1 _15166_ (.Y(_04804_),
    .B(net2806),
    .A_N(net2650));
 sg13g2_nand3_1 _15167_ (.B(_04803_),
    .C(_04804_),
    .A(_04802_),
    .Y(_04805_));
 sg13g2_xor2_1 _15168_ (.B(net2554),
    .A(net2551),
    .X(_04806_));
 sg13g2_nand2_1 _15169_ (.Y(_04807_),
    .A(net2551),
    .B(net2564));
 sg13g2_o21ai_1 _15170_ (.B1(_04807_),
    .Y(_04808_),
    .A1(net2564),
    .A2(_04806_));
 sg13g2_xor2_1 _15171_ (.B(_04808_),
    .A(_04805_),
    .X(_04809_));
 sg13g2_xnor2_1 _15172_ (.Y(_04810_),
    .A(_04801_),
    .B(_04809_));
 sg13g2_inv_1 _15173_ (.Y(_04811_),
    .A(_04810_));
 sg13g2_nor2_2 _15174_ (.A(\net.in[177] ),
    .B(net2250),
    .Y(_04812_));
 sg13g2_nor2_1 _15175_ (.A(net2445),
    .B(net2616),
    .Y(_04813_));
 sg13g2_xnor2_1 _15176_ (.Y(_04814_),
    .A(net2632),
    .B(_04813_));
 sg13g2_xor2_1 _15177_ (.B(net2390),
    .A(net2443),
    .X(_04815_));
 sg13g2_or2_1 _15178_ (.X(_04816_),
    .B(_04815_),
    .A(net2802));
 sg13g2_nor3_1 _15179_ (.A(net2802),
    .B(\net.in[65] ),
    .C(_04815_),
    .Y(_04817_));
 sg13g2_o21ai_1 _15180_ (.B1(_04814_),
    .Y(_04818_),
    .A1(\net.in[65] ),
    .A2(_04816_));
 sg13g2_nor2b_1 _15181_ (.A(_04814_),
    .B_N(_04817_),
    .Y(_04819_));
 sg13g2_xnor2_1 _15182_ (.Y(_04820_),
    .A(_04814_),
    .B(_04817_));
 sg13g2_xnor2_1 _15183_ (.Y(_04821_),
    .A(_04812_),
    .B(_04820_));
 sg13g2_inv_1 _15184_ (.Y(_04822_),
    .A(_04821_));
 sg13g2_nor2_1 _15185_ (.A(net2198),
    .B(\net.in[204] ),
    .Y(_04823_));
 sg13g2_nor2_1 _15186_ (.A(net2302),
    .B(net2744),
    .Y(_04824_));
 sg13g2_xnor2_1 _15187_ (.Y(_04825_),
    .A(_04823_),
    .B(_04824_));
 sg13g2_xor2_1 _15188_ (.B(_01155_),
    .A(net2302),
    .X(_04826_));
 sg13g2_nor2_1 _15189_ (.A(net2561),
    .B(net2616),
    .Y(_04827_));
 sg13g2_nor2_1 _15190_ (.A(net2632),
    .B(net2500),
    .Y(_04828_));
 sg13g2_xor2_1 _15191_ (.B(_04828_),
    .A(_04827_),
    .X(_04829_));
 sg13g2_nor2_1 _15192_ (.A(_04826_),
    .B(_04829_),
    .Y(_04830_));
 sg13g2_xor2_1 _15193_ (.B(_04829_),
    .A(_04826_),
    .X(_04831_));
 sg13g2_a21oi_1 _15194_ (.A1(_04826_),
    .A2(_04829_),
    .Y(_04832_),
    .B1(_04825_));
 sg13g2_nor2_1 _15195_ (.A(_04830_),
    .B(_04832_),
    .Y(_04833_));
 sg13g2_xnor2_1 _15196_ (.Y(_04834_),
    .A(_04825_),
    .B(_04831_));
 sg13g2_o21ai_1 _15197_ (.B1(_04834_),
    .Y(_04835_),
    .A1(_04811_),
    .A2(_04821_));
 sg13g2_o21ai_1 _15198_ (.B1(_04835_),
    .Y(_04836_),
    .A1(_04810_),
    .A2(_04822_));
 sg13g2_xor2_1 _15199_ (.B(net2261),
    .A(\net.in[159] ),
    .X(_04837_));
 sg13g2_nor2_1 _15200_ (.A(net2199),
    .B(_04837_),
    .Y(_04838_));
 sg13g2_inv_2 _15201_ (.Y(_04839_),
    .A(_04838_));
 sg13g2_xnor2_1 _15202_ (.Y(_04840_),
    .A(net2317),
    .B(\net.in[95] ));
 sg13g2_xnor2_1 _15203_ (.Y(_04841_),
    .A(net2777),
    .B(net2706));
 sg13g2_xnor2_1 _15204_ (.Y(_04842_),
    .A(net2771),
    .B(\net.in[79] ));
 sg13g2_a22oi_1 _15205_ (.Y(_04843_),
    .B1(_04842_),
    .B2(_00017_),
    .A2(_04841_),
    .A1(_04840_));
 sg13g2_nand4_1 _15206_ (.B(_04840_),
    .C(_04841_),
    .A(_00017_),
    .Y(_04844_),
    .D(_04842_));
 sg13g2_nor2b_1 _15207_ (.A(_04843_),
    .B_N(_04844_),
    .Y(_04845_));
 sg13g2_a21oi_2 _15208_ (.B1(_04843_),
    .Y(_04846_),
    .A2(_04844_),
    .A1(_04839_));
 sg13g2_xnor2_1 _15209_ (.Y(_04847_),
    .A(_04839_),
    .B(_04845_));
 sg13g2_xor2_1 _15210_ (.B(net2604),
    .A(net2708),
    .X(_04848_));
 sg13g2_xor2_1 _15211_ (.B(net2749),
    .A(net2659),
    .X(_04849_));
 sg13g2_nor2_1 _15212_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sg13g2_o21ai_1 _15213_ (.B1(_00020_),
    .Y(_04851_),
    .A1(net2337),
    .A2(net2632));
 sg13g2_a21oi_2 _15214_ (.B1(_04851_),
    .Y(_04852_),
    .A2(net2632),
    .A1(net2338));
 sg13g2_xnor2_1 _15215_ (.Y(_04853_),
    .A(_02504_),
    .B(_04852_));
 sg13g2_xnor2_1 _15216_ (.Y(_04854_),
    .A(_04850_),
    .B(_04853_));
 sg13g2_xor2_1 _15217_ (.B(net2727),
    .A(net2795),
    .X(_04855_));
 sg13g2_nor2_1 _15218_ (.A(net2266),
    .B(net2199),
    .Y(_04856_));
 sg13g2_xnor2_1 _15219_ (.Y(_04857_),
    .A(net2286),
    .B(_04856_));
 sg13g2_xor2_1 _15220_ (.B(\net.in[74] ),
    .A(net2688),
    .X(_04858_));
 sg13g2_nor2_1 _15221_ (.A(_04857_),
    .B(_04858_),
    .Y(_04859_));
 sg13g2_nand2_1 _15222_ (.Y(_04860_),
    .A(_04857_),
    .B(_04858_));
 sg13g2_nand2b_1 _15223_ (.Y(_04861_),
    .B(_04860_),
    .A_N(_04859_));
 sg13g2_xor2_1 _15224_ (.B(_04861_),
    .A(_04855_),
    .X(_04862_));
 sg13g2_a21o_1 _15225_ (.A2(_04854_),
    .A1(_04847_),
    .B1(_04862_),
    .X(_04863_));
 sg13g2_o21ai_1 _15226_ (.B1(_04863_),
    .Y(_04864_),
    .A1(_04847_),
    .A2(_04854_));
 sg13g2_a21o_1 _15227_ (.A2(_04836_),
    .A1(_04798_),
    .B1(_04864_),
    .X(_04865_));
 sg13g2_o21ai_1 _15228_ (.B1(_04865_),
    .Y(_04866_),
    .A1(_04798_),
    .A2(_04836_));
 sg13g2_nand3_1 _15229_ (.B(_04772_),
    .C(_04866_),
    .A(_04743_),
    .Y(_04867_));
 sg13g2_a21o_2 _15230_ (.A2(_04772_),
    .A1(_04743_),
    .B1(_04866_),
    .X(_04868_));
 sg13g2_nand2_1 _15231_ (.Y(_04869_),
    .A(_04867_),
    .B(_04868_));
 sg13g2_or3_1 _15232_ (.A(net2532),
    .B(net2399),
    .C(_04768_),
    .X(_04870_));
 sg13g2_o21ai_1 _15233_ (.B1(_04768_),
    .Y(_04871_),
    .A1(net2532),
    .A2(net2399));
 sg13g2_nand2_1 _15234_ (.Y(_04872_),
    .A(_04870_),
    .B(_04871_));
 sg13g2_xor2_1 _15235_ (.B(net2514),
    .A(net2358),
    .X(_04873_));
 sg13g2_inv_1 _15236_ (.Y(_04874_),
    .A(_04873_));
 sg13g2_xnor2_1 _15237_ (.Y(_04875_),
    .A(_04872_),
    .B(_04873_));
 sg13g2_nor2b_1 _15238_ (.A(net2396),
    .B_N(net2692),
    .Y(_04876_));
 sg13g2_nor2_1 _15239_ (.A(net2507),
    .B(net2459),
    .Y(_04877_));
 sg13g2_or2_2 _15240_ (.X(_04878_),
    .B(net2363),
    .A(\net.in[13] ));
 sg13g2_o21ai_1 _15241_ (.B1(_04876_),
    .Y(_04879_),
    .A1(_04877_),
    .A2(_04878_));
 sg13g2_inv_1 _15242_ (.Y(_04880_),
    .A(_04879_));
 sg13g2_or3_1 _15243_ (.A(_04876_),
    .B(_04877_),
    .C(_04878_),
    .X(_04881_));
 sg13g2_nand2_1 _15244_ (.Y(_04882_),
    .A(_04879_),
    .B(_04881_));
 sg13g2_nor2_1 _15245_ (.A(net2436),
    .B(net2626),
    .Y(_04883_));
 sg13g2_xor2_1 _15246_ (.B(net2660),
    .A(net2573),
    .X(_04884_));
 sg13g2_xnor2_1 _15247_ (.Y(_04885_),
    .A(_04883_),
    .B(_04884_));
 sg13g2_xor2_1 _15248_ (.B(_04885_),
    .A(_04882_),
    .X(_04886_));
 sg13g2_nand2_1 _15249_ (.Y(_04887_),
    .A(_04875_),
    .B(_04886_));
 sg13g2_or2_1 _15250_ (.X(_04888_),
    .B(_04886_),
    .A(_04875_));
 sg13g2_nor2_1 _15251_ (.A(net2749),
    .B(net2715),
    .Y(_04889_));
 sg13g2_nor2_1 _15252_ (.A(net2616),
    .B(net2784),
    .Y(_04890_));
 sg13g2_xor2_1 _15253_ (.B(_04890_),
    .A(_04889_),
    .X(_04891_));
 sg13g2_nand2b_1 _15254_ (.Y(_04892_),
    .B(net2747),
    .A_N(net2556));
 sg13g2_xnor2_1 _15255_ (.Y(_04893_),
    .A(net2598),
    .B(net2286));
 sg13g2_nand3_1 _15256_ (.B(_04892_),
    .C(_04893_),
    .A(_00563_),
    .Y(_04894_));
 sg13g2_or3_1 _15257_ (.A(net2196),
    .B(net2706),
    .C(_04894_),
    .X(_04895_));
 sg13g2_o21ai_1 _15258_ (.B1(_04894_),
    .Y(_04896_),
    .A1(net2196),
    .A2(net2706));
 sg13g2_nand2_1 _15259_ (.Y(_04897_),
    .A(_04895_),
    .B(_04896_));
 sg13g2_nand2_1 _15260_ (.Y(_04898_),
    .A(_04891_),
    .B(_04895_));
 sg13g2_nand2_2 _15261_ (.Y(_04899_),
    .A(_04896_),
    .B(_04898_));
 sg13g2_xnor2_1 _15262_ (.Y(_04900_),
    .A(_04891_),
    .B(_04897_));
 sg13g2_inv_2 _15263_ (.Y(_04901_),
    .A(_04900_));
 sg13g2_nand2_1 _15264_ (.Y(_04902_),
    .A(_04888_),
    .B(_04901_));
 sg13g2_nor2b_1 _15265_ (.A(net2709),
    .B_N(net2751),
    .Y(_04903_));
 sg13g2_nor2b_1 _15266_ (.A(net2751),
    .B_N(net2709),
    .Y(_04904_));
 sg13g2_nor4_2 _15267_ (.A(net2806),
    .B(\net.in[223] ),
    .C(_04903_),
    .Y(_04905_),
    .D(_04904_));
 sg13g2_nor2_1 _15268_ (.A(net2399),
    .B(net2375),
    .Y(_04906_));
 sg13g2_nor2_1 _15269_ (.A(net2538),
    .B(net2275),
    .Y(_04907_));
 sg13g2_xnor2_1 _15270_ (.Y(_04908_),
    .A(_04906_),
    .B(_04907_));
 sg13g2_a21o_1 _15271_ (.A2(_04905_),
    .A1(_04679_),
    .B1(_04908_),
    .X(_04909_));
 sg13g2_xor2_1 _15272_ (.B(_04905_),
    .A(_04679_),
    .X(_04910_));
 sg13g2_xnor2_1 _15273_ (.Y(_04911_),
    .A(_04908_),
    .B(_04910_));
 sg13g2_xnor2_1 _15274_ (.Y(_04912_),
    .A(net2610),
    .B(net2384));
 sg13g2_xor2_1 _15275_ (.B(net2636),
    .A(net2290),
    .X(_04913_));
 sg13g2_nand2b_1 _15276_ (.Y(_04914_),
    .B(net2574),
    .A_N(net2406));
 sg13g2_xnor2_1 _15277_ (.Y(_04915_),
    .A(net2607),
    .B(net2747));
 sg13g2_xnor2_1 _15278_ (.Y(_04916_),
    .A(_04914_),
    .B(_04915_));
 sg13g2_nand2b_1 _15279_ (.Y(_04917_),
    .B(_04913_),
    .A_N(_04916_));
 sg13g2_nor2b_1 _15280_ (.A(_04913_),
    .B_N(_04916_),
    .Y(_04918_));
 sg13g2_xnor2_1 _15281_ (.Y(_04919_),
    .A(_04913_),
    .B(_04916_));
 sg13g2_xnor2_1 _15282_ (.Y(_04920_),
    .A(_04912_),
    .B(_04919_));
 sg13g2_nand2b_1 _15283_ (.Y(_04921_),
    .B(_04911_),
    .A_N(_04920_));
 sg13g2_nand2b_1 _15284_ (.Y(_04922_),
    .B(_04920_),
    .A_N(_04911_));
 sg13g2_nor2_2 _15285_ (.A(net2440),
    .B(_05693_),
    .Y(_04923_));
 sg13g2_xor2_1 _15286_ (.B(net2803),
    .A(net2653),
    .X(_04924_));
 sg13g2_xor2_1 _15287_ (.B(net2709),
    .A(net2556),
    .X(_04925_));
 sg13g2_nor2_1 _15288_ (.A(_04924_),
    .B(_04925_),
    .Y(_04926_));
 sg13g2_xor2_1 _15289_ (.B(net2747),
    .A(net2659),
    .X(_04927_));
 sg13g2_nor2_2 _15290_ (.A(_02609_),
    .B(_04927_),
    .Y(_04928_));
 sg13g2_nand2_1 _15291_ (.Y(_04929_),
    .A(_04926_),
    .B(_04928_));
 sg13g2_or2_1 _15292_ (.X(_04930_),
    .B(_04928_),
    .A(_04926_));
 sg13g2_nand2_1 _15293_ (.Y(_04931_),
    .A(_04929_),
    .B(_04930_));
 sg13g2_xor2_1 _15294_ (.B(_04931_),
    .A(_04923_),
    .X(_04932_));
 sg13g2_nand2_1 _15295_ (.Y(_04933_),
    .A(_04921_),
    .B(_04932_));
 sg13g2_a22oi_1 _15296_ (.Y(_04934_),
    .B1(_04922_),
    .B2(_04933_),
    .A2(_04902_),
    .A1(_04887_));
 sg13g2_nand4_1 _15297_ (.B(_04902_),
    .C(_04922_),
    .A(_04887_),
    .Y(_04935_),
    .D(_04933_));
 sg13g2_nor2b_1 _15298_ (.A(net2676),
    .B_N(net2765),
    .Y(_04936_));
 sg13g2_xnor2_1 _15299_ (.Y(_04937_),
    .A(net2683),
    .B(_04936_));
 sg13g2_nor2_1 _15300_ (.A(net2366),
    .B(net2288),
    .Y(_04938_));
 sg13g2_xnor2_1 _15301_ (.Y(_04939_),
    .A(net2446),
    .B(net2702));
 sg13g2_xnor2_1 _15302_ (.Y(_04940_),
    .A(_04938_),
    .B(_04939_));
 sg13g2_nor2_1 _15303_ (.A(_04937_),
    .B(_04940_),
    .Y(_04941_));
 sg13g2_xnor2_1 _15304_ (.Y(_04942_),
    .A(_04937_),
    .B(_04940_));
 sg13g2_nor2_1 _15305_ (.A(net2177),
    .B(net2715),
    .Y(_04943_));
 sg13g2_xnor2_1 _15306_ (.Y(_04944_),
    .A(_02505_),
    .B(_04943_));
 sg13g2_xnor2_1 _15307_ (.Y(_04945_),
    .A(_04942_),
    .B(_04944_));
 sg13g2_nand2_1 _15308_ (.Y(_04946_),
    .A(_05033_),
    .B(net2464));
 sg13g2_o21ai_1 _15309_ (.B1(_04946_),
    .Y(_04947_),
    .A1(net2257),
    .A2(net2538));
 sg13g2_nand2b_1 _15310_ (.Y(_04948_),
    .B(net2780),
    .A_N(net2483));
 sg13g2_nand2b_1 _15311_ (.Y(_04949_),
    .B(net2483),
    .A_N(net2780));
 sg13g2_nand2b_1 _15312_ (.Y(_04950_),
    .B(net2808),
    .A_N(net2755));
 sg13g2_nand3_1 _15313_ (.B(_04949_),
    .C(_04950_),
    .A(_04948_),
    .Y(_04951_));
 sg13g2_xnor2_1 _15314_ (.Y(_04952_),
    .A(net2294),
    .B(net2649));
 sg13g2_inv_1 _15315_ (.Y(_04953_),
    .A(_04952_));
 sg13g2_nand2_1 _15316_ (.Y(_04954_),
    .A(_04951_),
    .B(_04953_));
 sg13g2_xnor2_1 _15317_ (.Y(_04955_),
    .A(_04951_),
    .B(_04952_));
 sg13g2_xnor2_1 _15318_ (.Y(_04956_),
    .A(_04947_),
    .B(_04955_));
 sg13g2_inv_1 _15319_ (.Y(_04957_),
    .A(_04956_));
 sg13g2_nand2_1 _15320_ (.Y(_04958_),
    .A(_04945_),
    .B(_04957_));
 sg13g2_nor2_1 _15321_ (.A(_04945_),
    .B(_04957_),
    .Y(_04959_));
 sg13g2_nor2b_1 _15322_ (.A(net2785),
    .B_N(net2459),
    .Y(_04960_));
 sg13g2_a22oi_1 _15323_ (.Y(_04961_),
    .B1(net2783),
    .B2(net2709),
    .A2(_05814_),
    .A1(net2444));
 sg13g2_o21ai_1 _15324_ (.B1(_04961_),
    .Y(_04962_),
    .A1(net2709),
    .A2(net2782));
 sg13g2_xor2_1 _15325_ (.B(net2399),
    .A(net2347),
    .X(_04963_));
 sg13g2_nand2_1 _15326_ (.Y(_04964_),
    .A(_04962_),
    .B(_04963_));
 sg13g2_xor2_1 _15327_ (.B(_04963_),
    .A(_04962_),
    .X(_04965_));
 sg13g2_xnor2_1 _15328_ (.Y(_04966_),
    .A(_04960_),
    .B(_04965_));
 sg13g2_a21oi_2 _15329_ (.B1(_04959_),
    .Y(_04967_),
    .A2(_04966_),
    .A1(_04958_));
 sg13g2_o21ai_1 _15330_ (.B1(_04935_),
    .Y(_04968_),
    .A1(_04934_),
    .A2(_04967_));
 sg13g2_xnor2_1 _15331_ (.Y(_04969_),
    .A(_04869_),
    .B(_04968_));
 sg13g2_nand2_1 _15332_ (.Y(_04970_),
    .A(_04887_),
    .B(_04888_));
 sg13g2_xnor2_1 _15333_ (.Y(_04971_),
    .A(_04901_),
    .B(_04970_));
 sg13g2_xor2_1 _15334_ (.B(_04763_),
    .A(_04756_),
    .X(_04972_));
 sg13g2_xnor2_1 _15335_ (.Y(_04973_),
    .A(_04770_),
    .B(_04972_));
 sg13g2_xnor2_1 _15336_ (.Y(_04974_),
    .A(_04911_),
    .B(_04920_));
 sg13g2_xnor2_1 _15337_ (.Y(_04975_),
    .A(_04932_),
    .B(_04974_));
 sg13g2_nand2_1 _15338_ (.Y(_04976_),
    .A(_04973_),
    .B(_04975_));
 sg13g2_or2_1 _15339_ (.X(_04977_),
    .B(_04975_),
    .A(_04973_));
 sg13g2_xor2_1 _15340_ (.B(_04975_),
    .A(_04973_),
    .X(_04978_));
 sg13g2_xnor2_1 _15341_ (.Y(_04979_),
    .A(_04971_),
    .B(_04978_));
 sg13g2_inv_1 _15342_ (.Y(_04980_),
    .A(_04979_));
 sg13g2_a21oi_1 _15343_ (.A1(_05341_),
    .A2(net2659),
    .Y(_04981_),
    .B1(net2747));
 sg13g2_a21oi_1 _15344_ (.A1(net2497),
    .A2(_05836_),
    .Y(_04982_),
    .B1(net2775));
 sg13g2_nand2_2 _15345_ (.Y(_04983_),
    .A(_04981_),
    .B(_04982_));
 sg13g2_xnor2_1 _15346_ (.Y(_04984_),
    .A(_04945_),
    .B(_04956_));
 sg13g2_xnor2_1 _15347_ (.Y(_04985_),
    .A(_04966_),
    .B(_04984_));
 sg13g2_nor2_2 _15348_ (.A(net2219),
    .B(net2314),
    .Y(_04986_));
 sg13g2_nor2b_1 _15349_ (.A(net2532),
    .B_N(net2610),
    .Y(_04987_));
 sg13g2_o21ai_1 _15350_ (.B1(_04806_),
    .Y(_04988_),
    .A1(_04986_),
    .A2(_04987_));
 sg13g2_nor3_1 _15351_ (.A(_04806_),
    .B(_04986_),
    .C(_04987_),
    .Y(_04989_));
 sg13g2_or3_1 _15352_ (.A(_04806_),
    .B(_04986_),
    .C(_04987_),
    .X(_04990_));
 sg13g2_and2_1 _15353_ (.A(_04988_),
    .B(_04990_),
    .X(_04991_));
 sg13g2_nor2_1 _15354_ (.A(net2440),
    .B(net2233),
    .Y(_04992_));
 sg13g2_nor2_1 _15355_ (.A(net2308),
    .B(net2355),
    .Y(_04993_));
 sg13g2_xor2_1 _15356_ (.B(_04993_),
    .A(_04992_),
    .X(_04994_));
 sg13g2_xnor2_1 _15357_ (.Y(_04995_),
    .A(_04991_),
    .B(_04994_));
 sg13g2_nand2b_1 _15358_ (.Y(_04996_),
    .B(net2617),
    .A_N(net2605));
 sg13g2_o21ai_1 _15359_ (.B1(_04996_),
    .Y(_04997_),
    .A1(_05462_),
    .A2(\net.in[229] ));
 sg13g2_a21oi_2 _15360_ (.B1(_04997_),
    .Y(_04998_),
    .A2(net2604),
    .A1(_05770_));
 sg13g2_xnor2_1 _15361_ (.Y(_04999_),
    .A(net2753),
    .B(net2670));
 sg13g2_a21oi_2 _15362_ (.B1(_04999_),
    .Y(_05001_),
    .A2(_05495_),
    .A1(net2184));
 sg13g2_nor2_1 _15363_ (.A(net2664),
    .B(net2464),
    .Y(_05002_));
 sg13g2_nor2_1 _15364_ (.A(net2498),
    .B(net2504),
    .Y(_05003_));
 sg13g2_xnor2_1 _15365_ (.Y(_05004_),
    .A(_05002_),
    .B(_05003_));
 sg13g2_nand2b_1 _15366_ (.Y(_05005_),
    .B(_05004_),
    .A_N(_05001_));
 sg13g2_nor2b_1 _15367_ (.A(_05004_),
    .B_N(_05001_),
    .Y(_05006_));
 sg13g2_xnor2_1 _15368_ (.Y(_05007_),
    .A(_05001_),
    .B(_05004_));
 sg13g2_xor2_1 _15369_ (.B(_05007_),
    .A(_04998_),
    .X(_05008_));
 sg13g2_xnor2_1 _15370_ (.Y(_05009_),
    .A(_04998_),
    .B(_05007_));
 sg13g2_nand2b_1 _15371_ (.Y(_05010_),
    .B(_05008_),
    .A_N(_04995_));
 sg13g2_xnor2_1 _15372_ (.Y(_05012_),
    .A(_04995_),
    .B(_05008_));
 sg13g2_nand2_1 _15373_ (.Y(_05013_),
    .A(net2679),
    .B(net2620));
 sg13g2_nor2_1 _15374_ (.A(net2679),
    .B(net2619),
    .Y(_05014_));
 sg13g2_o21ai_1 _15375_ (.B1(_05013_),
    .Y(_05015_),
    .A1(\net.in[139] ),
    .A2(_05561_));
 sg13g2_xor2_1 _15376_ (.B(net2667),
    .A(net2751),
    .X(_05016_));
 sg13g2_xnor2_1 _15377_ (.Y(_05017_),
    .A(_00485_),
    .B(_05016_));
 sg13g2_o21ai_1 _15378_ (.B1(_05017_),
    .Y(_05018_),
    .A1(_05014_),
    .A2(_05015_));
 sg13g2_nor3_1 _15379_ (.A(_05014_),
    .B(_05015_),
    .C(_05017_),
    .Y(_05019_));
 sg13g2_or3_1 _15380_ (.A(_05014_),
    .B(_05015_),
    .C(_05017_),
    .X(_05020_));
 sg13g2_nand2_1 _15381_ (.Y(_05021_),
    .A(_05018_),
    .B(_05020_));
 sg13g2_xnor2_1 _15382_ (.Y(_05023_),
    .A(net2636),
    .B(_02849_));
 sg13g2_xnor2_1 _15383_ (.Y(_05024_),
    .A(_05021_),
    .B(_05023_));
 sg13g2_xnor2_1 _15384_ (.Y(_05025_),
    .A(_05012_),
    .B(_05024_));
 sg13g2_nor2b_1 _15385_ (.A(_04985_),
    .B_N(_05025_),
    .Y(_05026_));
 sg13g2_nand2b_1 _15386_ (.Y(_05027_),
    .B(_04985_),
    .A_N(_05025_));
 sg13g2_xnor2_1 _15387_ (.Y(_05028_),
    .A(_04985_),
    .B(_05025_));
 sg13g2_a21o_1 _15388_ (.A2(_05027_),
    .A1(_04983_),
    .B1(_05026_),
    .X(_05029_));
 sg13g2_xnor2_1 _15389_ (.Y(_05030_),
    .A(_04983_),
    .B(_05028_));
 sg13g2_nor2_1 _15390_ (.A(_04980_),
    .B(_05030_),
    .Y(_05031_));
 sg13g2_nor2_1 _15391_ (.A(\net.in[10] ),
    .B(net2644),
    .Y(_05032_));
 sg13g2_xnor2_1 _15392_ (.Y(_05034_),
    .A(net2286),
    .B(_05032_));
 sg13g2_xor2_1 _15393_ (.B(net2568),
    .A(net2346),
    .X(_05035_));
 sg13g2_xnor2_1 _15394_ (.Y(_05036_),
    .A(net2636),
    .B(net2620));
 sg13g2_inv_1 _15395_ (.Y(_05037_),
    .A(_05036_));
 sg13g2_nand2b_1 _15396_ (.Y(_05038_),
    .B(_05036_),
    .A_N(_05035_));
 sg13g2_xnor2_1 _15397_ (.Y(_05039_),
    .A(_05035_),
    .B(_05036_));
 sg13g2_xnor2_1 _15398_ (.Y(_05040_),
    .A(_05034_),
    .B(_05039_));
 sg13g2_nor2b_1 _15399_ (.A(net2610),
    .B_N(net2723),
    .Y(_05041_));
 sg13g2_xor2_1 _15400_ (.B(net2604),
    .A(net2810),
    .X(_05042_));
 sg13g2_xnor2_1 _15401_ (.Y(_05043_),
    .A(_05041_),
    .B(_05042_));
 sg13g2_or2_1 _15402_ (.X(_05045_),
    .B(net2627),
    .A(net2719));
 sg13g2_a21oi_1 _15403_ (.A1(net2718),
    .A2(net2626),
    .Y(_05046_),
    .B1(net2456));
 sg13g2_nand2b_1 _15404_ (.Y(_05047_),
    .B(net2436),
    .A_N(net2487));
 sg13g2_and4_2 _15405_ (.A(_02814_),
    .B(_05045_),
    .C(_05046_),
    .D(_05047_),
    .X(_05048_));
 sg13g2_inv_1 _15406_ (.Y(_05049_),
    .A(_05048_));
 sg13g2_a22oi_1 _15407_ (.Y(_05050_),
    .B1(_05047_),
    .B2(_02814_),
    .A2(_05046_),
    .A1(_05045_));
 sg13g2_or3_1 _15408_ (.A(_05043_),
    .B(_05048_),
    .C(_05050_),
    .X(_05051_));
 sg13g2_o21ai_1 _15409_ (.B1(_05043_),
    .Y(_05052_),
    .A1(_05048_),
    .A2(_05050_));
 sg13g2_o21ai_1 _15410_ (.B1(_05049_),
    .Y(_05053_),
    .A1(_05043_),
    .A2(_05050_));
 sg13g2_and3_1 _15411_ (.X(_05054_),
    .A(_05040_),
    .B(_05051_),
    .C(_05052_));
 sg13g2_a21oi_1 _15412_ (.A1(_05051_),
    .A2(_05052_),
    .Y(_05056_),
    .B1(_05040_));
 sg13g2_nor2_1 _15413_ (.A(_05054_),
    .B(_05056_),
    .Y(_05057_));
 sg13g2_nand2_1 _15414_ (.Y(_05058_),
    .A(net2560),
    .B(net2179));
 sg13g2_xnor2_1 _15415_ (.Y(_05059_),
    .A(\net.in[209] ),
    .B(net2745));
 sg13g2_xnor2_1 _15416_ (.Y(_05060_),
    .A(_05058_),
    .B(_05059_));
 sg13g2_nor2_1 _15417_ (.A(net2594),
    .B(net2745),
    .Y(_05061_));
 sg13g2_xnor2_1 _15418_ (.Y(_05062_),
    .A(net2446),
    .B(_05061_));
 sg13g2_inv_1 _15419_ (.Y(_05063_),
    .A(_05062_));
 sg13g2_nor2b_1 _15420_ (.A(net2659),
    .B_N(net2205),
    .Y(_05064_));
 sg13g2_nor2_1 _15421_ (.A(_05836_),
    .B(net2205),
    .Y(_05065_));
 sg13g2_nor4_2 _15422_ (.A(net2745),
    .B(net2314),
    .C(_05064_),
    .Y(_05067_),
    .D(_05065_));
 sg13g2_nand2_1 _15423_ (.Y(_05068_),
    .A(_05063_),
    .B(_05067_));
 sg13g2_xnor2_1 _15424_ (.Y(_05069_),
    .A(_05062_),
    .B(_05067_));
 sg13g2_o21ai_1 _15425_ (.B1(_05060_),
    .Y(_05070_),
    .A1(_05063_),
    .A2(_05067_));
 sg13g2_and2_1 _15426_ (.A(_05068_),
    .B(_05070_),
    .X(_05071_));
 sg13g2_xnor2_1 _15427_ (.Y(_05072_),
    .A(_05060_),
    .B(_05069_));
 sg13g2_nor2b_1 _15428_ (.A(_05056_),
    .B_N(_05072_),
    .Y(_05073_));
 sg13g2_xnor2_1 _15429_ (.Y(_05074_),
    .A(_05057_),
    .B(_05072_));
 sg13g2_xnor2_1 _15430_ (.Y(_05075_),
    .A(net2626),
    .B(net2640));
 sg13g2_nor3_2 _15431_ (.A(net2610),
    .B(net2709),
    .C(_05075_),
    .Y(_05076_));
 sg13g2_xnor2_1 _15432_ (.Y(_05078_),
    .A(net2672),
    .B(net2784));
 sg13g2_nor2_1 _15433_ (.A(net2524),
    .B(net2780),
    .Y(_05079_));
 sg13g2_nor2_1 _15434_ (.A(net2514),
    .B(net2775),
    .Y(_05080_));
 sg13g2_xnor2_1 _15435_ (.Y(_05081_),
    .A(_05079_),
    .B(_05080_));
 sg13g2_nand2b_1 _15436_ (.Y(_05082_),
    .B(_05081_),
    .A_N(_05078_));
 sg13g2_nor2b_1 _15437_ (.A(_05081_),
    .B_N(_05078_),
    .Y(_05083_));
 sg13g2_o21ai_1 _15438_ (.B1(_05082_),
    .Y(_05084_),
    .A1(_05076_),
    .A2(_05083_));
 sg13g2_xor2_1 _15439_ (.B(_05081_),
    .A(_05078_),
    .X(_05085_));
 sg13g2_xnor2_1 _15440_ (.Y(_05086_),
    .A(_05076_),
    .B(_05085_));
 sg13g2_nor2_1 _15441_ (.A(net2676),
    .B(net2683),
    .Y(_05087_));
 sg13g2_xor2_1 _15442_ (.B(net2607),
    .A(net2712),
    .X(_05089_));
 sg13g2_xnor2_1 _15443_ (.Y(_05090_),
    .A(_05087_),
    .B(_05089_));
 sg13g2_xor2_1 _15444_ (.B(net2511),
    .A(net2414),
    .X(_05091_));
 sg13g2_nor2b_1 _15445_ (.A(net2712),
    .B_N(net2791),
    .Y(_05092_));
 sg13g2_nor2b_1 _15446_ (.A(net2617),
    .B_N(net2718),
    .Y(_05093_));
 sg13g2_xnor2_1 _15447_ (.Y(_05094_),
    .A(_05092_),
    .B(_05093_));
 sg13g2_a21o_1 _15448_ (.A2(_05094_),
    .A1(_05091_),
    .B1(_05090_),
    .X(_05095_));
 sg13g2_o21ai_1 _15449_ (.B1(_05095_),
    .Y(_05096_),
    .A1(_05091_),
    .A2(_05094_));
 sg13g2_xnor2_1 _15450_ (.Y(_05097_),
    .A(_05091_),
    .B(_05094_));
 sg13g2_xnor2_1 _15451_ (.Y(_05098_),
    .A(_05090_),
    .B(_05097_));
 sg13g2_nor2_1 _15452_ (.A(_05086_),
    .B(_05098_),
    .Y(_05100_));
 sg13g2_xnor2_1 _15453_ (.Y(_05101_),
    .A(net2514),
    .B(net2446));
 sg13g2_xnor2_1 _15454_ (.Y(_05102_),
    .A(net2323),
    .B(net2464));
 sg13g2_xor2_1 _15455_ (.B(_05102_),
    .A(_00018_),
    .X(_05103_));
 sg13g2_xnor2_1 _15456_ (.Y(_05104_),
    .A(_05101_),
    .B(_05103_));
 sg13g2_a21oi_1 _15457_ (.A1(_05086_),
    .A2(_05098_),
    .Y(_05105_),
    .B1(_05104_));
 sg13g2_xnor2_1 _15458_ (.Y(_05106_),
    .A(_05086_),
    .B(_05098_));
 sg13g2_xnor2_1 _15459_ (.Y(_05107_),
    .A(_05104_),
    .B(_05106_));
 sg13g2_or2_1 _15460_ (.X(_05108_),
    .B(_05107_),
    .A(_05074_));
 sg13g2_nand2_1 _15461_ (.Y(_05109_),
    .A(_05074_),
    .B(_05107_));
 sg13g2_xor2_1 _15462_ (.B(_05107_),
    .A(_05074_),
    .X(_05111_));
 sg13g2_xnor2_1 _15463_ (.Y(_05112_),
    .A(net2507),
    .B(net2424));
 sg13g2_xnor2_1 _15464_ (.Y(_05113_),
    .A(net2196),
    .B(net2659));
 sg13g2_xnor2_1 _15465_ (.Y(_05114_),
    .A(_04924_),
    .B(_05113_));
 sg13g2_nor2_1 _15466_ (.A(net2307),
    .B(net2225),
    .Y(_05115_));
 sg13g2_xnor2_1 _15467_ (.Y(_05116_),
    .A(_04815_),
    .B(_05115_));
 sg13g2_nor2_1 _15468_ (.A(_05114_),
    .B(_05116_),
    .Y(_05117_));
 sg13g2_nand2_1 _15469_ (.Y(_05118_),
    .A(_05114_),
    .B(_05116_));
 sg13g2_xnor2_1 _15470_ (.Y(_05119_),
    .A(_05114_),
    .B(_05116_));
 sg13g2_xnor2_1 _15471_ (.Y(_05120_),
    .A(_05112_),
    .B(_05119_));
 sg13g2_a21oi_2 _15472_ (.B1(net2808),
    .Y(_05122_),
    .A2(net2639),
    .A1(_05110_));
 sg13g2_a21oi_1 _15473_ (.A1(net2241),
    .A2(_05979_),
    .Y(_05123_),
    .B1(net2706));
 sg13g2_nand2_2 _15474_ (.Y(_05124_),
    .A(_05122_),
    .B(_05123_));
 sg13g2_xnor2_1 _15475_ (.Y(_05125_),
    .A(net2290),
    .B(net2736));
 sg13g2_nor2_1 _15476_ (.A(net2556),
    .B(net2500),
    .Y(_05126_));
 sg13g2_nor2_1 _15477_ (.A(net2551),
    .B(net2406),
    .Y(_05127_));
 sg13g2_xor2_1 _15478_ (.B(_05127_),
    .A(_05126_),
    .X(_05128_));
 sg13g2_nor2_1 _15479_ (.A(_05125_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_nand2_1 _15480_ (.Y(_05130_),
    .A(_05125_),
    .B(_05128_));
 sg13g2_xor2_1 _15481_ (.B(_05128_),
    .A(_05125_),
    .X(_05131_));
 sg13g2_a21oi_2 _15482_ (.B1(_05129_),
    .Y(_05133_),
    .A2(_05130_),
    .A1(_05124_));
 sg13g2_xnor2_1 _15483_ (.Y(_05134_),
    .A(_05124_),
    .B(_05131_));
 sg13g2_nor2_1 _15484_ (.A(_05120_),
    .B(_05134_),
    .Y(_05135_));
 sg13g2_nand2_1 _15485_ (.Y(_05136_),
    .A(_05120_),
    .B(_05134_));
 sg13g2_nand2b_1 _15486_ (.Y(_05137_),
    .B(_05136_),
    .A_N(_05135_));
 sg13g2_nor2_1 _15487_ (.A(net2607),
    .B(\net.in[28] ),
    .Y(_05138_));
 sg13g2_xnor2_1 _15488_ (.Y(_05139_),
    .A(net2708),
    .B(\net.in[191] ));
 sg13g2_xnor2_1 _15489_ (.Y(_05140_),
    .A(_05138_),
    .B(_05139_));
 sg13g2_xnor2_1 _15490_ (.Y(_05141_),
    .A(net2440),
    .B(net2616));
 sg13g2_and2_1 _15491_ (.A(net2663),
    .B(net2626),
    .X(_05142_));
 sg13g2_nor2_1 _15492_ (.A(net2664),
    .B(_02504_),
    .Y(_05144_));
 sg13g2_nor3_1 _15493_ (.A(_05141_),
    .B(_05142_),
    .C(_05144_),
    .Y(_05145_));
 sg13g2_o21ai_1 _15494_ (.B1(_05141_),
    .Y(_05146_),
    .A1(_05142_),
    .A2(_05144_));
 sg13g2_a21oi_2 _15495_ (.B1(_05145_),
    .Y(_05147_),
    .A2(_05146_),
    .A1(_05140_));
 sg13g2_or2_1 _15496_ (.X(_05148_),
    .B(_05146_),
    .A(_05140_));
 sg13g2_a22oi_1 _15497_ (.Y(_05149_),
    .B1(_05147_),
    .B2(_05148_),
    .A2(_05145_),
    .A1(_05140_));
 sg13g2_xnor2_1 _15498_ (.Y(_05150_),
    .A(_05137_),
    .B(_05149_));
 sg13g2_xnor2_1 _15499_ (.Y(_05151_),
    .A(_05111_),
    .B(_05150_));
 sg13g2_xnor2_1 _15500_ (.Y(_05152_),
    .A(net2653),
    .B(net2749));
 sg13g2_xor2_1 _15501_ (.B(net2806),
    .A(net2664),
    .X(_05153_));
 sg13g2_xnor2_1 _15502_ (.Y(_05155_),
    .A(_05152_),
    .B(_05153_));
 sg13g2_o21ai_1 _15503_ (.B1(_02834_),
    .Y(_05156_),
    .A1(net2507),
    .A2(_05836_));
 sg13g2_nand2_2 _15504_ (.Y(_05157_),
    .A(_00021_),
    .B(_02536_));
 sg13g2_nor2b_1 _15505_ (.A(_05157_),
    .B_N(_05156_),
    .Y(_05158_));
 sg13g2_nand2b_1 _15506_ (.Y(_05159_),
    .B(_05157_),
    .A_N(_05156_));
 sg13g2_xor2_1 _15507_ (.B(_05157_),
    .A(_05156_),
    .X(_05160_));
 sg13g2_xnor2_1 _15508_ (.Y(_05161_),
    .A(_05155_),
    .B(_05160_));
 sg13g2_nor2_1 _15509_ (.A(net2723),
    .B(net2709),
    .Y(_05162_));
 sg13g2_xnor2_1 _15510_ (.Y(_05163_),
    .A(net2712),
    .B(_05162_));
 sg13g2_nand2_1 _15511_ (.Y(_05164_),
    .A(net2733),
    .B(net2644));
 sg13g2_xor2_1 _15512_ (.B(_05164_),
    .A(net2240),
    .X(_05166_));
 sg13g2_xnor2_1 _15513_ (.Y(_05167_),
    .A(net2753),
    .B(net2672));
 sg13g2_a21oi_2 _15514_ (.B1(_05167_),
    .Y(_05168_),
    .A2(_05693_),
    .A1(_05594_));
 sg13g2_nor2b_1 _15515_ (.A(_05168_),
    .B_N(_05166_),
    .Y(_05169_));
 sg13g2_nor2b_1 _15516_ (.A(_05166_),
    .B_N(_05168_),
    .Y(_05170_));
 sg13g2_xnor2_1 _15517_ (.Y(_05171_),
    .A(_05166_),
    .B(_05168_));
 sg13g2_xnor2_1 _15518_ (.Y(_05172_),
    .A(_05163_),
    .B(_05171_));
 sg13g2_nand2_1 _15519_ (.Y(_05173_),
    .A(_05161_),
    .B(_05172_));
 sg13g2_xnor2_1 _15520_ (.Y(_05174_),
    .A(_05161_),
    .B(_05172_));
 sg13g2_and2_1 _15521_ (.A(net2679),
    .B(net2672),
    .X(_05175_));
 sg13g2_xor2_1 _15522_ (.B(net2774),
    .A(net2708),
    .X(_05177_));
 sg13g2_nor3_2 _15523_ (.A(_02773_),
    .B(_05175_),
    .C(_05177_),
    .Y(_05178_));
 sg13g2_xnor2_1 _15524_ (.Y(_05179_),
    .A(net2439),
    .B(_00007_));
 sg13g2_xnor2_1 _15525_ (.Y(_05180_),
    .A(net2350),
    .B(_05179_));
 sg13g2_or2_1 _15526_ (.X(_05181_),
    .B(net2254),
    .A(net2191));
 sg13g2_o21ai_1 _15527_ (.B1(_05181_),
    .Y(_05182_),
    .A1(net2659),
    .A2(net2727));
 sg13g2_nand2_2 _15528_ (.Y(_05183_),
    .A(_05180_),
    .B(_05182_));
 sg13g2_xor2_1 _15529_ (.B(_05182_),
    .A(_05180_),
    .X(_05184_));
 sg13g2_xnor2_1 _15530_ (.Y(_05185_),
    .A(_05178_),
    .B(_05184_));
 sg13g2_o21ai_1 _15531_ (.B1(_05185_),
    .Y(_05186_),
    .A1(_05161_),
    .A2(_05172_));
 sg13g2_xnor2_1 _15532_ (.Y(_05188_),
    .A(_05174_),
    .B(_05185_));
 sg13g2_xnor2_1 _15533_ (.Y(_05189_),
    .A(_04810_),
    .B(_04821_));
 sg13g2_xnor2_1 _15534_ (.Y(_05190_),
    .A(_04834_),
    .B(_05189_));
 sg13g2_nand2b_1 _15535_ (.Y(_05191_),
    .B(_05190_),
    .A_N(_05188_));
 sg13g2_nand2b_1 _15536_ (.Y(_05192_),
    .B(_05188_),
    .A_N(_05190_));
 sg13g2_xnor2_1 _15537_ (.Y(_05193_),
    .A(_05188_),
    .B(_05190_));
 sg13g2_xnor2_1 _15538_ (.Y(_05194_),
    .A(_04779_),
    .B(_04786_));
 sg13g2_xnor2_1 _15539_ (.Y(_05195_),
    .A(_04796_),
    .B(_05194_));
 sg13g2_xnor2_1 _15540_ (.Y(_05196_),
    .A(_05193_),
    .B(_05195_));
 sg13g2_nand2b_1 _15541_ (.Y(_05197_),
    .B(_05196_),
    .A_N(_05151_));
 sg13g2_nor2b_1 _15542_ (.A(_05196_),
    .B_N(_05151_),
    .Y(_05199_));
 sg13g2_xor2_1 _15543_ (.B(_04854_),
    .A(_04847_),
    .X(_05200_));
 sg13g2_xnor2_1 _15544_ (.Y(_05201_),
    .A(_04862_),
    .B(_05200_));
 sg13g2_xnor2_1 _15545_ (.Y(_05202_),
    .A(_04685_),
    .B(_04693_));
 sg13g2_xnor2_1 _15546_ (.Y(_05203_),
    .A(_04706_),
    .B(_05202_));
 sg13g2_nor2_1 _15547_ (.A(_05201_),
    .B(_05203_),
    .Y(_05204_));
 sg13g2_nand2_1 _15548_ (.Y(_05205_),
    .A(_05201_),
    .B(_05203_));
 sg13g2_nand2b_1 _15549_ (.Y(_05206_),
    .B(_05205_),
    .A_N(_05204_));
 sg13g2_xor2_1 _15550_ (.B(_04728_),
    .A(_04716_),
    .X(_05207_));
 sg13g2_xnor2_1 _15551_ (.Y(_05208_),
    .A(_04741_),
    .B(_05207_));
 sg13g2_xnor2_1 _15552_ (.Y(_05210_),
    .A(_05206_),
    .B(_05208_));
 sg13g2_a21o_1 _15553_ (.A2(_05210_),
    .A1(_05197_),
    .B1(_05199_),
    .X(_05211_));
 sg13g2_xor2_1 _15554_ (.B(_05030_),
    .A(_04979_),
    .X(_05212_));
 sg13g2_xor2_1 _15555_ (.B(_05196_),
    .A(_05151_),
    .X(_05213_));
 sg13g2_xnor2_1 _15556_ (.Y(_05214_),
    .A(_05210_),
    .B(_05213_));
 sg13g2_nor4_1 _15557_ (.A(_05197_),
    .B(_05199_),
    .C(_05210_),
    .D(_05212_),
    .Y(_05215_));
 sg13g2_nor2_1 _15558_ (.A(_05031_),
    .B(_05215_),
    .Y(_05216_));
 sg13g2_o21ai_1 _15559_ (.B1(_05211_),
    .Y(_05217_),
    .A1(_05212_),
    .A2(_05214_));
 sg13g2_nand2b_1 _15560_ (.Y(_05218_),
    .B(_05217_),
    .A_N(_05216_));
 sg13g2_o21ai_1 _15561_ (.B1(_04881_),
    .Y(_05219_),
    .A1(_04880_),
    .A2(_04885_));
 sg13g2_nand2_1 _15562_ (.Y(_05221_),
    .A(_04923_),
    .B(_04929_));
 sg13g2_nand2_1 _15563_ (.Y(_05222_),
    .A(_04870_),
    .B(_04874_));
 sg13g2_and4_1 _15564_ (.A(_04871_),
    .B(_04930_),
    .C(_05221_),
    .D(_05222_),
    .X(_05223_));
 sg13g2_a22oi_1 _15565_ (.Y(_05224_),
    .B1(_05222_),
    .B2(_04871_),
    .A2(_05221_),
    .A1(_04930_));
 sg13g2_nand2b_1 _15566_ (.Y(_05225_),
    .B(_05224_),
    .A_N(_05219_));
 sg13g2_nand2_1 _15567_ (.Y(_05226_),
    .A(_05219_),
    .B(_05223_));
 sg13g2_nor2_1 _15568_ (.A(_05219_),
    .B(_05223_),
    .Y(_05227_));
 sg13g2_nor2_2 _15569_ (.A(_05224_),
    .B(_05227_),
    .Y(_05228_));
 sg13g2_o21ai_1 _15570_ (.B1(_05225_),
    .Y(_05229_),
    .A1(_05224_),
    .A2(_05227_));
 sg13g2_a21oi_1 _15571_ (.A1(_04937_),
    .A2(_04940_),
    .Y(_05230_),
    .B1(_04944_));
 sg13g2_nor3_1 _15572_ (.A(_04899_),
    .B(_04941_),
    .C(_05230_),
    .Y(_05232_));
 sg13g2_o21ai_1 _15573_ (.B1(_04899_),
    .Y(_05233_),
    .A1(_04941_),
    .A2(_05230_));
 sg13g2_nor2b_1 _15574_ (.A(_05232_),
    .B_N(_05233_),
    .Y(_05234_));
 sg13g2_nand2_1 _15575_ (.Y(_05235_),
    .A(_04947_),
    .B(_04954_));
 sg13g2_o21ai_1 _15576_ (.B1(_05235_),
    .Y(_05236_),
    .A1(_04951_),
    .A2(_04953_));
 sg13g2_xnor2_1 _15577_ (.Y(_05237_),
    .A(_05234_),
    .B(_05236_));
 sg13g2_a21oi_1 _15578_ (.A1(_05226_),
    .A2(_05229_),
    .Y(_05238_),
    .B1(_05237_));
 sg13g2_and3_1 _15579_ (.X(_05239_),
    .A(_05226_),
    .B(_05229_),
    .C(_05237_));
 sg13g2_inv_1 _15580_ (.Y(_05240_),
    .A(_05239_));
 sg13g2_o21ai_1 _15581_ (.B1(_04988_),
    .Y(_05241_),
    .A1(_04989_),
    .A2(_04994_));
 sg13g2_o21ai_1 _15582_ (.B1(_04960_),
    .Y(_05243_),
    .A1(_04962_),
    .A2(_04963_));
 sg13g2_nand2_2 _15583_ (.Y(_05244_),
    .A(_04964_),
    .B(_05243_));
 sg13g2_nor2_1 _15584_ (.A(_05241_),
    .B(_05244_),
    .Y(_05245_));
 sg13g2_xnor2_1 _15585_ (.Y(_05246_),
    .A(_05241_),
    .B(_05244_));
 sg13g2_a21oi_2 _15586_ (.B1(_05006_),
    .Y(_05247_),
    .A2(_05005_),
    .A1(_04998_));
 sg13g2_xnor2_1 _15587_ (.Y(_05248_),
    .A(_05246_),
    .B(_05247_));
 sg13g2_o21ai_1 _15588_ (.B1(_05240_),
    .Y(_05249_),
    .A1(_05238_),
    .A2(_05248_));
 sg13g2_a21oi_1 _15589_ (.A1(_04718_),
    .A2(_04724_),
    .Y(_05250_),
    .B1(_04725_));
 sg13g2_nand2b_1 _15590_ (.Y(_05251_),
    .B(_04704_),
    .A_N(_05250_));
 sg13g2_nor2b_1 _15591_ (.A(_04704_),
    .B_N(_05250_),
    .Y(_05252_));
 sg13g2_xor2_1 _15592_ (.B(_05250_),
    .A(_04704_),
    .X(_05254_));
 sg13g2_o21ai_1 _15593_ (.B1(_04714_),
    .Y(_05255_),
    .A1(_04710_),
    .A2(_04713_));
 sg13g2_xnor2_1 _15594_ (.Y(_05256_),
    .A(_05254_),
    .B(_05255_));
 sg13g2_nand2_1 _15595_ (.Y(_05257_),
    .A(_04757_),
    .B(_04761_));
 sg13g2_or2_1 _15596_ (.X(_05258_),
    .B(_04738_),
    .A(_04731_));
 sg13g2_a22oi_1 _15597_ (.Y(_05259_),
    .B1(_05258_),
    .B2(_04737_),
    .A2(_05257_),
    .A1(_04760_));
 sg13g2_nand4_1 _15598_ (.B(_04760_),
    .C(_05257_),
    .A(_04737_),
    .Y(_05260_),
    .D(_05258_));
 sg13g2_nor2b_1 _15599_ (.A(_05259_),
    .B_N(_05260_),
    .Y(_05261_));
 sg13g2_a21oi_2 _15600_ (.B1(_04754_),
    .Y(_05262_),
    .A2(_04753_),
    .A1(_04747_));
 sg13g2_xnor2_1 _15601_ (.Y(_05263_),
    .A(_05261_),
    .B(_05262_));
 sg13g2_nor2b_1 _15602_ (.A(_05263_),
    .B_N(_05256_),
    .Y(_05265_));
 sg13g2_nand2b_1 _15603_ (.Y(_05266_),
    .B(_05263_),
    .A_N(_05256_));
 sg13g2_o21ai_1 _15604_ (.B1(_04909_),
    .Y(_05267_),
    .A1(_04679_),
    .A2(_04905_));
 sg13g2_a21oi_2 _15605_ (.B1(_04918_),
    .Y(_05268_),
    .A2(_04917_),
    .A1(_04912_));
 sg13g2_a21o_1 _15606_ (.A2(_04768_),
    .A1(_02704_),
    .B1(_04767_),
    .X(_05269_));
 sg13g2_o21ai_1 _15607_ (.B1(_05269_),
    .Y(_05270_),
    .A1(_02704_),
    .A2(_04768_));
 sg13g2_nand2_1 _15608_ (.Y(_05271_),
    .A(_05268_),
    .B(_05270_));
 sg13g2_nor2_1 _15609_ (.A(_05268_),
    .B(_05270_),
    .Y(_05272_));
 sg13g2_xor2_1 _15610_ (.B(_05270_),
    .A(_05268_),
    .X(_05273_));
 sg13g2_xnor2_1 _15611_ (.Y(_05274_),
    .A(_05267_),
    .B(_05273_));
 sg13g2_o21ai_1 _15612_ (.B1(_05266_),
    .Y(_05276_),
    .A1(_05265_),
    .A2(_05274_));
 sg13g2_or2_1 _15613_ (.X(_05277_),
    .B(_05276_),
    .A(_05249_));
 sg13g2_nand2_1 _15614_ (.Y(_05278_),
    .A(_05249_),
    .B(_05276_));
 sg13g2_nand2_1 _15615_ (.Y(_05279_),
    .A(_05277_),
    .B(_05278_));
 sg13g2_xor2_1 _15616_ (.B(_05279_),
    .A(_05218_),
    .X(_05280_));
 sg13g2_nand2_1 _15617_ (.Y(_05281_),
    .A(_04971_),
    .B(_04976_));
 sg13g2_a21oi_1 _15618_ (.A1(_04977_),
    .A2(_05281_),
    .Y(_05282_),
    .B1(_05029_));
 sg13g2_nand3_1 _15619_ (.B(_05029_),
    .C(_05281_),
    .A(_04977_),
    .Y(_05283_));
 sg13g2_nor2_1 _15620_ (.A(_05054_),
    .B(_05073_),
    .Y(_05284_));
 sg13g2_o21ai_1 _15621_ (.B1(_05283_),
    .Y(_05285_),
    .A1(_05282_),
    .A2(_05284_));
 sg13g2_nand2_1 _15622_ (.Y(_05287_),
    .A(_05192_),
    .B(_05195_));
 sg13g2_nand2_1 _15623_ (.Y(_05288_),
    .A(_05191_),
    .B(_05287_));
 sg13g2_nand2_1 _15624_ (.Y(_05289_),
    .A(_05109_),
    .B(_05150_));
 sg13g2_and3_1 _15625_ (.X(_05290_),
    .A(_05108_),
    .B(_05288_),
    .C(_05289_));
 sg13g2_a21oi_1 _15626_ (.A1(_05108_),
    .A2(_05289_),
    .Y(_05291_),
    .B1(_05288_));
 sg13g2_o21ai_1 _15627_ (.B1(_05205_),
    .Y(_05292_),
    .A1(_05204_),
    .A2(_05208_));
 sg13g2_nor2_1 _15628_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sg13g2_nor2_1 _15629_ (.A(_05290_),
    .B(_05293_),
    .Y(_05294_));
 sg13g2_nor2_1 _15630_ (.A(_05285_),
    .B(_05294_),
    .Y(_05295_));
 sg13g2_and2_1 _15631_ (.A(_05285_),
    .B(_05294_),
    .X(_05296_));
 sg13g2_nor2_1 _15632_ (.A(_05295_),
    .B(_05296_),
    .Y(_05298_));
 sg13g2_nor2_2 _15633_ (.A(_05100_),
    .B(_05105_),
    .Y(_05299_));
 sg13g2_a21oi_2 _15634_ (.B1(_05135_),
    .Y(_05300_),
    .A2(_05149_),
    .A1(_05136_));
 sg13g2_nand2_1 _15635_ (.Y(_05301_),
    .A(_05299_),
    .B(_05300_));
 sg13g2_nor2_1 _15636_ (.A(_05299_),
    .B(_05300_),
    .Y(_05302_));
 sg13g2_nand2_2 _15637_ (.Y(_05303_),
    .A(_05173_),
    .B(_05186_));
 sg13g2_a21oi_2 _15638_ (.B1(_05302_),
    .Y(_05304_),
    .A2(_05303_),
    .A1(_05301_));
 sg13g2_xnor2_1 _15639_ (.Y(_05305_),
    .A(_05298_),
    .B(_05304_));
 sg13g2_nand2_1 _15640_ (.Y(_05306_),
    .A(_05280_),
    .B(_05305_));
 sg13g2_xor2_1 _15641_ (.B(_05305_),
    .A(_05280_),
    .X(_05307_));
 sg13g2_o21ai_1 _15642_ (.B1(_04969_),
    .Y(_05309_),
    .A1(_05280_),
    .A2(_05305_));
 sg13g2_nand2_1 _15643_ (.Y(_05310_),
    .A(_05306_),
    .B(_05309_));
 sg13g2_xnor2_1 _15644_ (.Y(_05311_),
    .A(_04969_),
    .B(_05307_));
 sg13g2_a22oi_1 _15645_ (.Y(_05312_),
    .B1(_05216_),
    .B2(_05217_),
    .A2(_05211_),
    .A1(_05031_));
 sg13g2_nor2_1 _15646_ (.A(_05290_),
    .B(_05291_),
    .Y(_05313_));
 sg13g2_xnor2_1 _15647_ (.Y(_05314_),
    .A(_05292_),
    .B(_05313_));
 sg13g2_nor2_1 _15648_ (.A(_05312_),
    .B(_05314_),
    .Y(_05315_));
 sg13g2_xnor2_1 _15649_ (.Y(_05316_),
    .A(_05312_),
    .B(_05314_));
 sg13g2_nand2b_1 _15650_ (.Y(_05317_),
    .B(_05283_),
    .A_N(_05282_));
 sg13g2_xnor2_1 _15651_ (.Y(_05318_),
    .A(_05284_),
    .B(_05317_));
 sg13g2_xnor2_1 _15652_ (.Y(_05320_),
    .A(_05316_),
    .B(_05318_));
 sg13g2_xor2_1 _15653_ (.B(_05300_),
    .A(_05299_),
    .X(_05321_));
 sg13g2_xnor2_1 _15654_ (.Y(_05322_),
    .A(_05303_),
    .B(_05321_));
 sg13g2_xor2_1 _15655_ (.B(_04836_),
    .A(_04798_),
    .X(_05323_));
 sg13g2_xnor2_1 _15656_ (.Y(_05324_),
    .A(_04864_),
    .B(_05323_));
 sg13g2_and2_1 _15657_ (.A(_05322_),
    .B(_05324_),
    .X(_05325_));
 sg13g2_or2_1 _15658_ (.X(_05326_),
    .B(_05324_),
    .A(_05322_));
 sg13g2_nor2b_1 _15659_ (.A(_05325_),
    .B_N(_05326_),
    .Y(_05327_));
 sg13g2_nor2_1 _15660_ (.A(_04744_),
    .B(_04745_),
    .Y(_05328_));
 sg13g2_xnor2_1 _15661_ (.Y(_05329_),
    .A(_04771_),
    .B(_05328_));
 sg13g2_xnor2_1 _15662_ (.Y(_05331_),
    .A(_05327_),
    .B(_05329_));
 sg13g2_inv_1 _15663_ (.Y(_05332_),
    .A(_05331_));
 sg13g2_nand2_1 _15664_ (.Y(_05333_),
    .A(_05320_),
    .B(_05332_));
 sg13g2_or2_1 _15665_ (.X(_05334_),
    .B(_05084_),
    .A(_05071_));
 sg13g2_and2_1 _15666_ (.A(_05071_),
    .B(_05084_),
    .X(_05335_));
 sg13g2_inv_1 _15667_ (.Y(_05336_),
    .A(_05335_));
 sg13g2_nand2_1 _15668_ (.Y(_05337_),
    .A(_05334_),
    .B(_05336_));
 sg13g2_xnor2_1 _15669_ (.Y(_05338_),
    .A(_05096_),
    .B(_05337_));
 sg13g2_nand2b_1 _15670_ (.Y(_05339_),
    .B(_04935_),
    .A_N(_04934_));
 sg13g2_xnor2_1 _15671_ (.Y(_05340_),
    .A(_04967_),
    .B(_05339_));
 sg13g2_a21o_1 _15672_ (.A2(_05037_),
    .A1(_05035_),
    .B1(_05034_),
    .X(_05342_));
 sg13g2_a21o_1 _15673_ (.A2(_05009_),
    .A1(_04995_),
    .B1(_05024_),
    .X(_05343_));
 sg13g2_a22oi_1 _15674_ (.Y(_05344_),
    .B1(_05343_),
    .B2(_05010_),
    .A2(_05342_),
    .A1(_05038_));
 sg13g2_nand4_1 _15675_ (.B(_05038_),
    .C(_05342_),
    .A(_05010_),
    .Y(_05345_),
    .D(_05343_));
 sg13g2_nor2b_1 _15676_ (.A(_05344_),
    .B_N(_05345_),
    .Y(_05346_));
 sg13g2_xnor2_1 _15677_ (.Y(_05347_),
    .A(_05053_),
    .B(_05346_));
 sg13g2_nor2_1 _15678_ (.A(_05340_),
    .B(_05347_),
    .Y(_05348_));
 sg13g2_nand2_1 _15679_ (.Y(_05349_),
    .A(_05340_),
    .B(_05347_));
 sg13g2_nor2b_1 _15680_ (.A(_05348_),
    .B_N(_05349_),
    .Y(_05350_));
 sg13g2_xnor2_1 _15681_ (.Y(_05351_),
    .A(_05338_),
    .B(_05350_));
 sg13g2_o21ai_1 _15682_ (.B1(_05351_),
    .Y(_05353_),
    .A1(_05320_),
    .A2(_05332_));
 sg13g2_nand2_1 _15683_ (.Y(_05354_),
    .A(_05333_),
    .B(_05353_));
 sg13g2_nor2b_1 _15684_ (.A(_05265_),
    .B_N(_05266_),
    .Y(_05355_));
 sg13g2_xnor2_1 _15685_ (.Y(_05356_),
    .A(_05274_),
    .B(_05355_));
 sg13g2_nand2b_1 _15686_ (.Y(_05357_),
    .B(_04783_),
    .A_N(_04780_));
 sg13g2_a21oi_1 _15687_ (.A1(_04784_),
    .A2(_05357_),
    .Y(_05358_),
    .B1(_04833_));
 sg13g2_inv_1 _15688_ (.Y(_05359_),
    .A(_05358_));
 sg13g2_and3_1 _15689_ (.X(_05360_),
    .A(_04784_),
    .B(_04833_),
    .C(_05357_));
 sg13g2_nor2_1 _15690_ (.A(_05358_),
    .B(_05360_),
    .Y(_05361_));
 sg13g2_o21ai_1 _15691_ (.B1(_04773_),
    .Y(_05362_),
    .A1(_04775_),
    .A2(_04776_));
 sg13g2_nand2_1 _15692_ (.Y(_05364_),
    .A(_04777_),
    .B(_05362_));
 sg13g2_xnor2_1 _15693_ (.Y(_05365_),
    .A(_05361_),
    .B(_05364_));
 sg13g2_nor2_1 _15694_ (.A(_04792_),
    .B(_04795_),
    .Y(_05366_));
 sg13g2_a21o_1 _15695_ (.A2(_04852_),
    .A1(_02504_),
    .B1(_04850_),
    .X(_05367_));
 sg13g2_o21ai_1 _15696_ (.B1(_05367_),
    .Y(_05368_),
    .A1(_02504_),
    .A2(_04852_));
 sg13g2_nor2b_1 _15697_ (.A(_05366_),
    .B_N(_05368_),
    .Y(_05369_));
 sg13g2_nor2b_1 _15698_ (.A(_05368_),
    .B_N(_05366_),
    .Y(_05370_));
 sg13g2_nor2_1 _15699_ (.A(_05369_),
    .B(_05370_),
    .Y(_05371_));
 sg13g2_xnor2_1 _15700_ (.Y(_05372_),
    .A(_04846_),
    .B(_05371_));
 sg13g2_nand2_1 _15701_ (.Y(_05373_),
    .A(_05365_),
    .B(_05372_));
 sg13g2_xnor2_1 _15702_ (.Y(_05375_),
    .A(_05365_),
    .B(_05372_));
 sg13g2_o21ai_1 _15703_ (.B1(_04860_),
    .Y(_05376_),
    .A1(_04855_),
    .A2(_04859_));
 sg13g2_inv_1 _15704_ (.Y(_05377_),
    .A(_05376_));
 sg13g2_nand2_1 _15705_ (.Y(_05378_),
    .A(_04678_),
    .B(_04683_));
 sg13g2_nand2_2 _15706_ (.Y(_05379_),
    .A(_04682_),
    .B(_05378_));
 sg13g2_nor2_1 _15707_ (.A(_05377_),
    .B(_05379_),
    .Y(_05380_));
 sg13g2_nand2_1 _15708_ (.Y(_05381_),
    .A(_05377_),
    .B(_05379_));
 sg13g2_nor2b_1 _15709_ (.A(_05380_),
    .B_N(_05381_),
    .Y(_05382_));
 sg13g2_a21oi_1 _15710_ (.A1(_02703_),
    .A2(_04690_),
    .Y(_05383_),
    .B1(_04691_));
 sg13g2_inv_1 _15711_ (.Y(_05384_),
    .A(_05383_));
 sg13g2_xnor2_1 _15712_ (.Y(_05386_),
    .A(_05382_),
    .B(_05384_));
 sg13g2_xnor2_1 _15713_ (.Y(_05387_),
    .A(_05375_),
    .B(_05386_));
 sg13g2_nand2b_1 _15714_ (.Y(_05388_),
    .B(net2469),
    .A_N(_05102_));
 sg13g2_a22oi_1 _15715_ (.Y(_05389_),
    .B1(_05388_),
    .B2(_05101_),
    .A2(_05102_),
    .A1(_00018_));
 sg13g2_nand2_1 _15716_ (.Y(_05390_),
    .A(_05133_),
    .B(_05389_));
 sg13g2_nor2_1 _15717_ (.A(_05133_),
    .B(_05389_),
    .Y(_05391_));
 sg13g2_xor2_1 _15718_ (.B(_05389_),
    .A(_05133_),
    .X(_05392_));
 sg13g2_o21ai_1 _15719_ (.B1(_05118_),
    .Y(_05393_),
    .A1(_05112_),
    .A2(_05117_));
 sg13g2_xnor2_1 _15720_ (.Y(_05394_),
    .A(_05392_),
    .B(_05393_));
 sg13g2_a21oi_2 _15721_ (.B1(_05158_),
    .Y(_05395_),
    .A2(_05159_),
    .A1(_05155_));
 sg13g2_nor2_1 _15722_ (.A(_05163_),
    .B(_05169_),
    .Y(_05397_));
 sg13g2_nor3_1 _15723_ (.A(_05147_),
    .B(_05170_),
    .C(_05397_),
    .Y(_05398_));
 sg13g2_o21ai_1 _15724_ (.B1(_05147_),
    .Y(_05399_),
    .A1(_05170_),
    .A2(_05397_));
 sg13g2_nor2b_1 _15725_ (.A(_05398_),
    .B_N(_05399_),
    .Y(_05400_));
 sg13g2_xnor2_1 _15726_ (.Y(_05401_),
    .A(_05395_),
    .B(_05400_));
 sg13g2_nand2b_2 _15727_ (.Y(_05402_),
    .B(_05401_),
    .A_N(_05394_));
 sg13g2_nand2b_1 _15728_ (.Y(_05403_),
    .B(_05394_),
    .A_N(_05401_));
 sg13g2_nand2_1 _15729_ (.Y(_05404_),
    .A(_05402_),
    .B(_05403_));
 sg13g2_a21o_1 _15730_ (.A2(_04808_),
    .A1(_04805_),
    .B1(_04801_),
    .X(_05405_));
 sg13g2_o21ai_1 _15731_ (.B1(_05405_),
    .Y(_05406_),
    .A1(_04805_),
    .A2(_04808_));
 sg13g2_o21ai_1 _15732_ (.B1(_05178_),
    .Y(_05408_),
    .A1(_05180_),
    .A2(_05182_));
 sg13g2_nand2b_1 _15733_ (.Y(_05409_),
    .B(_04812_),
    .A_N(_04819_));
 sg13g2_a22oi_1 _15734_ (.Y(_05410_),
    .B1(_05409_),
    .B2(_04818_),
    .A2(_05408_),
    .A1(_05183_));
 sg13g2_nand4_1 _15735_ (.B(_05183_),
    .C(_05408_),
    .A(_04818_),
    .Y(_05411_),
    .D(_05409_));
 sg13g2_nand2b_1 _15736_ (.Y(_05412_),
    .B(_05411_),
    .A_N(_05410_));
 sg13g2_o21ai_1 _15737_ (.B1(_05411_),
    .Y(_05413_),
    .A1(_05406_),
    .A2(_05410_));
 sg13g2_xnor2_1 _15738_ (.Y(_05414_),
    .A(_05406_),
    .B(_05412_));
 sg13g2_xor2_1 _15739_ (.B(_05414_),
    .A(_05404_),
    .X(_05415_));
 sg13g2_nand2_1 _15740_ (.Y(_05416_),
    .A(_05387_),
    .B(_05415_));
 sg13g2_xor2_1 _15741_ (.B(_05415_),
    .A(_05387_),
    .X(_05417_));
 sg13g2_xnor2_1 _15742_ (.Y(_05419_),
    .A(_05356_),
    .B(_05417_));
 sg13g2_xnor2_1 _15743_ (.Y(_05420_),
    .A(_05320_),
    .B(_05331_));
 sg13g2_xnor2_1 _15744_ (.Y(_05421_),
    .A(_05351_),
    .B(_05420_));
 sg13g2_nand2b_1 _15745_ (.Y(_05422_),
    .B(_05419_),
    .A_N(_05421_));
 sg13g2_nor2b_1 _15746_ (.A(_05419_),
    .B_N(_05421_),
    .Y(_05423_));
 sg13g2_xnor2_1 _15747_ (.Y(_05424_),
    .A(_05419_),
    .B(_05421_));
 sg13g2_nor2_1 _15748_ (.A(_05238_),
    .B(_05239_),
    .Y(_05425_));
 sg13g2_xnor2_1 _15749_ (.Y(_05426_),
    .A(_05248_),
    .B(_05425_));
 sg13g2_xnor2_1 _15750_ (.Y(_05427_),
    .A(_05424_),
    .B(_05426_));
 sg13g2_a21o_2 _15751_ (.A2(_05023_),
    .A1(_05018_),
    .B1(_05019_),
    .X(_05428_));
 sg13g2_a21oi_1 _15752_ (.A1(_05422_),
    .A2(_05426_),
    .Y(_05430_),
    .B1(_05423_));
 sg13g2_o21ai_1 _15753_ (.B1(_05430_),
    .Y(_05431_),
    .A1(_05427_),
    .A2(_05428_));
 sg13g2_inv_1 _15754_ (.Y(_05432_),
    .A(_05431_));
 sg13g2_nand3b_1 _15755_ (.B(_05423_),
    .C(_05426_),
    .Y(_05433_),
    .A_N(_05428_));
 sg13g2_a21o_1 _15756_ (.A2(_05433_),
    .A1(_05431_),
    .B1(_05354_),
    .X(_05434_));
 sg13g2_nand3_1 _15757_ (.B(_05431_),
    .C(_05433_),
    .A(_05354_),
    .Y(_05435_));
 sg13g2_o21ai_1 _15758_ (.B1(_05326_),
    .Y(_05436_),
    .A1(_05325_),
    .A2(_05329_));
 sg13g2_o21ai_1 _15759_ (.B1(_05356_),
    .Y(_05437_),
    .A1(_05387_),
    .A2(_05415_));
 sg13g2_nand2_1 _15760_ (.Y(_05438_),
    .A(_05416_),
    .B(_05437_));
 sg13g2_inv_1 _15761_ (.Y(_05439_),
    .A(_05438_));
 sg13g2_a21oi_1 _15762_ (.A1(_05312_),
    .A2(_05314_),
    .Y(_05441_),
    .B1(_05318_));
 sg13g2_nor2_2 _15763_ (.A(_05315_),
    .B(_05441_),
    .Y(_05442_));
 sg13g2_nor2_1 _15764_ (.A(_05439_),
    .B(_05442_),
    .Y(_05443_));
 sg13g2_xnor2_1 _15765_ (.Y(_05444_),
    .A(_05438_),
    .B(_05442_));
 sg13g2_xnor2_1 _15766_ (.Y(_05445_),
    .A(_05436_),
    .B(_05444_));
 sg13g2_a21o_1 _15767_ (.A2(_05435_),
    .A1(_05434_),
    .B1(_05445_),
    .X(_05446_));
 sg13g2_nand3_1 _15768_ (.B(_05435_),
    .C(_05445_),
    .A(_05434_),
    .Y(_05447_));
 sg13g2_o21ai_1 _15769_ (.B1(_05386_),
    .Y(_05448_),
    .A1(_05365_),
    .A2(_05372_));
 sg13g2_nand2_2 _15770_ (.Y(_05449_),
    .A(_05373_),
    .B(_05448_));
 sg13g2_nand2b_2 _15771_ (.Y(_05450_),
    .B(_05403_),
    .A_N(_05414_));
 sg13g2_a21oi_1 _15772_ (.A1(_05338_),
    .A2(_05349_),
    .Y(_05452_),
    .B1(_05348_));
 sg13g2_nand3_1 _15773_ (.B(_05450_),
    .C(_05452_),
    .A(_05402_),
    .Y(_05453_));
 sg13g2_a21o_1 _15774_ (.A2(_05450_),
    .A1(_05402_),
    .B1(_05452_),
    .X(_05454_));
 sg13g2_nand2_1 _15775_ (.Y(_05455_),
    .A(_05453_),
    .B(_05454_));
 sg13g2_nand2_1 _15776_ (.Y(_05456_),
    .A(_05449_),
    .B(_05453_));
 sg13g2_nand2_2 _15777_ (.Y(_05457_),
    .A(_05454_),
    .B(_05456_));
 sg13g2_inv_1 _15778_ (.Y(_05458_),
    .A(_05457_));
 sg13g2_xor2_1 _15779_ (.B(_05455_),
    .A(_05449_),
    .X(_05459_));
 sg13g2_nand3_1 _15780_ (.B(_05447_),
    .C(_05459_),
    .A(_05446_),
    .Y(_05460_));
 sg13g2_a21o_1 _15781_ (.A2(_05447_),
    .A1(_05446_),
    .B1(_05459_),
    .X(_05461_));
 sg13g2_nand3_1 _15782_ (.B(_05460_),
    .C(_05461_),
    .A(_05311_),
    .Y(_05463_));
 sg13g2_a21oi_1 _15783_ (.A1(_05460_),
    .A2(_05461_),
    .Y(_05464_),
    .B1(_05311_));
 sg13g2_a21o_1 _15784_ (.A2(_05461_),
    .A1(_05460_),
    .B1(_05311_),
    .X(_05465_));
 sg13g2_a21oi_2 _15785_ (.B1(_05398_),
    .Y(_05466_),
    .A2(_05399_),
    .A1(_05395_));
 sg13g2_nand2_1 _15786_ (.Y(_05467_),
    .A(_05413_),
    .B(_05466_));
 sg13g2_xor2_1 _15787_ (.B(_05466_),
    .A(_05413_),
    .X(_05468_));
 sg13g2_o21ai_1 _15788_ (.B1(_05359_),
    .Y(_05469_),
    .A1(_05360_),
    .A2(_05364_));
 sg13g2_xnor2_1 _15789_ (.Y(_05470_),
    .A(_05468_),
    .B(_05469_));
 sg13g2_o21ai_1 _15790_ (.B1(_05334_),
    .Y(_05471_),
    .A1(_05096_),
    .A2(_05335_));
 sg13g2_a21oi_1 _15791_ (.A1(_05053_),
    .A2(_05345_),
    .Y(_05472_),
    .B1(_05344_));
 sg13g2_nor2_1 _15792_ (.A(_05471_),
    .B(_05472_),
    .Y(_05474_));
 sg13g2_and2_1 _15793_ (.A(_05471_),
    .B(_05472_),
    .X(_05475_));
 sg13g2_nor2_1 _15794_ (.A(_05474_),
    .B(_05475_),
    .Y(_05476_));
 sg13g2_a21oi_2 _15795_ (.B1(_05391_),
    .Y(_05477_),
    .A2(_05393_),
    .A1(_05390_));
 sg13g2_xor2_1 _15796_ (.B(_05477_),
    .A(_05476_),
    .X(_05478_));
 sg13g2_nand2_1 _15797_ (.Y(_05479_),
    .A(_05470_),
    .B(_05478_));
 sg13g2_nor2_1 _15798_ (.A(_05470_),
    .B(_05478_),
    .Y(_05480_));
 sg13g2_inv_1 _15799_ (.Y(_05481_),
    .A(_05480_));
 sg13g2_nand2_1 _15800_ (.Y(_05482_),
    .A(_05479_),
    .B(_05481_));
 sg13g2_nor2_1 _15801_ (.A(_04846_),
    .B(_05370_),
    .Y(_05483_));
 sg13g2_o21ai_1 _15802_ (.B1(_05381_),
    .Y(_05485_),
    .A1(_05380_),
    .A2(_05384_));
 sg13g2_o21ai_1 _15803_ (.B1(_05485_),
    .Y(_05486_),
    .A1(_05369_),
    .A2(_05483_));
 sg13g2_or3_1 _15804_ (.A(_05369_),
    .B(_05483_),
    .C(_05485_),
    .X(_05487_));
 sg13g2_nand2_1 _15805_ (.Y(_05488_),
    .A(_05486_),
    .B(_05487_));
 sg13g2_o21ai_1 _15806_ (.B1(_05251_),
    .Y(_05489_),
    .A1(_05252_),
    .A2(_05255_));
 sg13g2_xnor2_1 _15807_ (.Y(_05490_),
    .A(_05488_),
    .B(_05489_));
 sg13g2_xor2_1 _15808_ (.B(_05490_),
    .A(_05482_),
    .X(_05491_));
 sg13g2_inv_1 _15809_ (.Y(_05492_),
    .A(_05491_));
 sg13g2_and3_1 _15810_ (.X(_05493_),
    .A(_05463_),
    .B(_05465_),
    .C(_05492_));
 sg13g2_a21oi_1 _15811_ (.A1(_05463_),
    .A2(_05465_),
    .Y(_05494_),
    .B1(_05492_));
 sg13g2_nor2_1 _15812_ (.A(_05493_),
    .B(_05494_),
    .Y(_05496_));
 sg13g2_o21ai_1 _15813_ (.B1(_05233_),
    .Y(_05497_),
    .A1(_05232_),
    .A2(_05236_));
 sg13g2_a21oi_2 _15814_ (.B1(_05259_),
    .Y(_05498_),
    .A2(_05262_),
    .A1(_05260_));
 sg13g2_a21oi_2 _15815_ (.B1(_05272_),
    .Y(_05499_),
    .A2(_05271_),
    .A1(_05267_));
 sg13g2_nand2b_1 _15816_ (.Y(_05500_),
    .B(_05499_),
    .A_N(_05498_));
 sg13g2_inv_1 _15817_ (.Y(_05501_),
    .A(_05500_));
 sg13g2_nand2b_1 _15818_ (.Y(_05502_),
    .B(_05498_),
    .A_N(_05499_));
 sg13g2_and2_1 _15819_ (.A(_05500_),
    .B(_05502_),
    .X(_05503_));
 sg13g2_xnor2_1 _15820_ (.Y(_05504_),
    .A(_05228_),
    .B(_05503_));
 sg13g2_nor2_1 _15821_ (.A(_05497_),
    .B(_05504_),
    .Y(_05505_));
 sg13g2_nand2_1 _15822_ (.Y(_05507_),
    .A(_05497_),
    .B(_05504_));
 sg13g2_nand2b_1 _15823_ (.Y(_05508_),
    .B(_05507_),
    .A_N(_05505_));
 sg13g2_a21oi_1 _15824_ (.A1(_05241_),
    .A2(_05244_),
    .Y(_05509_),
    .B1(_05247_));
 sg13g2_nor2_1 _15825_ (.A(_05245_),
    .B(_05509_),
    .Y(_05510_));
 sg13g2_xnor2_1 _15826_ (.Y(_05511_),
    .A(_05508_),
    .B(_05510_));
 sg13g2_nor3_1 _15827_ (.A(_05493_),
    .B(_05494_),
    .C(_05511_),
    .Y(_05512_));
 sg13g2_a21oi_1 _15828_ (.A1(_05463_),
    .A2(_05492_),
    .Y(_05513_),
    .B1(_05464_));
 sg13g2_nor2b_1 _15829_ (.A(_05512_),
    .B_N(_05513_),
    .Y(_05514_));
 sg13g2_nor3_1 _15830_ (.A(_05465_),
    .B(_05491_),
    .C(_05511_),
    .Y(_05515_));
 sg13g2_nand2_1 _15831_ (.Y(_05516_),
    .A(_05446_),
    .B(_05459_));
 sg13g2_and2_1 _15832_ (.A(_05447_),
    .B(_05516_),
    .X(_05518_));
 sg13g2_nor2_1 _15833_ (.A(_05515_),
    .B(_05518_),
    .Y(_05519_));
 sg13g2_a21o_1 _15834_ (.A2(_05490_),
    .A1(_05479_),
    .B1(_05480_),
    .X(_05520_));
 sg13g2_or2_1 _15835_ (.X(_05521_),
    .B(_05520_),
    .A(_05310_));
 sg13g2_and2_1 _15836_ (.A(_05310_),
    .B(_05520_),
    .X(_05522_));
 sg13g2_o21ai_1 _15837_ (.B1(_05507_),
    .Y(_05523_),
    .A1(_05505_),
    .A2(_05510_));
 sg13g2_a21oi_2 _15838_ (.B1(_05522_),
    .Y(_05524_),
    .A2(_05523_),
    .A1(_05521_));
 sg13g2_o21ai_1 _15839_ (.B1(_05524_),
    .Y(_05525_),
    .A1(_05514_),
    .A2(_05519_));
 sg13g2_or3_1 _15840_ (.A(_05514_),
    .B(_05519_),
    .C(_05524_),
    .X(_05526_));
 sg13g2_o21ai_1 _15841_ (.B1(_05433_),
    .Y(_05527_),
    .A1(_05354_),
    .A2(_05432_));
 sg13g2_nor2_1 _15842_ (.A(_05436_),
    .B(_05443_),
    .Y(_05529_));
 sg13g2_a21oi_2 _15843_ (.B1(_05529_),
    .Y(_05530_),
    .A2(_05442_),
    .A1(_05439_));
 sg13g2_nor2_1 _15844_ (.A(_05527_),
    .B(_05530_),
    .Y(_05531_));
 sg13g2_nand2_1 _15845_ (.Y(_05532_),
    .A(_05527_),
    .B(_05530_));
 sg13g2_o21ai_1 _15846_ (.B1(_05532_),
    .Y(_05533_),
    .A1(_05458_),
    .A2(_05531_));
 sg13g2_nand2_1 _15847_ (.Y(_05534_),
    .A(_05525_),
    .B(_05533_));
 sg13g2_nand2_2 _15848_ (.Y(_05535_),
    .A(_05526_),
    .B(_05534_));
 sg13g2_nand2_1 _15849_ (.Y(_05536_),
    .A(_05525_),
    .B(_05526_));
 sg13g2_xor2_1 _15850_ (.B(_05536_),
    .A(_05533_),
    .X(_05537_));
 sg13g2_xor2_1 _15851_ (.B(_05513_),
    .A(_05512_),
    .X(_05538_));
 sg13g2_xor2_1 _15852_ (.B(_05538_),
    .A(_05518_),
    .X(_05540_));
 sg13g2_or2_1 _15853_ (.X(_05541_),
    .B(_05523_),
    .A(_05521_));
 sg13g2_a22oi_1 _15854_ (.Y(_05542_),
    .B1(_05524_),
    .B2(_05541_),
    .A2(_05523_),
    .A1(_05522_));
 sg13g2_nor2b_1 _15855_ (.A(_05531_),
    .B_N(_05532_),
    .Y(_05543_));
 sg13g2_xnor2_1 _15856_ (.Y(_05544_),
    .A(_05457_),
    .B(_05543_));
 sg13g2_a21o_1 _15857_ (.A2(_05542_),
    .A1(_05540_),
    .B1(_05544_),
    .X(_05545_));
 sg13g2_o21ai_1 _15858_ (.B1(_05545_),
    .Y(_05546_),
    .A1(_05540_),
    .A2(_05542_));
 sg13g2_xor2_1 _15859_ (.B(_05542_),
    .A(_05540_),
    .X(_05547_));
 sg13g2_xnor2_1 _15860_ (.Y(_05548_),
    .A(_05544_),
    .B(_05547_));
 sg13g2_o21ai_1 _15861_ (.B1(_05469_),
    .Y(_05549_),
    .A1(_05413_),
    .A2(_05466_));
 sg13g2_nand2_1 _15862_ (.Y(_05551_),
    .A(_05467_),
    .B(_05549_));
 sg13g2_nor2_1 _15863_ (.A(_05475_),
    .B(_05477_),
    .Y(_05552_));
 sg13g2_nor3_1 _15864_ (.A(_05474_),
    .B(_05551_),
    .C(_05552_),
    .Y(_05553_));
 sg13g2_o21ai_1 _15865_ (.B1(_05551_),
    .Y(_05554_),
    .A1(_05474_),
    .A2(_05552_));
 sg13g2_nor2b_1 _15866_ (.A(_05553_),
    .B_N(_05554_),
    .Y(_05555_));
 sg13g2_nand2_1 _15867_ (.Y(_05556_),
    .A(_05487_),
    .B(_05489_));
 sg13g2_nand2_2 _15868_ (.Y(_05557_),
    .A(_05486_),
    .B(_05556_));
 sg13g2_inv_1 _15869_ (.Y(_05558_),
    .A(_05557_));
 sg13g2_xnor2_1 _15870_ (.Y(_05559_),
    .A(_05555_),
    .B(_05557_));
 sg13g2_nor2_1 _15871_ (.A(_05295_),
    .B(_05304_),
    .Y(_05560_));
 sg13g2_nor2_1 _15872_ (.A(_05296_),
    .B(_05560_),
    .Y(_05562_));
 sg13g2_nand2b_1 _15873_ (.Y(_05563_),
    .B(_05277_),
    .A_N(_05218_));
 sg13g2_a21oi_1 _15874_ (.A1(_05278_),
    .A2(_05563_),
    .Y(_05564_),
    .B1(_05562_));
 sg13g2_nand3_1 _15875_ (.B(_05562_),
    .C(_05563_),
    .A(_05278_),
    .Y(_05565_));
 sg13g2_nor2b_1 _15876_ (.A(_05564_),
    .B_N(_05565_),
    .Y(_05566_));
 sg13g2_nand2_1 _15877_ (.Y(_05567_),
    .A(_04867_),
    .B(_04968_));
 sg13g2_nand2_1 _15878_ (.Y(_05568_),
    .A(_04868_),
    .B(_05567_));
 sg13g2_xnor2_1 _15879_ (.Y(_05569_),
    .A(_05566_),
    .B(_05568_));
 sg13g2_nor2_1 _15880_ (.A(_05559_),
    .B(_05569_),
    .Y(_05570_));
 sg13g2_nand2_1 _15881_ (.Y(_05571_),
    .A(_05559_),
    .B(_05569_));
 sg13g2_nor2b_1 _15882_ (.A(_05570_),
    .B_N(_05571_),
    .Y(_05573_));
 sg13g2_o21ai_1 _15883_ (.B1(_05502_),
    .Y(_05574_),
    .A1(_05228_),
    .A2(_05501_));
 sg13g2_xnor2_1 _15884_ (.Y(_05575_),
    .A(_05573_),
    .B(_05574_));
 sg13g2_inv_1 _15885_ (.Y(_05576_),
    .A(_05575_));
 sg13g2_a21o_1 _15886_ (.A2(_05576_),
    .A1(_05548_),
    .B1(_05546_),
    .X(_05577_));
 sg13g2_nand3_1 _15887_ (.B(_05548_),
    .C(_05576_),
    .A(_05546_),
    .Y(_05578_));
 sg13g2_o21ai_1 _15888_ (.B1(_05571_),
    .Y(_05579_),
    .A1(_05570_),
    .A2(_05574_));
 sg13g2_nand3_1 _15889_ (.B(_05578_),
    .C(_05579_),
    .A(_05577_),
    .Y(_05580_));
 sg13g2_a21o_1 _15890_ (.A2(_05578_),
    .A1(_05577_),
    .B1(_05579_),
    .X(_05581_));
 sg13g2_and3_1 _15891_ (.X(_05582_),
    .A(_05537_),
    .B(_05580_),
    .C(_05581_));
 sg13g2_nand3_1 _15892_ (.B(_05580_),
    .C(_05581_),
    .A(_05537_),
    .Y(_05584_));
 sg13g2_a21oi_2 _15893_ (.B1(_05537_),
    .Y(_05585_),
    .A2(_05581_),
    .A1(_05580_));
 sg13g2_a21oi_2 _15894_ (.B1(_05564_),
    .Y(_05586_),
    .A2(_05568_),
    .A1(_05565_));
 sg13g2_inv_1 _15895_ (.Y(_05587_),
    .A(_05586_));
 sg13g2_nor3_1 _15896_ (.A(_05582_),
    .B(_05585_),
    .C(_05586_),
    .Y(_05588_));
 sg13g2_o21ai_1 _15897_ (.B1(_05586_),
    .Y(_05589_),
    .A1(_05582_),
    .A2(_05585_));
 sg13g2_nor2b_1 _15898_ (.A(_05588_),
    .B_N(_05589_),
    .Y(_05590_));
 sg13g2_o21ai_1 _15899_ (.B1(_05554_),
    .Y(_05591_),
    .A1(_05553_),
    .A2(_05558_));
 sg13g2_nand3b_1 _15900_ (.B(_05589_),
    .C(_05591_),
    .Y(_05592_),
    .A_N(_05588_));
 sg13g2_o21ai_1 _15901_ (.B1(_05584_),
    .Y(_05593_),
    .A1(_05585_),
    .A2(_05587_));
 sg13g2_nand4_1 _15902_ (.B(_05585_),
    .C(_05587_),
    .A(_05584_),
    .Y(_05595_),
    .D(_05591_));
 sg13g2_xnor2_1 _15903_ (.Y(_05596_),
    .A(_05592_),
    .B(_05593_));
 sg13g2_nand2_1 _15904_ (.Y(_05597_),
    .A(_05578_),
    .B(_05579_));
 sg13g2_and2_1 _15905_ (.A(_05577_),
    .B(_05597_),
    .X(_05598_));
 sg13g2_inv_1 _15906_ (.Y(_05599_),
    .A(_05598_));
 sg13g2_xnor2_1 _15907_ (.Y(_05600_),
    .A(_05596_),
    .B(_05599_));
 sg13g2_xnor2_1 _15908_ (.Y(_05601_),
    .A(_05596_),
    .B(_05598_));
 sg13g2_and2_1 _15909_ (.A(_05595_),
    .B(_05599_),
    .X(_05602_));
 sg13g2_a21oi_2 _15910_ (.B1(_05602_),
    .Y(_05603_),
    .A2(_05593_),
    .A1(_05592_));
 sg13g2_a21oi_2 _15911_ (.B1(_05603_),
    .Y(_05604_),
    .A2(_05601_),
    .A1(_05535_));
 sg13g2_a21o_2 _15912_ (.A2(_05601_),
    .A1(_05535_),
    .B1(_05603_),
    .X(_05606_));
 sg13g2_xnor2_1 _15913_ (.Y(_05607_),
    .A(_05535_),
    .B(_05600_));
 sg13g2_xnor2_1 _15914_ (.Y(_05608_),
    .A(_05535_),
    .B(_05601_));
 sg13g2_xnor2_1 _15915_ (.Y(_05609_),
    .A(_05548_),
    .B(_05575_));
 sg13g2_inv_1 _15916_ (.Y(_05610_),
    .A(_05609_));
 sg13g2_xnor2_1 _15917_ (.Y(_05611_),
    .A(_04631_),
    .B(_04643_));
 sg13g2_inv_1 _15918_ (.Y(_05612_),
    .A(_05611_));
 sg13g2_xnor2_1 _15919_ (.Y(_05613_),
    .A(_03962_),
    .B(_04586_));
 sg13g2_inv_1 _15920_ (.Y(_05614_),
    .A(_05613_));
 sg13g2_xnor2_1 _15921_ (.Y(_05615_),
    .A(_05496_),
    .B(_05511_));
 sg13g2_inv_1 _15922_ (.Y(_05617_),
    .A(_05615_));
 sg13g2_xnor2_1 _15923_ (.Y(_05618_),
    .A(_04496_),
    .B(_04497_));
 sg13g2_xnor2_1 _15924_ (.Y(_05619_),
    .A(_04341_),
    .B(_04383_));
 sg13g2_xnor2_1 _15925_ (.Y(_05620_),
    .A(_05212_),
    .B(_05214_));
 sg13g2_nand2b_1 _15926_ (.Y(_05621_),
    .B(_05620_),
    .A_N(_05619_));
 sg13g2_xnor2_1 _15927_ (.Y(_05622_),
    .A(_05427_),
    .B(_05428_));
 sg13g2_inv_1 _15928_ (.Y(_05623_),
    .A(_05622_));
 sg13g2_nor2_1 _15929_ (.A(_05618_),
    .B(_05621_),
    .Y(_05624_));
 sg13g2_nor2_1 _15930_ (.A(_05622_),
    .B(_05624_),
    .Y(_05625_));
 sg13g2_a221oi_1 _15931_ (.B2(_05621_),
    .C1(_05625_),
    .B1(_05618_),
    .A1(_05613_),
    .Y(_05626_),
    .A2(_05615_));
 sg13g2_a221oi_1 _15932_ (.B2(_05617_),
    .C1(_05626_),
    .B1(_05614_),
    .A1(_05610_),
    .Y(_05628_),
    .A2(_05612_));
 sg13g2_a21oi_1 _15933_ (.A1(_05609_),
    .A2(_05611_),
    .Y(_05629_),
    .B1(_05628_));
 sg13g2_xor2_1 _15934_ (.B(_05591_),
    .A(_05590_),
    .X(_05630_));
 sg13g2_inv_1 _15935_ (.Y(_05631_),
    .A(_05630_));
 sg13g2_xnor2_1 _15936_ (.Y(_05632_),
    .A(_04663_),
    .B(_04665_));
 sg13g2_nand2_1 _15937_ (.Y(_05633_),
    .A(_05630_),
    .B(_05632_));
 sg13g2_nor2_1 _15938_ (.A(_05630_),
    .B(_05632_),
    .Y(_05634_));
 sg13g2_a21oi_1 _15939_ (.A1(_05629_),
    .A2(_05633_),
    .Y(_05635_),
    .B1(_05634_));
 sg13g2_o21ai_1 _15940_ (.B1(_04672_),
    .Y(_05636_),
    .A1(_05607_),
    .A2(_05635_));
 sg13g2_a22oi_1 _15941_ (.Y(_05637_),
    .B1(_05607_),
    .B2(_05635_),
    .A2(_05606_),
    .A1(_04675_));
 sg13g2_a21o_2 _15942_ (.A2(_05607_),
    .A1(_04672_),
    .B1(_05635_),
    .X(_05639_));
 sg13g2_a22oi_1 _15943_ (.Y(_05640_),
    .B1(_05608_),
    .B2(_04671_),
    .A2(_05604_),
    .A1(_04676_));
 sg13g2_a22oi_1 _15944_ (.Y(_05641_),
    .B1(_05636_),
    .B2(_05637_),
    .A2(_05604_),
    .A1(_04676_));
 sg13g2_a22oi_1 _15945_ (.Y(_05642_),
    .B1(_05639_),
    .B2(_05640_),
    .A2(_05606_),
    .A1(_04675_));
 sg13g2_a221oi_1 _15946_ (.B2(_05640_),
    .C1(_04672_),
    .B1(_05639_),
    .A1(_04675_),
    .Y(_05643_),
    .A2(_05606_));
 sg13g2_a221oi_1 _15947_ (.B2(_05640_),
    .C1(_04671_),
    .B1(_05639_),
    .A1(_04675_),
    .Y(_05644_),
    .A2(_05606_));
 sg13g2_a21oi_1 _15948_ (.A1(_05607_),
    .A2(_05641_),
    .Y(_05645_),
    .B1(_05643_));
 sg13g2_o21ai_1 _15949_ (.B1(_03766_),
    .Y(_05646_),
    .A1(net2176),
    .A2(net2173));
 sg13g2_or4_1 _15950_ (.A(_03359_),
    .B(net2175),
    .C(_03768_),
    .D(net2174),
    .X(_05647_));
 sg13g2_o21ai_1 _15951_ (.B1(_03767_),
    .Y(_05648_),
    .A1(net2175),
    .A2(net2173));
 sg13g2_or3_1 _15952_ (.A(net2175),
    .B(_03769_),
    .C(net2173),
    .X(_05650_));
 sg13g2_nand2_1 _15953_ (.Y(_05651_),
    .A(_05648_),
    .B(_05650_));
 sg13g2_a221oi_1 _15954_ (.B2(_05650_),
    .C1(_05644_),
    .B1(_05648_),
    .A1(_05608_),
    .Y(_05652_),
    .A2(_05641_));
 sg13g2_a221oi_1 _15955_ (.B2(_03765_),
    .C1(_03798_),
    .B1(_03800_),
    .A1(_03756_),
    .Y(_05653_),
    .A2(_03794_));
 sg13g2_o21ai_1 _15956_ (.B1(_03795_),
    .Y(_05654_),
    .A1(net2176),
    .A2(net2174));
 sg13g2_nor3_1 _15957_ (.A(net2175),
    .B(_03791_),
    .C(net2173),
    .Y(_05655_));
 sg13g2_or3_1 _15958_ (.A(net2175),
    .B(_03791_),
    .C(net2173),
    .X(_05656_));
 sg13g2_nand2_1 _15959_ (.Y(_05657_),
    .A(_05654_),
    .B(_05656_));
 sg13g2_a221oi_1 _15960_ (.B2(_05637_),
    .C1(_05630_),
    .B1(_05636_),
    .A1(_04676_),
    .Y(_05658_),
    .A2(_05604_));
 sg13g2_a221oi_1 _15961_ (.B2(_05640_),
    .C1(_05632_),
    .B1(_05639_),
    .A1(_04675_),
    .Y(_05659_),
    .A2(_05606_));
 sg13g2_a221oi_1 _15962_ (.B2(_05637_),
    .C1(_05631_),
    .B1(_05636_),
    .A1(_04676_),
    .Y(_05661_),
    .A2(_05604_));
 sg13g2_nor2_1 _15963_ (.A(_05659_),
    .B(_05661_),
    .Y(_05662_));
 sg13g2_a221oi_1 _15964_ (.B2(_05656_),
    .C1(_05658_),
    .B1(_05654_),
    .A1(_05632_),
    .Y(_05663_),
    .A2(_05642_));
 sg13g2_nor2_1 _15965_ (.A(_05652_),
    .B(_05663_),
    .Y(_05664_));
 sg13g2_a221oi_1 _15966_ (.B2(_05647_),
    .C1(_05643_),
    .B1(_05646_),
    .A1(_05607_),
    .Y(_05665_),
    .A2(_05641_));
 sg13g2_nor4_1 _15967_ (.A(_05653_),
    .B(_05655_),
    .C(_05659_),
    .D(_05661_),
    .Y(_05666_));
 sg13g2_nor4_2 _15968_ (.A(_05652_),
    .B(_05663_),
    .C(_05665_),
    .Y(_05667_),
    .D(_05666_));
 sg13g2_mux2_1 _15969_ (.A0(_05609_),
    .A1(_05612_),
    .S(_05642_),
    .X(_05668_));
 sg13g2_mux2_1 _15970_ (.A0(_05610_),
    .A1(_05611_),
    .S(_05642_),
    .X(_05669_));
 sg13g2_or3_1 _15971_ (.A(net2175),
    .B(_03771_),
    .C(net2173),
    .X(_05670_));
 sg13g2_o21ai_1 _15972_ (.B1(_05670_),
    .Y(_05672_),
    .A1(_03789_),
    .A2(_03802_));
 sg13g2_mux2_1 _15973_ (.A0(_03789_),
    .A1(_03771_),
    .S(_03802_),
    .X(_05673_));
 sg13g2_mux2_1 _15974_ (.A0(_05613_),
    .A1(_05617_),
    .S(_05641_),
    .X(_05674_));
 sg13g2_mux2_1 _15975_ (.A0(_05614_),
    .A1(_05615_),
    .S(_05641_),
    .X(_05675_));
 sg13g2_or3_1 _15976_ (.A(net2175),
    .B(_03783_),
    .C(net2173),
    .X(_05676_));
 sg13g2_o21ai_1 _15977_ (.B1(_05676_),
    .Y(_05677_),
    .A1(_03781_),
    .A2(_03802_));
 sg13g2_mux2_1 _15978_ (.A0(_03781_),
    .A1(_03783_),
    .S(_03802_),
    .X(_05678_));
 sg13g2_a22oi_1 _15979_ (.Y(_05679_),
    .B1(_05675_),
    .B2(_05677_),
    .A2(_05672_),
    .A1(_05668_));
 sg13g2_nand2_1 _15980_ (.Y(_05680_),
    .A(_05669_),
    .B(_05673_));
 sg13g2_a22oi_1 _15981_ (.Y(_05681_),
    .B1(_05674_),
    .B2(_05678_),
    .A2(_05673_),
    .A1(_05669_));
 sg13g2_and3_1 _15982_ (.X(_05683_),
    .A(_05667_),
    .B(_05679_),
    .C(_05681_));
 sg13g2_nor3_1 _15983_ (.A(net2176),
    .B(_03772_),
    .C(net2174),
    .Y(_05684_));
 sg13g2_or3_1 _15984_ (.A(net2176),
    .B(_03772_),
    .C(net2174),
    .X(_05685_));
 sg13g2_a221oi_1 _15985_ (.B2(_03765_),
    .C1(_03798_),
    .B1(_03800_),
    .A1(_03654_),
    .Y(_05686_),
    .A2(_03773_));
 sg13g2_o21ai_1 _15986_ (.B1(_03774_),
    .Y(_05687_),
    .A1(net2176),
    .A2(net2174));
 sg13g2_nand2_1 _15987_ (.Y(_05688_),
    .A(_05685_),
    .B(_05687_));
 sg13g2_a221oi_1 _15988_ (.B2(_05637_),
    .C1(_05622_),
    .B1(_05636_),
    .A1(_04676_),
    .Y(_05689_),
    .A2(_05604_));
 sg13g2_a221oi_1 _15989_ (.B2(_05640_),
    .C1(_05618_),
    .B1(_05639_),
    .A1(_04675_),
    .Y(_05690_),
    .A2(_05606_));
 sg13g2_a221oi_1 _15990_ (.B2(_05637_),
    .C1(_05623_),
    .B1(_05636_),
    .A1(_04676_),
    .Y(_05691_),
    .A2(_05604_));
 sg13g2_nor2_1 _15991_ (.A(_05689_),
    .B(_05690_),
    .Y(_05692_));
 sg13g2_or4_1 _15992_ (.A(_05684_),
    .B(_05686_),
    .C(_05689_),
    .D(_05690_),
    .X(_05694_));
 sg13g2_a221oi_1 _15993_ (.B2(_05637_),
    .C1(_05620_),
    .B1(_05636_),
    .A1(_04676_),
    .Y(_05695_),
    .A2(_05604_));
 sg13g2_a221oi_1 _15994_ (.B2(_05640_),
    .C1(_05619_),
    .B1(_05639_),
    .A1(_04675_),
    .Y(_05696_),
    .A2(_05606_));
 sg13g2_nor2_1 _15995_ (.A(_05695_),
    .B(_05696_),
    .Y(_05697_));
 sg13g2_or4_1 _15996_ (.A(_03803_),
    .B(_03804_),
    .C(_05695_),
    .D(_05696_),
    .X(_05698_));
 sg13g2_nand2_1 _15997_ (.Y(_05699_),
    .A(_05694_),
    .B(_05698_));
 sg13g2_a221oi_1 _15998_ (.B2(_05687_),
    .C1(_05691_),
    .B1(_05685_),
    .A1(_05618_),
    .Y(_05700_),
    .A2(_05642_));
 sg13g2_a21o_1 _15999_ (.A2(_05698_),
    .A1(_05694_),
    .B1(_05700_),
    .X(_05701_));
 sg13g2_nand4_1 _16000_ (.B(_05679_),
    .C(_05681_),
    .A(_05667_),
    .Y(_05702_),
    .D(_05701_));
 sg13g2_nand3b_1 _16001_ (.B(_05680_),
    .C(_05667_),
    .Y(_05703_),
    .A_N(_05679_));
 sg13g2_nand2b_2 _16002_ (.Y(_05705_),
    .B(_03763_),
    .A_N(_03361_));
 sg13g2_nor2_2 _16003_ (.A(_04676_),
    .B(_05606_),
    .Y(_05706_));
 sg13g2_nor2_1 _16004_ (.A(_05705_),
    .B(_05706_),
    .Y(_05707_));
 sg13g2_or2_1 _16005_ (.X(_05708_),
    .B(_05706_),
    .A(_05705_));
 sg13g2_or2_1 _16006_ (.X(_05709_),
    .B(_05665_),
    .A(_05664_));
 sg13g2_nand4_1 _16007_ (.B(_05703_),
    .C(_05708_),
    .A(_05702_),
    .Y(_05710_),
    .D(_05709_));
 sg13g2_nor2_1 _16008_ (.A(_03805_),
    .B(_05697_),
    .Y(_05711_));
 sg13g2_nor4_1 _16009_ (.A(_05699_),
    .B(_05700_),
    .C(_05707_),
    .D(_05711_),
    .Y(_05712_));
 sg13g2_a22oi_1 _16010_ (.Y(_05713_),
    .B1(_05712_),
    .B2(_05683_),
    .A2(_05706_),
    .A1(_05705_));
 sg13g2_and2_2 _16011_ (.A(_05710_),
    .B(_05713_),
    .X(_05714_));
 sg13g2_inv_2 _16012_ (.Y(_05716_),
    .A(_05714_));
 sg13g2_a21oi_2 _16013_ (.B1(_03805_),
    .Y(_05717_),
    .A2(_05713_),
    .A1(_05710_));
 sg13g2_nand3_1 _16014_ (.B(_05710_),
    .C(_05713_),
    .A(_05697_),
    .Y(_05718_));
 sg13g2_nand2b_1 _16015_ (.Y(_05719_),
    .B(_05718_),
    .A_N(_05717_));
 sg13g2_inv_1 _16016_ (.Y(_05720_),
    .A(_05719_));
 sg13g2_nand2b_1 _16017_ (.Y(_05721_),
    .B(net2616),
    .A_N(net2428));
 sg13g2_nor2_1 _16018_ (.A(net2710),
    .B(net2777),
    .Y(_05722_));
 sg13g2_xnor2_1 _16019_ (.Y(_05723_),
    .A(_05721_),
    .B(_05722_));
 sg13g2_xor2_1 _16020_ (.B(net2643),
    .A(net2593),
    .X(_05724_));
 sg13g2_xor2_1 _16021_ (.B(\net.in[174] ),
    .A(net2527),
    .X(_05725_));
 sg13g2_and2_1 _16022_ (.A(_05724_),
    .B(_05725_),
    .X(_05727_));
 sg13g2_xnor2_1 _16023_ (.Y(_05728_),
    .A(net2688),
    .B(net2770));
 sg13g2_nor3_1 _16024_ (.A(\net.in[34] ),
    .B(_06694_),
    .C(_05728_),
    .Y(_05729_));
 sg13g2_o21ai_1 _16025_ (.B1(_05728_),
    .Y(_05730_),
    .A1(\net.in[34] ),
    .A2(_06694_));
 sg13g2_nor2b_1 _16026_ (.A(_05729_),
    .B_N(_05730_),
    .Y(_05731_));
 sg13g2_xnor2_1 _16027_ (.Y(_05732_),
    .A(_05727_),
    .B(_05731_));
 sg13g2_xor2_1 _16028_ (.B(net2723),
    .A(net2751),
    .X(_05733_));
 sg13g2_nand2b_1 _16029_ (.Y(_05734_),
    .B(net2683),
    .A_N(net2643));
 sg13g2_o21ai_1 _16030_ (.B1(_05734_),
    .Y(_05735_),
    .A1(net2519),
    .A2(net2577));
 sg13g2_a21oi_2 _16031_ (.B1(_05735_),
    .Y(_05736_),
    .A2(net2643),
    .A1(net2177));
 sg13g2_xnor2_1 _16032_ (.Y(_05738_),
    .A(net2307),
    .B(net2358));
 sg13g2_nor2_1 _16033_ (.A(_05736_),
    .B(_05738_),
    .Y(_05739_));
 sg13g2_xnor2_1 _16034_ (.Y(_05740_),
    .A(_05736_),
    .B(_05738_));
 sg13g2_xnor2_1 _16035_ (.Y(_05741_),
    .A(_05733_),
    .B(_05740_));
 sg13g2_nand2_1 _16036_ (.Y(_05742_),
    .A(_05732_),
    .B(_05741_));
 sg13g2_xnor2_1 _16037_ (.Y(_05743_),
    .A(_05732_),
    .B(_05741_));
 sg13g2_nor2_1 _16038_ (.A(net2487),
    .B(net2589),
    .Y(_05744_));
 sg13g2_xnor2_1 _16039_ (.Y(_05745_),
    .A(net2641),
    .B(_05744_));
 sg13g2_nand2b_1 _16040_ (.Y(_05746_),
    .B(\net.in[201] ),
    .A_N(net2374));
 sg13g2_nand2b_1 _16041_ (.Y(_05747_),
    .B(net2374),
    .A_N(net2288));
 sg13g2_nand2b_1 _16042_ (.Y(_05749_),
    .B(net2537),
    .A_N(net2619));
 sg13g2_nand3_1 _16043_ (.B(_05747_),
    .C(_05749_),
    .A(_05746_),
    .Y(_05750_));
 sg13g2_nand4_1 _16044_ (.B(_05746_),
    .C(_05747_),
    .A(_05745_),
    .Y(_05751_),
    .D(_05749_));
 sg13g2_nor2b_1 _16045_ (.A(_05745_),
    .B_N(_05750_),
    .Y(_05752_));
 sg13g2_xor2_1 _16046_ (.B(_05750_),
    .A(_05745_),
    .X(_05753_));
 sg13g2_xnor2_1 _16047_ (.Y(_05754_),
    .A(net2333),
    .B(net2342));
 sg13g2_xnor2_1 _16048_ (.Y(_05755_),
    .A(_05753_),
    .B(_05754_));
 sg13g2_xnor2_1 _16049_ (.Y(_05756_),
    .A(_05743_),
    .B(_05755_));
 sg13g2_nor2_2 _16050_ (.A(net2552),
    .B(net2600),
    .Y(_05757_));
 sg13g2_o21ai_1 _16051_ (.B1(_05757_),
    .Y(_05758_),
    .A1(net2698),
    .A2(net2768));
 sg13g2_a21o_1 _16052_ (.A2(net2767),
    .A1(net2698),
    .B1(_05758_),
    .X(_05760_));
 sg13g2_or2_1 _16053_ (.X(_05761_),
    .B(net2773),
    .A(net2361));
 sg13g2_xor2_1 _16054_ (.B(net2643),
    .A(net2577),
    .X(_05762_));
 sg13g2_nor3_1 _16055_ (.A(_03818_),
    .B(_05761_),
    .C(_05762_),
    .Y(_05763_));
 sg13g2_o21ai_1 _16056_ (.B1(_05762_),
    .Y(_05764_),
    .A1(_03818_),
    .A2(_05761_));
 sg13g2_nand2b_1 _16057_ (.Y(_05765_),
    .B(_05764_),
    .A_N(_05763_));
 sg13g2_xor2_1 _16058_ (.B(_05765_),
    .A(_05760_),
    .X(_05766_));
 sg13g2_nor2b_1 _16059_ (.A(net2236),
    .B_N(net2205),
    .Y(_05767_));
 sg13g2_nor2b_1 _16060_ (.A(net2205),
    .B_N(net2236),
    .Y(_05768_));
 sg13g2_nor2_1 _16061_ (.A(net2379),
    .B(net2374),
    .Y(_05769_));
 sg13g2_nor3_1 _16062_ (.A(_05767_),
    .B(_05768_),
    .C(_05769_),
    .Y(_05771_));
 sg13g2_nor2_1 _16063_ (.A(_05286_),
    .B(net2201),
    .Y(_05772_));
 sg13g2_nor2_1 _16064_ (.A(_05771_),
    .B(_05772_),
    .Y(_05773_));
 sg13g2_a22oi_1 _16065_ (.Y(_05774_),
    .B1(net2363),
    .B2(net2531),
    .A2(\net.in[225] ),
    .A1(_05429_));
 sg13g2_o21ai_1 _16066_ (.B1(_05774_),
    .Y(_05775_),
    .A1(_05429_),
    .A2(\net.in[225] ));
 sg13g2_and2_1 _16067_ (.A(_05773_),
    .B(_05775_),
    .X(_05776_));
 sg13g2_nand2_1 _16068_ (.Y(_05777_),
    .A(_05771_),
    .B(_05772_));
 sg13g2_a21oi_2 _16069_ (.B1(_05773_),
    .Y(_05778_),
    .A2(_05777_),
    .A1(_05775_));
 sg13g2_inv_1 _16070_ (.Y(_05779_),
    .A(_05778_));
 sg13g2_or2_1 _16071_ (.X(_05780_),
    .B(_05777_),
    .A(_05775_));
 sg13g2_o21ai_1 _16072_ (.B1(_05780_),
    .Y(_05782_),
    .A1(_05776_),
    .A2(_05778_));
 sg13g2_nand2b_1 _16073_ (.Y(_05783_),
    .B(_05766_),
    .A_N(_05782_));
 sg13g2_nor2b_1 _16074_ (.A(_05766_),
    .B_N(_05782_),
    .Y(_05784_));
 sg13g2_xor2_1 _16075_ (.B(_05782_),
    .A(_05766_),
    .X(_05785_));
 sg13g2_a21oi_1 _16076_ (.A1(_05517_),
    .A2(_05957_),
    .Y(_05786_),
    .B1(_08421_));
 sg13g2_nand4_1 _16077_ (.B(net2223),
    .C(net2250),
    .A(_05506_),
    .Y(_05787_),
    .D(_05924_));
 sg13g2_nand2_1 _16078_ (.Y(_05788_),
    .A(net2687),
    .B(net2363));
 sg13g2_xor2_1 _16079_ (.B(_05788_),
    .A(_00010_),
    .X(_05789_));
 sg13g2_nand2b_1 _16080_ (.Y(_05790_),
    .B(_05789_),
    .A_N(_05787_));
 sg13g2_nor2b_1 _16081_ (.A(_05789_),
    .B_N(_05787_),
    .Y(_05791_));
 sg13g2_xnor2_1 _16082_ (.Y(_05793_),
    .A(_05787_),
    .B(_05789_));
 sg13g2_xnor2_1 _16083_ (.Y(_05794_),
    .A(_05786_),
    .B(_05793_));
 sg13g2_xnor2_1 _16084_ (.Y(_05795_),
    .A(_05785_),
    .B(_05794_));
 sg13g2_inv_1 _16085_ (.Y(_05796_),
    .A(_05795_));
 sg13g2_nand2_1 _16086_ (.Y(_05797_),
    .A(_05756_),
    .B(_05796_));
 sg13g2_xor2_1 _16087_ (.B(_05795_),
    .A(_05756_),
    .X(_05798_));
 sg13g2_xnor2_1 _16088_ (.Y(_05799_),
    .A(_05723_),
    .B(_05798_));
 sg13g2_xor2_1 _16089_ (.B(net2350),
    .A(net2339),
    .X(_05800_));
 sg13g2_nor2_1 _16090_ (.A(net2401),
    .B(net2600),
    .Y(_05801_));
 sg13g2_xnor2_1 _16091_ (.Y(_05802_),
    .A(_05800_),
    .B(_05801_));
 sg13g2_nor2_1 _16092_ (.A(net2428),
    .B(net2802),
    .Y(_05804_));
 sg13g2_xnor2_1 _16093_ (.Y(_05805_),
    .A(net2346),
    .B(_05804_));
 sg13g2_xnor2_1 _16094_ (.Y(_05806_),
    .A(net2648),
    .B(_00009_));
 sg13g2_xnor2_1 _16095_ (.Y(_05807_),
    .A(net2346),
    .B(_05806_));
 sg13g2_nand2_1 _16096_ (.Y(_05808_),
    .A(_05805_),
    .B(_05807_));
 sg13g2_nor2_1 _16097_ (.A(_05805_),
    .B(_05807_),
    .Y(_05809_));
 sg13g2_xor2_1 _16098_ (.B(_05806_),
    .A(_05804_),
    .X(_05810_));
 sg13g2_xnor2_1 _16099_ (.Y(_05811_),
    .A(_05802_),
    .B(_05810_));
 sg13g2_xor2_1 _16100_ (.B(net2318),
    .A(\net.in[209] ),
    .X(_05812_));
 sg13g2_xor2_1 _16101_ (.B(net2556),
    .A(net2323),
    .X(_05813_));
 sg13g2_xnor2_1 _16102_ (.Y(_05815_),
    .A(_05812_),
    .B(_05813_));
 sg13g2_xnor2_1 _16103_ (.Y(_05816_),
    .A(net2692),
    .B(net2650));
 sg13g2_xnor2_1 _16104_ (.Y(_05817_),
    .A(net2401),
    .B(net2708));
 sg13g2_xnor2_1 _16105_ (.Y(_05818_),
    .A(net2298),
    .B(net2290));
 sg13g2_and3_1 _16106_ (.X(_05819_),
    .A(_05816_),
    .B(_05817_),
    .C(_05818_));
 sg13g2_inv_1 _16107_ (.Y(_05820_),
    .A(_05819_));
 sg13g2_a21oi_1 _16108_ (.A1(_05816_),
    .A2(_05817_),
    .Y(_05821_),
    .B1(_05818_));
 sg13g2_nand2b_1 _16109_ (.Y(_05822_),
    .B(_05819_),
    .A_N(_05815_));
 sg13g2_o21ai_1 _16110_ (.B1(_05820_),
    .Y(_05823_),
    .A1(_05815_),
    .A2(_05821_));
 sg13g2_a21o_1 _16111_ (.A2(_05821_),
    .A1(_05815_),
    .B1(_05823_),
    .X(_05824_));
 sg13g2_nor2_1 _16112_ (.A(net2182),
    .B(net2504),
    .Y(_05826_));
 sg13g2_xnor2_1 _16113_ (.Y(_05827_),
    .A(net2573),
    .B(net2641));
 sg13g2_inv_1 _16114_ (.Y(_05828_),
    .A(_05827_));
 sg13g2_nand2b_1 _16115_ (.Y(_05829_),
    .B(net2472),
    .A_N(net2540));
 sg13g2_nor2_2 _16116_ (.A(net2654),
    .B(_05682_),
    .Y(_05830_));
 sg13g2_xnor2_1 _16117_ (.Y(_05831_),
    .A(_05829_),
    .B(_05830_));
 sg13g2_nand2_1 _16118_ (.Y(_05832_),
    .A(_05828_),
    .B(_05831_));
 sg13g2_xnor2_1 _16119_ (.Y(_05833_),
    .A(_05827_),
    .B(_05831_));
 sg13g2_xnor2_1 _16120_ (.Y(_05834_),
    .A(_05826_),
    .B(_05833_));
 sg13g2_a21oi_1 _16121_ (.A1(_05822_),
    .A2(_05824_),
    .Y(_05835_),
    .B1(_05834_));
 sg13g2_nand3_1 _16122_ (.B(_05824_),
    .C(_05834_),
    .A(_05822_),
    .Y(_05837_));
 sg13g2_nor2b_1 _16123_ (.A(_05835_),
    .B_N(_05837_),
    .Y(_05838_));
 sg13g2_xor2_1 _16124_ (.B(_05838_),
    .A(_05811_),
    .X(_05839_));
 sg13g2_nor2_1 _16125_ (.A(net2390),
    .B(net2556),
    .Y(_05840_));
 sg13g2_nor2_1 _16126_ (.A(net2261),
    .B(_05264_),
    .Y(_05841_));
 sg13g2_xnor2_1 _16127_ (.Y(_05842_),
    .A(_05840_),
    .B(_05841_));
 sg13g2_a22oi_1 _16128_ (.Y(_05843_),
    .B1(net2395),
    .B2(net2272),
    .A2(_05913_),
    .A1(net2536));
 sg13g2_xor2_1 _16129_ (.B(net2563),
    .A(net2637),
    .X(_05844_));
 sg13g2_nand2_1 _16130_ (.Y(_05845_),
    .A(_05843_),
    .B(_05844_));
 sg13g2_or2_1 _16131_ (.X(_05846_),
    .B(_05844_),
    .A(_05843_));
 sg13g2_nand2_1 _16132_ (.Y(_05848_),
    .A(_05845_),
    .B(_05846_));
 sg13g2_xor2_1 _16133_ (.B(_05848_),
    .A(_05842_),
    .X(_05849_));
 sg13g2_xnor2_1 _16134_ (.Y(_05850_),
    .A(net2383),
    .B(net2330));
 sg13g2_nand2b_2 _16135_ (.Y(_05851_),
    .B(net2201),
    .A_N(net2303));
 sg13g2_nor2_1 _16136_ (.A(\net.in[176] ),
    .B(\net.in[18] ),
    .Y(_05852_));
 sg13g2_xnor2_1 _16137_ (.Y(_05853_),
    .A(_05851_),
    .B(_05852_));
 sg13g2_nor2b_1 _16138_ (.A(net2531),
    .B_N(net2326),
    .Y(_05854_));
 sg13g2_xor2_1 _16139_ (.B(net2773),
    .A(\net.in[65] ),
    .X(_05855_));
 sg13g2_xnor2_1 _16140_ (.Y(_05856_),
    .A(_05854_),
    .B(_05855_));
 sg13g2_nor2_1 _16141_ (.A(_05853_),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_nand2_1 _16142_ (.Y(_05859_),
    .A(_05853_),
    .B(_05856_));
 sg13g2_xor2_1 _16143_ (.B(_05856_),
    .A(_05853_),
    .X(_05860_));
 sg13g2_xnor2_1 _16144_ (.Y(_05861_),
    .A(_05850_),
    .B(_05860_));
 sg13g2_xor2_1 _16145_ (.B(net2424),
    .A(net2333),
    .X(_05862_));
 sg13g2_xnor2_1 _16146_ (.Y(_05863_),
    .A(net2486),
    .B(net2436));
 sg13g2_nor2b_2 _16147_ (.A(net2554),
    .B_N(net2573),
    .Y(_05864_));
 sg13g2_nand2_1 _16148_ (.Y(_05865_),
    .A(_05863_),
    .B(_05864_));
 sg13g2_xnor2_1 _16149_ (.Y(_05866_),
    .A(_05863_),
    .B(_05864_));
 sg13g2_xor2_1 _16150_ (.B(_05866_),
    .A(_05862_),
    .X(_05867_));
 sg13g2_nand2_1 _16151_ (.Y(_05868_),
    .A(_05861_),
    .B(_05867_));
 sg13g2_nor2_1 _16152_ (.A(_05861_),
    .B(_05867_),
    .Y(_05870_));
 sg13g2_xnor2_1 _16153_ (.Y(_05871_),
    .A(_05861_),
    .B(_05867_));
 sg13g2_o21ai_1 _16154_ (.B1(_05868_),
    .Y(_05872_),
    .A1(_05849_),
    .A2(_05870_));
 sg13g2_xnor2_1 _16155_ (.Y(_05873_),
    .A(_05849_),
    .B(_05871_));
 sg13g2_xor2_1 _16156_ (.B(net2640),
    .A(net2648),
    .X(_05874_));
 sg13g2_xnor2_1 _16157_ (.Y(_05875_),
    .A(net2599),
    .B(_05874_));
 sg13g2_nor2_1 _16158_ (.A(_05363_),
    .B(net2598),
    .Y(_05876_));
 sg13g2_nor2b_1 _16159_ (.A(net2383),
    .B_N(net2598),
    .Y(_05877_));
 sg13g2_nor2b_1 _16160_ (.A(net2688),
    .B_N(net2649),
    .Y(_05878_));
 sg13g2_nor3_2 _16161_ (.A(_05876_),
    .B(_05877_),
    .C(_05878_),
    .Y(_05879_));
 sg13g2_xnor2_1 _16162_ (.Y(_05881_),
    .A(net2390),
    .B(net2401));
 sg13g2_xnor2_1 _16163_ (.Y(_05882_),
    .A(net2523),
    .B(net2648));
 sg13g2_xnor2_1 _16164_ (.Y(_05883_),
    .A(_05881_),
    .B(_05882_));
 sg13g2_nand2b_1 _16165_ (.Y(_05884_),
    .B(_05883_),
    .A_N(_05879_));
 sg13g2_nor2b_1 _16166_ (.A(_05883_),
    .B_N(_05879_),
    .Y(_05885_));
 sg13g2_xnor2_1 _16167_ (.Y(_05886_),
    .A(_05879_),
    .B(_05883_));
 sg13g2_xnor2_1 _16168_ (.Y(_05887_),
    .A(_05875_),
    .B(_05886_));
 sg13g2_nand2_1 _16169_ (.Y(_05888_),
    .A(net2486),
    .B(net2182));
 sg13g2_o21ai_1 _16170_ (.B1(_05888_),
    .Y(_05889_),
    .A1(net2225),
    .A2(net2563));
 sg13g2_inv_1 _16171_ (.Y(_05890_),
    .A(_05889_));
 sg13g2_xor2_1 _16172_ (.B(net2767),
    .A(net2507),
    .X(_05892_));
 sg13g2_nor2_1 _16173_ (.A(net2692),
    .B(net2601),
    .Y(_05893_));
 sg13g2_nor2_1 _16174_ (.A(net2683),
    .B(net2650),
    .Y(_05894_));
 sg13g2_xnor2_1 _16175_ (.Y(_05895_),
    .A(_05893_),
    .B(_05894_));
 sg13g2_nor2_1 _16176_ (.A(_05892_),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_xor2_1 _16177_ (.B(_05895_),
    .A(_05892_),
    .X(_05897_));
 sg13g2_xnor2_1 _16178_ (.Y(_05898_),
    .A(_05889_),
    .B(_05897_));
 sg13g2_o21ai_1 _16179_ (.B1(_05418_),
    .Y(_05899_),
    .A1(net2797),
    .A2(net2314));
 sg13g2_xnor2_1 _16180_ (.Y(_05900_),
    .A(net2298),
    .B(net2411));
 sg13g2_nand2_1 _16181_ (.Y(_05901_),
    .A(net2643),
    .B(net2317));
 sg13g2_xor2_1 _16182_ (.B(net2208),
    .A(net2275),
    .X(_05903_));
 sg13g2_xnor2_1 _16183_ (.Y(_05904_),
    .A(_05901_),
    .B(_05903_));
 sg13g2_nand2_1 _16184_ (.Y(_05905_),
    .A(_05900_),
    .B(_05904_));
 sg13g2_nor2_1 _16185_ (.A(_05900_),
    .B(_05904_),
    .Y(_05906_));
 sg13g2_xor2_1 _16186_ (.B(_05904_),
    .A(_05900_),
    .X(_05907_));
 sg13g2_xnor2_1 _16187_ (.Y(_05908_),
    .A(_05899_),
    .B(_05907_));
 sg13g2_nor2_1 _16188_ (.A(_05898_),
    .B(_05908_),
    .Y(_05909_));
 sg13g2_nand2_1 _16189_ (.Y(_05910_),
    .A(_05898_),
    .B(_05908_));
 sg13g2_o21ai_1 _16190_ (.B1(_05910_),
    .Y(_05911_),
    .A1(_05887_),
    .A2(_05909_));
 sg13g2_xor2_1 _16191_ (.B(_05908_),
    .A(_05898_),
    .X(_05912_));
 sg13g2_xnor2_1 _16192_ (.Y(_05914_),
    .A(_05887_),
    .B(_05912_));
 sg13g2_nand2_1 _16193_ (.Y(_05915_),
    .A(_05873_),
    .B(_05914_));
 sg13g2_or2_1 _16194_ (.X(_05916_),
    .B(_05914_),
    .A(_05873_));
 sg13g2_nand2_1 _16195_ (.Y(_05917_),
    .A(_05915_),
    .B(_05916_));
 sg13g2_xnor2_1 _16196_ (.Y(_05918_),
    .A(_05839_),
    .B(_05917_));
 sg13g2_and2_1 _16197_ (.A(_05799_),
    .B(_05918_),
    .X(_05919_));
 sg13g2_xor2_1 _16198_ (.B(_05918_),
    .A(_05799_),
    .X(_05920_));
 sg13g2_nor2b_1 _16199_ (.A(\net.in[80] ),
    .B_N(net2540),
    .Y(_05921_));
 sg13g2_xnor2_1 _16200_ (.Y(_05922_),
    .A(net2351),
    .B(net2589));
 sg13g2_xnor2_1 _16201_ (.Y(_05923_),
    .A(_05921_),
    .B(_05922_));
 sg13g2_nand2b_1 _16202_ (.Y(_05925_),
    .B(net2472),
    .A_N(net2536));
 sg13g2_nor2_1 _16203_ (.A(_05693_),
    .B(net2650),
    .Y(_05926_));
 sg13g2_xnor2_1 _16204_ (.Y(_05927_),
    .A(_05925_),
    .B(_05926_));
 sg13g2_nand2b_1 _16205_ (.Y(_05928_),
    .B(net2678),
    .A_N(net2342));
 sg13g2_xnor2_1 _16206_ (.Y(_05929_),
    .A(_00577_),
    .B(_05928_));
 sg13g2_nand2_1 _16207_ (.Y(_05930_),
    .A(_05927_),
    .B(_05929_));
 sg13g2_nor2_1 _16208_ (.A(_05927_),
    .B(_05929_),
    .Y(_05931_));
 sg13g2_xor2_1 _16209_ (.B(_05929_),
    .A(_05927_),
    .X(_05932_));
 sg13g2_xnor2_1 _16210_ (.Y(_05933_),
    .A(_05923_),
    .B(_05932_));
 sg13g2_nand2b_1 _16211_ (.Y(_05934_),
    .B(net2383),
    .A_N(net2307));
 sg13g2_xnor2_1 _16212_ (.Y(_05936_),
    .A(_04815_),
    .B(_05934_));
 sg13g2_nor3_1 _16213_ (.A(_05044_),
    .B(net2500),
    .C(_05936_),
    .Y(_05937_));
 sg13g2_o21ai_1 _16214_ (.B1(_05936_),
    .Y(_05938_),
    .A1(_05044_),
    .A2(net2500));
 sg13g2_nand2b_1 _16215_ (.Y(_05939_),
    .B(_05938_),
    .A_N(_05937_));
 sg13g2_nor2_1 _16216_ (.A(net2523),
    .B(net2556),
    .Y(_05940_));
 sg13g2_xnor2_1 _16217_ (.Y(_05941_),
    .A(_05724_),
    .B(_05940_));
 sg13g2_xnor2_1 _16218_ (.Y(_05942_),
    .A(_05939_),
    .B(_05941_));
 sg13g2_nor2_1 _16219_ (.A(_05933_),
    .B(_05942_),
    .Y(_05943_));
 sg13g2_nand2_1 _16220_ (.Y(_05944_),
    .A(_00006_),
    .B(_05816_));
 sg13g2_nand2_1 _16221_ (.Y(_05945_),
    .A(_00006_),
    .B(_05881_));
 sg13g2_nor2_1 _16222_ (.A(net2182),
    .B(net2590),
    .Y(_05947_));
 sg13g2_nor2_1 _16223_ (.A(net2616),
    .B(_05979_),
    .Y(_05948_));
 sg13g2_xnor2_1 _16224_ (.Y(_05949_),
    .A(_05947_),
    .B(_05948_));
 sg13g2_nand2_1 _16225_ (.Y(_05950_),
    .A(_05945_),
    .B(_05949_));
 sg13g2_xnor2_1 _16226_ (.Y(_05951_),
    .A(_05945_),
    .B(_05949_));
 sg13g2_xnor2_1 _16227_ (.Y(_05952_),
    .A(_05944_),
    .B(_05951_));
 sg13g2_nor2_1 _16228_ (.A(_05943_),
    .B(_05952_),
    .Y(_05953_));
 sg13g2_a21oi_1 _16229_ (.A1(_05933_),
    .A2(_05942_),
    .Y(_05954_),
    .B1(_05953_));
 sg13g2_xnor2_1 _16230_ (.Y(_05955_),
    .A(_05933_),
    .B(_05942_));
 sg13g2_xnor2_1 _16231_ (.Y(_05956_),
    .A(_05952_),
    .B(_05955_));
 sg13g2_a22oi_1 _16232_ (.Y(_05958_),
    .B1(_06001_),
    .B2(net2663),
    .A2(net2573),
    .A1(net2326));
 sg13g2_o21ai_1 _16233_ (.B1(_05958_),
    .Y(_05959_),
    .A1(net2663),
    .A2(_06001_));
 sg13g2_nor2b_1 _16234_ (.A(net2266),
    .B_N(net2201),
    .Y(_05960_));
 sg13g2_nor2b_1 _16235_ (.A(net2201),
    .B_N(net2266),
    .Y(_05961_));
 sg13g2_nor2b_1 _16236_ (.A(net2755),
    .B_N(net2342),
    .Y(_05962_));
 sg13g2_nor3_2 _16237_ (.A(_05960_),
    .B(_05961_),
    .C(_05962_),
    .Y(_05963_));
 sg13g2_o21ai_1 _16238_ (.B1(_05963_),
    .Y(_05964_),
    .A1(net2540),
    .A2(_01230_));
 sg13g2_or3_1 _16239_ (.A(net2541),
    .B(_01230_),
    .C(_05963_),
    .X(_05965_));
 sg13g2_and2_1 _16240_ (.A(_05964_),
    .B(_05965_),
    .X(_05966_));
 sg13g2_xnor2_1 _16241_ (.Y(_05967_),
    .A(_05959_),
    .B(_05966_));
 sg13g2_xnor2_1 _16242_ (.Y(_05969_),
    .A(\net.in[75] ),
    .B(net2780));
 sg13g2_xnor2_1 _16243_ (.Y(_05970_),
    .A(net2641),
    .B(_05969_));
 sg13g2_nand2_1 _16244_ (.Y(_05971_),
    .A(_04750_),
    .B(_05970_));
 sg13g2_xor2_1 _16245_ (.B(_05970_),
    .A(_04750_),
    .X(_05972_));
 sg13g2_xor2_1 _16246_ (.B(net2281),
    .A(net2288),
    .X(_05973_));
 sg13g2_xnor2_1 _16247_ (.Y(_05974_),
    .A(_05972_),
    .B(_05973_));
 sg13g2_o21ai_1 _16248_ (.B1(_02823_),
    .Y(_05975_),
    .A1(net2741),
    .A2(_05660_));
 sg13g2_a21oi_2 _16249_ (.B1(_05975_),
    .Y(_05976_),
    .A2(_05660_),
    .A1(net2741));
 sg13g2_nand2b_1 _16250_ (.Y(_05977_),
    .B(net2784),
    .A_N(net2432));
 sg13g2_nand2b_1 _16251_ (.Y(_05978_),
    .B(net2767),
    .A_N(net2293));
 sg13g2_xnor2_1 _16252_ (.Y(_05980_),
    .A(net2583),
    .B(net2619));
 sg13g2_and3_1 _16253_ (.X(_05981_),
    .A(_05977_),
    .B(_05978_),
    .C(_05980_));
 sg13g2_a21oi_1 _16254_ (.A1(_05977_),
    .A2(_05978_),
    .Y(_05982_),
    .B1(_05980_));
 sg13g2_inv_1 _16255_ (.Y(_05983_),
    .A(_05982_));
 sg13g2_nor2_1 _16256_ (.A(_05981_),
    .B(_05982_),
    .Y(_05984_));
 sg13g2_xnor2_1 _16257_ (.Y(_05985_),
    .A(_05976_),
    .B(_05984_));
 sg13g2_nor2b_1 _16258_ (.A(_05985_),
    .B_N(_05974_),
    .Y(_05986_));
 sg13g2_nand2b_1 _16259_ (.Y(_05987_),
    .B(_05985_),
    .A_N(_05974_));
 sg13g2_xnor2_1 _16260_ (.Y(_05988_),
    .A(_05974_),
    .B(_05985_));
 sg13g2_o21ai_1 _16261_ (.B1(_05987_),
    .Y(_05989_),
    .A1(_05967_),
    .A2(_05986_));
 sg13g2_xnor2_1 _16262_ (.Y(_05991_),
    .A(_05967_),
    .B(_05988_));
 sg13g2_xor2_1 _16263_ (.B(net2476),
    .A(net2753),
    .X(_05992_));
 sg13g2_nor2_1 _16264_ (.A(net2432),
    .B(net2379),
    .Y(_05993_));
 sg13g2_nand2b_1 _16265_ (.Y(_05994_),
    .B(net2199),
    .A_N(net2257));
 sg13g2_xnor2_1 _16266_ (.Y(_05995_),
    .A(_05993_),
    .B(_05994_));
 sg13g2_nor2_1 _16267_ (.A(_05992_),
    .B(_05995_),
    .Y(_05996_));
 sg13g2_nand2_1 _16268_ (.Y(_05997_),
    .A(_05992_),
    .B(_05995_));
 sg13g2_nor2b_1 _16269_ (.A(_05996_),
    .B_N(_05997_),
    .Y(_05998_));
 sg13g2_nor2b_1 _16270_ (.A(net2198),
    .B_N(net2254),
    .Y(_05999_));
 sg13g2_nor2b_1 _16271_ (.A(net2500),
    .B_N(net2221),
    .Y(_06000_));
 sg13g2_xnor2_1 _16272_ (.Y(_06002_),
    .A(_05999_),
    .B(_06000_));
 sg13g2_xnor2_1 _16273_ (.Y(_06003_),
    .A(_05998_),
    .B(_06002_));
 sg13g2_a22oi_1 _16274_ (.Y(_06004_),
    .B1(_06045_),
    .B2(net2666),
    .A2(net2760),
    .A1(_05077_));
 sg13g2_o21ai_1 _16275_ (.B1(_06004_),
    .Y(_06005_),
    .A1(net2666),
    .A2(_06045_));
 sg13g2_nor2_2 _16276_ (.A(net2736),
    .B(net2621),
    .Y(_06006_));
 sg13g2_nor2_1 _16277_ (.A(net2795),
    .B(net2650),
    .Y(_06007_));
 sg13g2_xnor2_1 _16278_ (.Y(_06008_),
    .A(_06006_),
    .B(_06007_));
 sg13g2_nand2b_1 _16279_ (.Y(_06009_),
    .B(net2523),
    .A_N(net2383));
 sg13g2_xnor2_1 _16280_ (.Y(_06010_),
    .A(net2508),
    .B(\net.in[49] ));
 sg13g2_xnor2_1 _16281_ (.Y(_06011_),
    .A(_06009_),
    .B(_06010_));
 sg13g2_nor2_1 _16282_ (.A(_06008_),
    .B(_06011_),
    .Y(_06013_));
 sg13g2_nand2_1 _16283_ (.Y(_06014_),
    .A(_06008_),
    .B(_06011_));
 sg13g2_xnor2_1 _16284_ (.Y(_06015_),
    .A(_06008_),
    .B(_06011_));
 sg13g2_o21ai_1 _16285_ (.B1(_06014_),
    .Y(_06016_),
    .A1(_06005_),
    .A2(_06013_));
 sg13g2_xnor2_1 _16286_ (.Y(_06017_),
    .A(_06005_),
    .B(_06015_));
 sg13g2_xnor2_1 _16287_ (.Y(_06018_),
    .A(net2330),
    .B(net2701));
 sg13g2_xnor2_1 _16288_ (.Y(_06019_),
    .A(net2772),
    .B(_06018_));
 sg13g2_xor2_1 _16289_ (.B(net2198),
    .A(net2784),
    .X(_06020_));
 sg13g2_nand2_1 _16290_ (.Y(_06021_),
    .A(_06019_),
    .B(_06020_));
 sg13g2_xor2_1 _16291_ (.B(_06020_),
    .A(_06019_),
    .X(_06022_));
 sg13g2_nor2_1 _16292_ (.A(net2473),
    .B(net2575),
    .Y(_06024_));
 sg13g2_a21oi_2 _16293_ (.B1(_06024_),
    .Y(_06025_),
    .A2(_06177_),
    .A1(net2473));
 sg13g2_xnor2_1 _16294_ (.Y(_06026_),
    .A(_06022_),
    .B(_06025_));
 sg13g2_inv_1 _16295_ (.Y(_06027_),
    .A(_06026_));
 sg13g2_nand2_1 _16296_ (.Y(_06028_),
    .A(_06017_),
    .B(_06027_));
 sg13g2_xor2_1 _16297_ (.B(_06026_),
    .A(_06017_),
    .X(_06029_));
 sg13g2_xnor2_1 _16298_ (.Y(_06030_),
    .A(_06003_),
    .B(_06029_));
 sg13g2_nand2_1 _16299_ (.Y(_06031_),
    .A(_05991_),
    .B(_06030_));
 sg13g2_or2_1 _16300_ (.X(_06032_),
    .B(_06030_),
    .A(_05991_));
 sg13g2_xor2_1 _16301_ (.B(_06030_),
    .A(_05991_),
    .X(_06033_));
 sg13g2_xnor2_1 _16302_ (.Y(_06035_),
    .A(_05956_),
    .B(_06033_));
 sg13g2_nor2_1 _16303_ (.A(net2540),
    .B(net2495),
    .Y(_06036_));
 sg13g2_xnor2_1 _16304_ (.Y(_06037_),
    .A(net2191),
    .B(net2254));
 sg13g2_xnor2_1 _16305_ (.Y(_06038_),
    .A(net2199),
    .B(net2321));
 sg13g2_nand2_1 _16306_ (.Y(_06039_),
    .A(_06037_),
    .B(_06038_));
 sg13g2_nor2_1 _16307_ (.A(_06037_),
    .B(_06038_),
    .Y(_06040_));
 sg13g2_xnor2_1 _16308_ (.Y(_06041_),
    .A(_06037_),
    .B(_06038_));
 sg13g2_xor2_1 _16309_ (.B(_06041_),
    .A(_06036_),
    .X(_06042_));
 sg13g2_xor2_1 _16310_ (.B(net2387),
    .A(net2697),
    .X(_06043_));
 sg13g2_nor3_2 _16311_ (.A(net2439),
    .B(net2657),
    .C(_06043_),
    .Y(_06044_));
 sg13g2_xor2_1 _16312_ (.B(net2302),
    .A(net2357),
    .X(_06046_));
 sg13g2_nor2_2 _16313_ (.A(net2500),
    .B(_06046_),
    .Y(_06047_));
 sg13g2_nor2_1 _16314_ (.A(net2739),
    .B(net2773),
    .Y(_06048_));
 sg13g2_o21ai_1 _16315_ (.B1(_06048_),
    .Y(_06049_),
    .A1(net2483),
    .A2(_05814_));
 sg13g2_xnor2_1 _16316_ (.Y(_06050_),
    .A(_06047_),
    .B(_06049_));
 sg13g2_xnor2_1 _16317_ (.Y(_06051_),
    .A(_06044_),
    .B(_06050_));
 sg13g2_inv_1 _16318_ (.Y(_06052_),
    .A(_06051_));
 sg13g2_nand2b_1 _16319_ (.Y(_06053_),
    .B(_06051_),
    .A_N(_06042_));
 sg13g2_nand2_1 _16320_ (.Y(_06054_),
    .A(_06042_),
    .B(_06052_));
 sg13g2_xor2_1 _16321_ (.B(_06051_),
    .A(_06042_),
    .X(_06055_));
 sg13g2_nand2b_1 _16322_ (.Y(_06057_),
    .B(net2333),
    .A_N(net2480));
 sg13g2_xnor2_1 _16323_ (.Y(_06058_),
    .A(net2346),
    .B(net2650));
 sg13g2_xnor2_1 _16324_ (.Y(_06059_),
    .A(_06057_),
    .B(_06058_));
 sg13g2_nor2_2 _16325_ (.A(net2317),
    .B(net2321),
    .Y(_06060_));
 sg13g2_xor2_1 _16326_ (.B(net2545),
    .A(net2326),
    .X(_06061_));
 sg13g2_xor2_1 _16327_ (.B(_06061_),
    .A(_06060_),
    .X(_06062_));
 sg13g2_xnor2_1 _16328_ (.Y(_06063_),
    .A(_06060_),
    .B(_06061_));
 sg13g2_nand2b_1 _16329_ (.Y(_06064_),
    .B(_06062_),
    .A_N(_06059_));
 sg13g2_xnor2_1 _16330_ (.Y(_06065_),
    .A(_06059_),
    .B(_06062_));
 sg13g2_xor2_1 _16331_ (.B(net2293),
    .A(net2424),
    .X(_06066_));
 sg13g2_xor2_1 _16332_ (.B(_06066_),
    .A(_06065_),
    .X(_06068_));
 sg13g2_xnor2_1 _16333_ (.Y(_06069_),
    .A(_06055_),
    .B(_06068_));
 sg13g2_xor2_1 _16334_ (.B(net2770),
    .A(net2698),
    .X(_06070_));
 sg13g2_nor2_1 _16335_ (.A(net2788),
    .B(net2556),
    .Y(_06071_));
 sg13g2_nor2_1 _16336_ (.A(net2203),
    .B(net2281),
    .Y(_06072_));
 sg13g2_xor2_1 _16337_ (.B(_06072_),
    .A(_06071_),
    .X(_06073_));
 sg13g2_nor2_1 _16338_ (.A(_06070_),
    .B(_06073_),
    .Y(_06074_));
 sg13g2_nand2_1 _16339_ (.Y(_06075_),
    .A(_06070_),
    .B(_06073_));
 sg13g2_nor2b_1 _16340_ (.A(_06074_),
    .B_N(_06075_),
    .Y(_06076_));
 sg13g2_nor2_1 _16341_ (.A(net2537),
    .B(net2601),
    .Y(_06077_));
 sg13g2_xnor2_1 _16342_ (.Y(_06079_),
    .A(_00812_),
    .B(_06077_));
 sg13g2_xor2_1 _16343_ (.B(_06079_),
    .A(_06076_),
    .X(_06080_));
 sg13g2_and2_1 _16344_ (.A(net2758),
    .B(net2318),
    .X(_06081_));
 sg13g2_nor3_1 _16345_ (.A(net2351),
    .B(net2545),
    .C(_06081_),
    .Y(_06082_));
 sg13g2_o21ai_1 _16346_ (.B1(_06082_),
    .Y(_06083_),
    .A1(net2758),
    .A2(net2318));
 sg13g2_o21ai_1 _16347_ (.B1(_00645_),
    .Y(_06084_),
    .A1(net2712),
    .A2(_05880_));
 sg13g2_xnor2_1 _16348_ (.Y(_06085_),
    .A(net2797),
    .B(_06562_));
 sg13g2_nand2b_1 _16349_ (.Y(_06086_),
    .B(_06085_),
    .A_N(_06084_));
 sg13g2_nor2b_1 _16350_ (.A(_06085_),
    .B_N(_06084_),
    .Y(_06087_));
 sg13g2_xnor2_1 _16351_ (.Y(_06088_),
    .A(_06084_),
    .B(_06085_));
 sg13g2_o21ai_1 _16352_ (.B1(_06086_),
    .Y(_06090_),
    .A1(_06083_),
    .A2(_06087_));
 sg13g2_xnor2_1 _16353_ (.Y(_06091_),
    .A(_06083_),
    .B(_06088_));
 sg13g2_xnor2_1 _16354_ (.Y(_06092_),
    .A(net2507),
    .B(net2627));
 sg13g2_nor2_1 _16355_ (.A(net2519),
    .B(net2637),
    .Y(_06093_));
 sg13g2_o21ai_1 _16356_ (.B1(_06093_),
    .Y(_06094_),
    .A1(net2351),
    .A2(_06092_));
 sg13g2_nor3_1 _16357_ (.A(net2351),
    .B(_06092_),
    .C(_06093_),
    .Y(_06095_));
 sg13g2_or3_1 _16358_ (.A(net2350),
    .B(_06092_),
    .C(_06093_),
    .X(_06096_));
 sg13g2_nand2_1 _16359_ (.Y(_06097_),
    .A(_06094_),
    .B(_06096_));
 sg13g2_nor2_1 _16360_ (.A(net2480),
    .B(net2536),
    .Y(_06098_));
 sg13g2_nand2_1 _16361_ (.Y(_06099_),
    .A(net2568),
    .B(_05473_));
 sg13g2_xnor2_1 _16362_ (.Y(_06101_),
    .A(_06098_),
    .B(_06099_));
 sg13g2_xnor2_1 _16363_ (.Y(_06102_),
    .A(_06097_),
    .B(_06101_));
 sg13g2_nand2_1 _16364_ (.Y(_06103_),
    .A(_06091_),
    .B(_06102_));
 sg13g2_nor2_1 _16365_ (.A(_06091_),
    .B(_06102_),
    .Y(_06104_));
 sg13g2_xnor2_1 _16366_ (.Y(_06105_),
    .A(_06091_),
    .B(_06102_));
 sg13g2_xnor2_1 _16367_ (.Y(_06106_),
    .A(_06080_),
    .B(_06105_));
 sg13g2_nor2_1 _16368_ (.A(net2298),
    .B(net2366),
    .Y(_06107_));
 sg13g2_xnor2_1 _16369_ (.Y(_06108_),
    .A(net2383),
    .B(_06107_));
 sg13g2_xor2_1 _16370_ (.B(net2545),
    .A(net2640),
    .X(_06109_));
 sg13g2_xor2_1 _16371_ (.B(net2428),
    .A(net2697),
    .X(_06110_));
 sg13g2_and3_1 _16372_ (.X(_06112_),
    .A(_00895_),
    .B(_06109_),
    .C(_06110_));
 sg13g2_nand3_1 _16373_ (.B(_06109_),
    .C(_06110_),
    .A(_00895_),
    .Y(_06113_));
 sg13g2_a21oi_1 _16374_ (.A1(_06109_),
    .A2(_06110_),
    .Y(_06114_),
    .B1(_00895_));
 sg13g2_nor2_1 _16375_ (.A(_06112_),
    .B(_06114_),
    .Y(_06115_));
 sg13g2_xnor2_1 _16376_ (.Y(_06116_),
    .A(_06108_),
    .B(_06115_));
 sg13g2_and2_1 _16377_ (.A(net2810),
    .B(net2730),
    .X(_06117_));
 sg13g2_nor2_1 _16378_ (.A(net2810),
    .B(net2730),
    .Y(_06118_));
 sg13g2_nor4_2 _16379_ (.A(net2500),
    .B(net2544),
    .C(_06117_),
    .Y(_06119_),
    .D(_06118_));
 sg13g2_nor2b_1 _16380_ (.A(net2649),
    .B_N(net2688),
    .Y(_06120_));
 sg13g2_nor4_2 _16381_ (.A(net2443),
    .B(net2439),
    .C(_05878_),
    .Y(_06121_),
    .D(_06120_));
 sg13g2_nand2_1 _16382_ (.Y(_06123_),
    .A(_06119_),
    .B(_06121_));
 sg13g2_or2_1 _16383_ (.X(_06124_),
    .B(_06121_),
    .A(_06119_));
 sg13g2_xnor2_1 _16384_ (.Y(_06125_),
    .A(_06119_),
    .B(_06121_));
 sg13g2_xnor2_1 _16385_ (.Y(_06126_),
    .A(net2583),
    .B(net2692));
 sg13g2_xnor2_1 _16386_ (.Y(_06127_),
    .A(_06125_),
    .B(_06126_));
 sg13g2_nor2_1 _16387_ (.A(_06116_),
    .B(_06127_),
    .Y(_06128_));
 sg13g2_xnor2_1 _16388_ (.Y(_06129_),
    .A(_06116_),
    .B(_06127_));
 sg13g2_and2_1 _16389_ (.A(net2540),
    .B(net2589),
    .X(_06130_));
 sg13g2_nor3_1 _16390_ (.A(net2808),
    .B(net2797),
    .C(_06130_),
    .Y(_06131_));
 sg13g2_o21ai_1 _16391_ (.B1(_06131_),
    .Y(_06132_),
    .A1(net2540),
    .A2(net2589));
 sg13g2_nand2b_1 _16392_ (.Y(_06134_),
    .B(net2718),
    .A_N(net2708));
 sg13g2_nor2_1 _16393_ (.A(net2445),
    .B(net2777),
    .Y(_06135_));
 sg13g2_xnor2_1 _16394_ (.Y(_06136_),
    .A(_06134_),
    .B(_06135_));
 sg13g2_nor2_1 _16395_ (.A(net2401),
    .B(net2648),
    .Y(_06137_));
 sg13g2_nand2b_1 _16396_ (.Y(_06138_),
    .B(net2527),
    .A_N(net2598));
 sg13g2_xnor2_1 _16397_ (.Y(_06139_),
    .A(_06137_),
    .B(_06138_));
 sg13g2_nor2_1 _16398_ (.A(_06136_),
    .B(_06139_),
    .Y(_06140_));
 sg13g2_and2_1 _16399_ (.A(_06136_),
    .B(_06139_),
    .X(_06141_));
 sg13g2_nor2_1 _16400_ (.A(_06140_),
    .B(_06141_),
    .Y(_06142_));
 sg13g2_xnor2_1 _16401_ (.Y(_06143_),
    .A(_06132_),
    .B(_06142_));
 sg13g2_xnor2_1 _16402_ (.Y(_06145_),
    .A(_06129_),
    .B(_06143_));
 sg13g2_nor2_1 _16403_ (.A(_06106_),
    .B(_06145_),
    .Y(_06146_));
 sg13g2_nand2_1 _16404_ (.Y(_06147_),
    .A(_06106_),
    .B(_06145_));
 sg13g2_xnor2_1 _16405_ (.Y(_06148_),
    .A(_06106_),
    .B(_06145_));
 sg13g2_xnor2_1 _16406_ (.Y(_06149_),
    .A(_06069_),
    .B(_06148_));
 sg13g2_nor2_1 _16407_ (.A(_06035_),
    .B(_06149_),
    .Y(_06150_));
 sg13g2_nand2_1 _16408_ (.Y(_06151_),
    .A(_06035_),
    .B(_06149_));
 sg13g2_xor2_1 _16409_ (.B(_06149_),
    .A(_06035_),
    .X(_06152_));
 sg13g2_xnor2_1 _16410_ (.Y(_06153_),
    .A(net2794),
    .B(net2697));
 sg13g2_nor2_1 _16411_ (.A(net2184),
    .B(net2428),
    .Y(_06154_));
 sg13g2_xnor2_1 _16412_ (.Y(_06156_),
    .A(net2751),
    .B(net2683));
 sg13g2_xnor2_1 _16413_ (.Y(_06157_),
    .A(_06154_),
    .B(_06156_));
 sg13g2_xnor2_1 _16414_ (.Y(_06158_),
    .A(_06153_),
    .B(_06157_));
 sg13g2_nor2_1 _16415_ (.A(net2432),
    .B(net2445),
    .Y(_06159_));
 sg13g2_nor2_1 _16416_ (.A(net2439),
    .B(net2379),
    .Y(_06160_));
 sg13g2_xor2_1 _16417_ (.B(_06160_),
    .A(_06159_),
    .X(_06161_));
 sg13g2_a22oi_1 _16418_ (.Y(_06162_),
    .B1(_05440_),
    .B2(net2560),
    .A2(net2810),
    .A1(net2753));
 sg13g2_o21ai_1 _16419_ (.B1(_06162_),
    .Y(_06163_),
    .A1(net2560),
    .A2(_05440_));
 sg13g2_nand2_1 _16420_ (.Y(_06164_),
    .A(net2339),
    .B(net2636));
 sg13g2_xnor2_1 _16421_ (.Y(_06165_),
    .A(_00910_),
    .B(_06164_));
 sg13g2_nand2_1 _16422_ (.Y(_06167_),
    .A(_06163_),
    .B(_06165_));
 sg13g2_nor2_1 _16423_ (.A(_06163_),
    .B(_06165_),
    .Y(_06168_));
 sg13g2_xnor2_1 _16424_ (.Y(_06169_),
    .A(_06163_),
    .B(_06165_));
 sg13g2_o21ai_1 _16425_ (.B1(_06167_),
    .Y(_06170_),
    .A1(_06161_),
    .A2(_06168_));
 sg13g2_xnor2_1 _16426_ (.Y(_06171_),
    .A(_06161_),
    .B(_06169_));
 sg13g2_nand2_1 _16427_ (.Y(_06172_),
    .A(_06158_),
    .B(_06171_));
 sg13g2_nor2_1 _16428_ (.A(_06158_),
    .B(_06171_),
    .Y(_06173_));
 sg13g2_xor2_1 _16429_ (.B(_06171_),
    .A(_06158_),
    .X(_06174_));
 sg13g2_xor2_1 _16430_ (.B(net2712),
    .A(net2797),
    .X(_06175_));
 sg13g2_nand3_1 _16431_ (.B(_05539_),
    .C(_06175_),
    .A(_05418_),
    .Y(_06176_));
 sg13g2_nor2b_1 _16432_ (.A(net2733),
    .B_N(net2810),
    .Y(_06178_));
 sg13g2_nor3_1 _16433_ (.A(net2770),
    .B(\net.in[192] ),
    .C(_06178_),
    .Y(_06179_));
 sg13g2_nand2_1 _16434_ (.Y(_06180_),
    .A(net2599),
    .B(_06001_));
 sg13g2_xnor2_1 _16435_ (.Y(_06181_),
    .A(_05757_),
    .B(_06180_));
 sg13g2_nor2b_1 _16436_ (.A(_06181_),
    .B_N(_06179_),
    .Y(_06182_));
 sg13g2_nand2b_1 _16437_ (.Y(_06183_),
    .B(_06181_),
    .A_N(_06179_));
 sg13g2_nor2b_1 _16438_ (.A(_06182_),
    .B_N(_06183_),
    .Y(_06184_));
 sg13g2_xnor2_1 _16439_ (.Y(_06185_),
    .A(_06176_),
    .B(_06184_));
 sg13g2_xnor2_1 _16440_ (.Y(_06186_),
    .A(_06174_),
    .B(_06185_));
 sg13g2_xnor2_1 _16441_ (.Y(_06187_),
    .A(net2307),
    .B(net2205));
 sg13g2_nand2_1 _16442_ (.Y(_06189_),
    .A(_00007_),
    .B(_06187_));
 sg13g2_nor4_2 _16443_ (.A(\net.in[35] ),
    .B(net2815),
    .C(net2205),
    .Y(_06190_),
    .D(\net.in[176] ));
 sg13g2_xnor2_1 _16444_ (.Y(_06191_),
    .A(net2251),
    .B(\net.in[209] ));
 sg13g2_xnor2_1 _16445_ (.Y(_06192_),
    .A(net2217),
    .B(_06191_));
 sg13g2_nand2b_1 _16446_ (.Y(_06193_),
    .B(_06190_),
    .A_N(_06192_));
 sg13g2_nor2b_1 _16447_ (.A(_06190_),
    .B_N(_06192_),
    .Y(_06194_));
 sg13g2_xnor2_1 _16448_ (.Y(_06195_),
    .A(_06190_),
    .B(_06192_));
 sg13g2_xnor2_1 _16449_ (.Y(_06196_),
    .A(_06189_),
    .B(_06195_));
 sg13g2_xnor2_1 _16450_ (.Y(_06197_),
    .A(net2316),
    .B(net2314));
 sg13g2_o21ai_1 _16451_ (.B1(_06197_),
    .Y(_06198_),
    .A1(_05132_),
    .A2(net2648));
 sg13g2_inv_1 _16452_ (.Y(_06200_),
    .A(_06198_));
 sg13g2_nor2_1 _16453_ (.A(net2594),
    .B(\net.in[191] ),
    .Y(_06201_));
 sg13g2_xnor2_1 _16454_ (.Y(_06202_),
    .A(net2697),
    .B(net2654));
 sg13g2_a21oi_1 _16455_ (.A1(_00003_),
    .A2(_06201_),
    .Y(_06203_),
    .B1(_06202_));
 sg13g2_nand3_1 _16456_ (.B(_06201_),
    .C(_06202_),
    .A(_00003_),
    .Y(_06204_));
 sg13g2_o21ai_1 _16457_ (.B1(_06204_),
    .Y(_06205_),
    .A1(_06200_),
    .A2(_06203_));
 sg13g2_nand2b_1 _16458_ (.Y(_06206_),
    .B(_06198_),
    .A_N(_06204_));
 sg13g2_a22oi_1 _16459_ (.Y(_06207_),
    .B1(_06205_),
    .B2(_06206_),
    .A2(_06203_),
    .A1(_06200_));
 sg13g2_xor2_1 _16460_ (.B(net2707),
    .A(net2445),
    .X(_06208_));
 sg13g2_a21oi_2 _16461_ (.B1(_06208_),
    .Y(_06209_),
    .A2(net2600),
    .A1(_05187_));
 sg13g2_xnor2_1 _16462_ (.Y(_06211_),
    .A(net2643),
    .B(net2411));
 sg13g2_xnor2_1 _16463_ (.Y(_06212_),
    .A(net2346),
    .B(_06211_));
 sg13g2_nor2_1 _16464_ (.A(net2727),
    .B(net2318),
    .Y(_06213_));
 sg13g2_nor2_1 _16465_ (.A(net2490),
    .B(net2783),
    .Y(_06214_));
 sg13g2_xnor2_1 _16466_ (.Y(_06215_),
    .A(_06213_),
    .B(_06214_));
 sg13g2_nand2_1 _16467_ (.Y(_06216_),
    .A(_06212_),
    .B(_06215_));
 sg13g2_nor2_1 _16468_ (.A(_06212_),
    .B(_06215_),
    .Y(_06217_));
 sg13g2_xnor2_1 _16469_ (.Y(_06218_),
    .A(_06212_),
    .B(_06215_));
 sg13g2_xnor2_1 _16470_ (.Y(_06219_),
    .A(_06209_),
    .B(_06218_));
 sg13g2_nand2_1 _16471_ (.Y(_06220_),
    .A(_06207_),
    .B(_06219_));
 sg13g2_xnor2_1 _16472_ (.Y(_06222_),
    .A(_06207_),
    .B(_06219_));
 sg13g2_nand2_1 _16473_ (.Y(_06223_),
    .A(_06196_),
    .B(_06220_));
 sg13g2_o21ai_1 _16474_ (.B1(_06223_),
    .Y(_06224_),
    .A1(_06207_),
    .A2(_06219_));
 sg13g2_xor2_1 _16475_ (.B(_06222_),
    .A(_06196_),
    .X(_06225_));
 sg13g2_nand2b_1 _16476_ (.Y(_06226_),
    .B(_06225_),
    .A_N(_06186_));
 sg13g2_nand2b_1 _16477_ (.Y(_06227_),
    .B(_06186_),
    .A_N(_06225_));
 sg13g2_nor2_1 _16478_ (.A(net2540),
    .B(_05724_),
    .Y(_06228_));
 sg13g2_a22oi_1 _16479_ (.Y(_06229_),
    .B1(net2374),
    .B2(_05176_),
    .A2(_05187_),
    .A1(net2698));
 sg13g2_o21ai_1 _16480_ (.B1(_06229_),
    .Y(_06230_),
    .A1(_05176_),
    .A2(net2374));
 sg13g2_nand2b_1 _16481_ (.Y(_06231_),
    .B(_06230_),
    .A_N(_06228_));
 sg13g2_nor3_1 _16482_ (.A(net2540),
    .B(_05724_),
    .C(_06230_),
    .Y(_06233_));
 sg13g2_xnor2_1 _16483_ (.Y(_06234_),
    .A(_06228_),
    .B(_06230_));
 sg13g2_nor2_1 _16484_ (.A(net2810),
    .B(net2797),
    .Y(_06235_));
 sg13g2_xnor2_1 _16485_ (.Y(_06236_),
    .A(_06551_),
    .B(_06235_));
 sg13g2_xnor2_1 _16486_ (.Y(_06237_),
    .A(_06234_),
    .B(_06236_));
 sg13g2_or2_1 _16487_ (.X(_06238_),
    .B(net2399),
    .A(net2445));
 sg13g2_nand2_1 _16488_ (.Y(_06239_),
    .A(net2445),
    .B(net2399));
 sg13g2_xnor2_1 _16489_ (.Y(_06240_),
    .A(net2338),
    .B(_00008_));
 sg13g2_xnor2_1 _16490_ (.Y(_06241_),
    .A(net2519),
    .B(_06240_));
 sg13g2_a21oi_1 _16491_ (.A1(_06238_),
    .A2(_06239_),
    .Y(_06242_),
    .B1(_06241_));
 sg13g2_nand3_1 _16492_ (.B(_06239_),
    .C(_06241_),
    .A(_06238_),
    .Y(_06244_));
 sg13g2_nor2b_1 _16493_ (.A(_06242_),
    .B_N(_06244_),
    .Y(_06245_));
 sg13g2_xor2_1 _16494_ (.B(net2627),
    .A(net2465),
    .X(_06246_));
 sg13g2_xnor2_1 _16495_ (.Y(_06247_),
    .A(_06245_),
    .B(_06246_));
 sg13g2_or2_1 _16496_ (.X(_06248_),
    .B(_06247_),
    .A(_06237_));
 sg13g2_nand2_1 _16497_ (.Y(_06249_),
    .A(_06237_),
    .B(_06247_));
 sg13g2_nand2_1 _16498_ (.Y(_06250_),
    .A(_06248_),
    .B(_06249_));
 sg13g2_a21oi_2 _16499_ (.B1(_02427_),
    .Y(_06251_),
    .A2(net2777),
    .A1(_05759_));
 sg13g2_xnor2_1 _16500_ (.Y(_06252_),
    .A(net2390),
    .B(_01113_));
 sg13g2_xnor2_1 _16501_ (.Y(_06253_),
    .A(net2445),
    .B(_06252_));
 sg13g2_nand2b_1 _16502_ (.Y(_06255_),
    .B(_06251_),
    .A_N(_06253_));
 sg13g2_nand2b_1 _16503_ (.Y(_06256_),
    .B(net2266),
    .A_N(net2741));
 sg13g2_nor2_1 _16504_ (.A(_05451_),
    .B(net2293),
    .Y(_06257_));
 sg13g2_xnor2_1 _16505_ (.Y(_06258_),
    .A(_06256_),
    .B(_06257_));
 sg13g2_nor2b_1 _16506_ (.A(_06251_),
    .B_N(_06253_),
    .Y(_06259_));
 sg13g2_a21oi_2 _16507_ (.B1(_06259_),
    .Y(_06260_),
    .A2(_06258_),
    .A1(_06255_));
 sg13g2_xor2_1 _16508_ (.B(_06253_),
    .A(_06251_),
    .X(_06261_));
 sg13g2_xnor2_1 _16509_ (.Y(_06262_),
    .A(_06258_),
    .B(_06261_));
 sg13g2_xnor2_1 _16510_ (.Y(_06263_),
    .A(_06250_),
    .B(_06262_));
 sg13g2_nand2_1 _16511_ (.Y(_06264_),
    .A(_06227_),
    .B(_06263_));
 sg13g2_xnor2_1 _16512_ (.Y(_06266_),
    .A(_06186_),
    .B(_06225_));
 sg13g2_xnor2_1 _16513_ (.Y(_06267_),
    .A(_06263_),
    .B(_06266_));
 sg13g2_xnor2_1 _16514_ (.Y(_06268_),
    .A(_06152_),
    .B(_06267_));
 sg13g2_xnor2_1 _16515_ (.Y(_06269_),
    .A(_05920_),
    .B(_06268_));
 sg13g2_nand2_1 _16516_ (.Y(_06270_),
    .A(net2513),
    .B(_05297_));
 sg13g2_nor2_1 _16517_ (.A(net2539),
    .B(net2602),
    .Y(_06271_));
 sg13g2_xnor2_1 _16518_ (.Y(_06272_),
    .A(_06270_),
    .B(_06271_));
 sg13g2_nand2_1 _16519_ (.Y(_06273_),
    .A(net2566),
    .B(net2702));
 sg13g2_or2_1 _16520_ (.X(_06274_),
    .B(net2702),
    .A(net2566));
 sg13g2_nand2b_1 _16521_ (.Y(_06275_),
    .B(net2381),
    .A_N(net2559));
 sg13g2_nand3_1 _16522_ (.B(_06274_),
    .C(_06275_),
    .A(_06273_),
    .Y(_06277_));
 sg13g2_nor2b_1 _16523_ (.A(net2332),
    .B_N(net2463),
    .Y(_06278_));
 sg13g2_xnor2_1 _16524_ (.Y(_06279_),
    .A(_00005_),
    .B(_06278_));
 sg13g2_nand2b_1 _16525_ (.Y(_06280_),
    .B(_06279_),
    .A_N(_06277_));
 sg13g2_nor2b_1 _16526_ (.A(_06279_),
    .B_N(_06277_),
    .Y(_06281_));
 sg13g2_xnor2_1 _16527_ (.Y(_06282_),
    .A(_06277_),
    .B(_06279_));
 sg13g2_xnor2_1 _16528_ (.Y(_06283_),
    .A(_06272_),
    .B(_06282_));
 sg13g2_xor2_1 _16529_ (.B(net2224),
    .A(net2473),
    .X(_06284_));
 sg13g2_xnor2_1 _16530_ (.Y(_06285_),
    .A(net2368),
    .B(net2329));
 sg13g2_xnor2_1 _16531_ (.Y(_06286_),
    .A(net2453),
    .B(_06285_));
 sg13g2_nor2_1 _16532_ (.A(net2553),
    .B(net2270),
    .Y(_06288_));
 sg13g2_xnor2_1 _16533_ (.Y(_06289_),
    .A(net2354),
    .B(net2255));
 sg13g2_xnor2_1 _16534_ (.Y(_06290_),
    .A(_06288_),
    .B(_06289_));
 sg13g2_nand2_1 _16535_ (.Y(_06291_),
    .A(_06286_),
    .B(_06290_));
 sg13g2_nor2_1 _16536_ (.A(_06286_),
    .B(_06290_),
    .Y(_06292_));
 sg13g2_xor2_1 _16537_ (.B(_06290_),
    .A(_06286_),
    .X(_06293_));
 sg13g2_xnor2_1 _16538_ (.Y(_06294_),
    .A(_06284_),
    .B(_06293_));
 sg13g2_nand2_1 _16539_ (.Y(_06295_),
    .A(_06283_),
    .B(_06294_));
 sg13g2_xor2_1 _16540_ (.B(net2457),
    .A(net2553),
    .X(_06296_));
 sg13g2_nor2_1 _16541_ (.A(net2449),
    .B(net2797),
    .Y(_06297_));
 sg13g2_xnor2_1 _16542_ (.Y(_06299_),
    .A(net2449),
    .B(net2797));
 sg13g2_xnor2_1 _16543_ (.Y(_06300_),
    .A(net2521),
    .B(net2488));
 sg13g2_xnor2_1 _16544_ (.Y(_06301_),
    .A(_06299_),
    .B(_06300_));
 sg13g2_nand2b_1 _16545_ (.Y(_06302_),
    .B(_06301_),
    .A_N(_06296_));
 sg13g2_nor2b_1 _16546_ (.A(_06301_),
    .B_N(_06296_),
    .Y(_06303_));
 sg13g2_xnor2_1 _16547_ (.Y(_06304_),
    .A(_06296_),
    .B(_06301_));
 sg13g2_xor2_1 _16548_ (.B(net2318),
    .A(net2239),
    .X(_06305_));
 sg13g2_xor2_1 _16549_ (.B(net2808),
    .A(net2453),
    .X(_06306_));
 sg13g2_xnor2_1 _16550_ (.Y(_06307_),
    .A(_06305_),
    .B(_06306_));
 sg13g2_xnor2_1 _16551_ (.Y(_06308_),
    .A(_06304_),
    .B(_06307_));
 sg13g2_or2_1 _16552_ (.X(_06310_),
    .B(_06294_),
    .A(_06283_));
 sg13g2_nand2_1 _16553_ (.Y(_06311_),
    .A(_06295_),
    .B(_06308_));
 sg13g2_nor2b_1 _16554_ (.A(net2752),
    .B_N(net2388),
    .Y(_06312_));
 sg13g2_xnor2_1 _16555_ (.Y(_06313_),
    .A(net2571),
    .B(_06312_));
 sg13g2_nor2_1 _16556_ (.A(net2473),
    .B(net2365),
    .Y(_06314_));
 sg13g2_xnor2_1 _16557_ (.Y(_06315_),
    .A(net2316),
    .B(_06314_));
 sg13g2_nand2b_1 _16558_ (.Y(_06316_),
    .B(_06315_),
    .A_N(_06313_));
 sg13g2_xnor2_1 _16559_ (.Y(_06317_),
    .A(net2241),
    .B(net2318));
 sg13g2_a21oi_2 _16560_ (.B1(_06317_),
    .Y(_06318_),
    .A2(net2666),
    .A1(net2200));
 sg13g2_nand2b_1 _16561_ (.Y(_06319_),
    .B(_06313_),
    .A_N(_06315_));
 sg13g2_nand2_1 _16562_ (.Y(_06321_),
    .A(_06316_),
    .B(_06318_));
 sg13g2_nand4_1 _16563_ (.B(_06311_),
    .C(_06319_),
    .A(_06310_),
    .Y(_06322_),
    .D(_06321_));
 sg13g2_inv_1 _16564_ (.Y(_06323_),
    .A(_06322_));
 sg13g2_xor2_1 _16565_ (.B(net2272),
    .A(net2630),
    .X(_06324_));
 sg13g2_a21oi_2 _16566_ (.B1(_06324_),
    .Y(_06325_),
    .A2(_06012_),
    .A1(net2382));
 sg13g2_xor2_1 _16567_ (.B(net2231),
    .A(net2359),
    .X(_06326_));
 sg13g2_and2_1 _16568_ (.A(net2639),
    .B(net2700),
    .X(_06327_));
 sg13g2_nor3_2 _16569_ (.A(_09433_),
    .B(_06326_),
    .C(_06327_),
    .Y(_06328_));
 sg13g2_nand3_1 _16570_ (.B(_06012_),
    .C(_06324_),
    .A(net2381),
    .Y(_06329_));
 sg13g2_o21ai_1 _16571_ (.B1(_06329_),
    .Y(_06330_),
    .A1(_06325_),
    .A2(_06328_));
 sg13g2_a22oi_1 _16572_ (.Y(_06332_),
    .B1(_06319_),
    .B2(_06321_),
    .A2(_06311_),
    .A1(_06310_));
 sg13g2_a21oi_2 _16573_ (.B1(_06332_),
    .Y(_06333_),
    .A2(_06330_),
    .A1(_06322_));
 sg13g2_nand2_1 _16574_ (.Y(_06334_),
    .A(net2195),
    .B(net2328));
 sg13g2_nor2_1 _16575_ (.A(net2195),
    .B(net2328),
    .Y(_06335_));
 sg13g2_o21ai_1 _16576_ (.B1(_06334_),
    .Y(_06336_),
    .A1(net2305),
    .A2(_05550_));
 sg13g2_nor2b_1 _16577_ (.A(net2434),
    .B_N(net2760),
    .Y(_06337_));
 sg13g2_xor2_1 _16578_ (.B(\net.in[191] ),
    .A(net2354),
    .X(_06338_));
 sg13g2_xnor2_1 _16579_ (.Y(_06339_),
    .A(_06337_),
    .B(_06338_));
 sg13g2_o21ai_1 _16580_ (.B1(_06339_),
    .Y(_06340_),
    .A1(_06335_),
    .A2(_06336_));
 sg13g2_xnor2_1 _16581_ (.Y(_06341_),
    .A(net2496),
    .B(_00305_));
 sg13g2_or3_2 _16582_ (.A(_06335_),
    .B(_06336_),
    .C(_06339_),
    .X(_06343_));
 sg13g2_nand2_1 _16583_ (.Y(_06344_),
    .A(_06340_),
    .B(_06341_));
 sg13g2_nand2_2 _16584_ (.Y(_06345_),
    .A(_06343_),
    .B(_06344_));
 sg13g2_nor2_2 _16585_ (.A(net2498),
    .B(net2278),
    .Y(_06346_));
 sg13g2_xnor2_1 _16586_ (.Y(_06347_),
    .A(net2361),
    .B(_06346_));
 sg13g2_a22oi_1 _16587_ (.Y(_06348_),
    .B1(_05858_),
    .B2(_05440_),
    .A2(net2377),
    .A1(_05132_));
 sg13g2_nor2b_1 _16588_ (.A(_06347_),
    .B_N(_06348_),
    .Y(_06349_));
 sg13g2_a21oi_1 _16589_ (.A1(net2326),
    .A2(_05385_),
    .Y(_06350_),
    .B1(_05800_));
 sg13g2_nand2b_1 _16590_ (.Y(_06351_),
    .B(_06347_),
    .A_N(_06348_));
 sg13g2_o21ai_1 _16591_ (.B1(_06351_),
    .Y(_06352_),
    .A1(_06349_),
    .A2(_06350_));
 sg13g2_or2_1 _16592_ (.X(_06354_),
    .B(_06352_),
    .A(_06345_));
 sg13g2_and2_1 _16593_ (.A(_06345_),
    .B(_06352_),
    .X(_06355_));
 sg13g2_xor2_1 _16594_ (.B(net2374),
    .A(net2346),
    .X(_06356_));
 sg13g2_nor2_1 _16595_ (.A(net2191),
    .B(net2203),
    .Y(_06357_));
 sg13g2_xnor2_1 _16596_ (.Y(_06358_),
    .A(net2225),
    .B(net2210));
 sg13g2_xnor2_1 _16597_ (.Y(_06359_),
    .A(_06357_),
    .B(_06358_));
 sg13g2_nor2_1 _16598_ (.A(_06356_),
    .B(_06359_),
    .Y(_06360_));
 sg13g2_xor2_1 _16599_ (.B(net2251),
    .A(net2419),
    .X(_06361_));
 sg13g2_nor2_1 _16600_ (.A(net2817),
    .B(_06361_),
    .Y(_06362_));
 sg13g2_nand2_1 _16601_ (.Y(_06363_),
    .A(_06356_),
    .B(_06359_));
 sg13g2_o21ai_1 _16602_ (.B1(_06363_),
    .Y(_06365_),
    .A1(_06360_),
    .A2(_06362_));
 sg13g2_a21oi_1 _16603_ (.A1(_06354_),
    .A2(_06365_),
    .Y(_06366_),
    .B1(_06355_));
 sg13g2_nand2_1 _16604_ (.Y(_06367_),
    .A(_06333_),
    .B(_06366_));
 sg13g2_nor2_1 _16605_ (.A(_06333_),
    .B(_06366_),
    .Y(_06368_));
 sg13g2_xnor2_1 _16606_ (.Y(_06369_),
    .A(net2643),
    .B(net2600));
 sg13g2_xor2_1 _16607_ (.B(net2238),
    .A(net2593),
    .X(_06370_));
 sg13g2_xnor2_1 _16608_ (.Y(_06371_),
    .A(_06369_),
    .B(_06370_));
 sg13g2_nand2b_1 _16609_ (.Y(_06372_),
    .B(net2554),
    .A_N(net2745));
 sg13g2_xnor2_1 _16610_ (.Y(_06373_),
    .A(net2465),
    .B(net2377));
 sg13g2_xnor2_1 _16611_ (.Y(_06374_),
    .A(_06372_),
    .B(_06373_));
 sg13g2_inv_1 _16612_ (.Y(_06376_),
    .A(_06374_));
 sg13g2_nand2_1 _16613_ (.Y(_06377_),
    .A(_06371_),
    .B(_06376_));
 sg13g2_nor2b_2 _16614_ (.A(\net.in[28] ),
    .B_N(net2512),
    .Y(_06378_));
 sg13g2_nor2_1 _16615_ (.A(net2631),
    .B(net2544),
    .Y(_06379_));
 sg13g2_xnor2_1 _16616_ (.Y(_06380_),
    .A(_06378_),
    .B(_06379_));
 sg13g2_o21ai_1 _16617_ (.B1(_06380_),
    .Y(_06381_),
    .A1(_06371_),
    .A2(_06376_));
 sg13g2_nand2_2 _16618_ (.Y(_06382_),
    .A(_06377_),
    .B(_06381_));
 sg13g2_xor2_1 _16619_ (.B(net2318),
    .A(net2577),
    .X(_06383_));
 sg13g2_nor2_1 _16620_ (.A(net2326),
    .B(net2784),
    .Y(_06384_));
 sg13g2_nand2b_1 _16621_ (.Y(_06385_),
    .B(net2568),
    .A_N(net2426));
 sg13g2_xnor2_1 _16622_ (.Y(_06387_),
    .A(_06384_),
    .B(_06385_));
 sg13g2_nand2_1 _16623_ (.Y(_06388_),
    .A(_06383_),
    .B(_06387_));
 sg13g2_a22oi_1 _16624_ (.Y(_06389_),
    .B1(net2227),
    .B2(_05561_),
    .A2(_05319_),
    .A1(net2523));
 sg13g2_o21ai_1 _16625_ (.B1(_06389_),
    .Y(_06390_),
    .A1(net2523),
    .A2(_05319_));
 sg13g2_nor2_1 _16626_ (.A(_06383_),
    .B(_06387_),
    .Y(_06391_));
 sg13g2_a21oi_2 _16627_ (.B1(_06391_),
    .Y(_06392_),
    .A2(_06390_),
    .A1(_06388_));
 sg13g2_nor2_1 _16628_ (.A(_06382_),
    .B(_06392_),
    .Y(_06393_));
 sg13g2_nor2_1 _16629_ (.A(net2349),
    .B(net2310),
    .Y(_06394_));
 sg13g2_xnor2_1 _16630_ (.Y(_06395_),
    .A(_00002_),
    .B(_06394_));
 sg13g2_nor2b_1 _16631_ (.A(net2640),
    .B_N(net2261),
    .Y(_06396_));
 sg13g2_xnor2_1 _16632_ (.Y(_06398_),
    .A(net2313),
    .B(\net.in[175] ));
 sg13g2_xnor2_1 _16633_ (.Y(_06399_),
    .A(_06396_),
    .B(_06398_));
 sg13g2_nor2_1 _16634_ (.A(_06395_),
    .B(_06399_),
    .Y(_06400_));
 sg13g2_xor2_1 _16635_ (.B(net2583),
    .A(net2541),
    .X(_06401_));
 sg13g2_xnor2_1 _16636_ (.Y(_06402_),
    .A(net2203),
    .B(\net.in[129] ));
 sg13g2_xnor2_1 _16637_ (.Y(_06403_),
    .A(_06401_),
    .B(_06402_));
 sg13g2_nand2_1 _16638_ (.Y(_06404_),
    .A(_06395_),
    .B(_06399_));
 sg13g2_o21ai_1 _16639_ (.B1(_06404_),
    .Y(_06405_),
    .A1(_06400_),
    .A2(_06403_));
 sg13g2_nor2_1 _16640_ (.A(_06393_),
    .B(_06405_),
    .Y(_06406_));
 sg13g2_a21oi_2 _16641_ (.B1(_06406_),
    .Y(_06407_),
    .A2(_06392_),
    .A1(_06382_));
 sg13g2_a21o_1 _16642_ (.A2(_06407_),
    .A1(_06367_),
    .B1(_06368_),
    .X(_06409_));
 sg13g2_xnor2_1 _16643_ (.Y(_06410_),
    .A(net2470),
    .B(net2563));
 sg13g2_xnor2_1 _16644_ (.Y(_06411_),
    .A(net2531),
    .B(net2495));
 sg13g2_nor2_1 _16645_ (.A(_06410_),
    .B(_06411_),
    .Y(_06412_));
 sg13g2_nor2_1 _16646_ (.A(net2198),
    .B(net2210),
    .Y(_06413_));
 sg13g2_xor2_1 _16647_ (.B(net2188),
    .A(net2663),
    .X(_06414_));
 sg13g2_xnor2_1 _16648_ (.Y(_06415_),
    .A(_06413_),
    .B(_06414_));
 sg13g2_nand2_1 _16649_ (.Y(_06416_),
    .A(_06410_),
    .B(_06411_));
 sg13g2_a21o_1 _16650_ (.A2(_06416_),
    .A1(_06415_),
    .B1(_06412_),
    .X(_06417_));
 sg13g2_xnor2_1 _16651_ (.Y(_06418_),
    .A(net2733),
    .B(net2812));
 sg13g2_xnor2_1 _16652_ (.Y(_06420_),
    .A(net2495),
    .B(_06418_));
 sg13g2_xor2_1 _16653_ (.B(net2369),
    .A(net2758),
    .X(_06421_));
 sg13g2_xor2_1 _16654_ (.B(net2706),
    .A(net2544),
    .X(_06422_));
 sg13g2_xor2_1 _16655_ (.B(net2536),
    .A(net2527),
    .X(_06423_));
 sg13g2_nor2_2 _16656_ (.A(_06422_),
    .B(_06423_),
    .Y(_06424_));
 sg13g2_nand2_1 _16657_ (.Y(_06425_),
    .A(_06420_),
    .B(_06421_));
 sg13g2_o21ai_1 _16658_ (.B1(_06424_),
    .Y(_06426_),
    .A1(_06420_),
    .A2(_06421_));
 sg13g2_nand3_1 _16659_ (.B(_06425_),
    .C(_06426_),
    .A(_06417_),
    .Y(_06427_));
 sg13g2_inv_1 _16660_ (.Y(_06428_),
    .A(_06427_));
 sg13g2_a21oi_1 _16661_ (.A1(_06425_),
    .A2(_06426_),
    .Y(_06429_),
    .B1(_06417_));
 sg13g2_nor2b_1 _16662_ (.A(net2261),
    .B_N(net2360),
    .Y(_06431_));
 sg13g2_nor2b_1 _16663_ (.A(net2360),
    .B_N(net2261),
    .Y(_06432_));
 sg13g2_nor2b_1 _16664_ (.A(net2544),
    .B_N(\net.in[143] ),
    .Y(_06433_));
 sg13g2_nor3_2 _16665_ (.A(_06431_),
    .B(_06432_),
    .C(_06433_),
    .Y(_06434_));
 sg13g2_xor2_1 _16666_ (.B(net2227),
    .A(net2476),
    .X(_06435_));
 sg13g2_nand2b_1 _16667_ (.Y(_06436_),
    .B(_06435_),
    .A_N(_06434_));
 sg13g2_xnor2_1 _16668_ (.Y(_06437_),
    .A(net2575),
    .B(net2549));
 sg13g2_xor2_1 _16669_ (.B(net2206),
    .A(net2646),
    .X(_06438_));
 sg13g2_xnor2_1 _16670_ (.Y(_06439_),
    .A(_06437_),
    .B(_06438_));
 sg13g2_nor2b_1 _16671_ (.A(_06435_),
    .B_N(_06434_),
    .Y(_06440_));
 sg13g2_o21ai_1 _16672_ (.B1(_06436_),
    .Y(_06442_),
    .A1(_06439_),
    .A2(_06440_));
 sg13g2_a21oi_1 _16673_ (.A1(_06427_),
    .A2(_06442_),
    .Y(_06443_),
    .B1(_06429_));
 sg13g2_nor2_1 _16674_ (.A(_05297_),
    .B(net2230),
    .Y(_06444_));
 sg13g2_xnor2_1 _16675_ (.Y(_06445_),
    .A(net2527),
    .B(_06444_));
 sg13g2_nor2_1 _16676_ (.A(net2452),
    .B(net2241),
    .Y(_06446_));
 sg13g2_xnor2_1 _16677_ (.Y(_06447_),
    .A(_00001_),
    .B(_06446_));
 sg13g2_xnor2_1 _16678_ (.Y(_06448_),
    .A(net2536),
    .B(net2544));
 sg13g2_nand2_1 _16679_ (.Y(_06449_),
    .A(_06445_),
    .B(_06447_));
 sg13g2_o21ai_1 _16680_ (.B1(_06448_),
    .Y(_06450_),
    .A1(_06445_),
    .A2(_06447_));
 sg13g2_nand2_1 _16681_ (.Y(_06451_),
    .A(net2350),
    .B(net2283));
 sg13g2_or2_1 _16682_ (.X(_06453_),
    .B(net2283),
    .A(net2350));
 sg13g2_nand2b_1 _16683_ (.Y(_06454_),
    .B(net2593),
    .A_N(net2432));
 sg13g2_nand3_1 _16684_ (.B(_06453_),
    .C(_06454_),
    .A(_06451_),
    .Y(_06455_));
 sg13g2_nor2_1 _16685_ (.A(net2361),
    .B(net2545),
    .Y(_06456_));
 sg13g2_xor2_1 _16686_ (.B(net2515),
    .A(net2531),
    .X(_06457_));
 sg13g2_xnor2_1 _16687_ (.Y(_06458_),
    .A(_06456_),
    .B(_06457_));
 sg13g2_nand2_1 _16688_ (.Y(_06459_),
    .A(_06455_),
    .B(_06458_));
 sg13g2_nand2b_1 _16689_ (.Y(_06460_),
    .B(net2432),
    .A_N(net2663));
 sg13g2_nor2_1 _16690_ (.A(net2307),
    .B(net2400),
    .Y(_06461_));
 sg13g2_xnor2_1 _16691_ (.Y(_06462_),
    .A(_06460_),
    .B(_06461_));
 sg13g2_or2_1 _16692_ (.X(_06464_),
    .B(_06458_),
    .A(_06455_));
 sg13g2_nand2_1 _16693_ (.Y(_06465_),
    .A(_06459_),
    .B(_06462_));
 sg13g2_nand4_1 _16694_ (.B(_06450_),
    .C(_06464_),
    .A(_06449_),
    .Y(_06466_),
    .D(_06465_));
 sg13g2_inv_1 _16695_ (.Y(_06467_),
    .A(_06466_));
 sg13g2_a22oi_1 _16696_ (.Y(_06468_),
    .B1(_06464_),
    .B2(_06465_),
    .A2(_06450_),
    .A1(_06449_));
 sg13g2_nand2b_1 _16697_ (.Y(_06469_),
    .B(net2326),
    .A_N(net2470));
 sg13g2_nand2b_1 _16698_ (.Y(_06470_),
    .B(net2342),
    .A_N(net2203));
 sg13g2_xnor2_1 _16699_ (.Y(_06471_),
    .A(net2323),
    .B(\net.in[218] ));
 sg13g2_and3_1 _16700_ (.X(_06472_),
    .A(_06469_),
    .B(_06470_),
    .C(_06471_));
 sg13g2_nor2b_1 _16701_ (.A(net2532),
    .B_N(net2542),
    .Y(_06473_));
 sg13g2_xor2_1 _16702_ (.B(net2541),
    .A(net2531),
    .X(_06475_));
 sg13g2_xor2_1 _16703_ (.B(net2210),
    .A(net2577),
    .X(_06476_));
 sg13g2_xnor2_1 _16704_ (.Y(_06477_),
    .A(_06475_),
    .B(_06476_));
 sg13g2_a21oi_1 _16705_ (.A1(_06469_),
    .A2(_06470_),
    .Y(_06478_),
    .B1(_06471_));
 sg13g2_nor2_1 _16706_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sg13g2_nor2_1 _16707_ (.A(_06472_),
    .B(_06479_),
    .Y(_06480_));
 sg13g2_a21oi_1 _16708_ (.A1(_06466_),
    .A2(_06480_),
    .Y(_06481_),
    .B1(_06468_));
 sg13g2_nand2_1 _16709_ (.Y(_06482_),
    .A(_06443_),
    .B(_06481_));
 sg13g2_inv_1 _16710_ (.Y(_06483_),
    .A(_06482_));
 sg13g2_nor2_1 _16711_ (.A(_06443_),
    .B(_06481_),
    .Y(_06484_));
 sg13g2_nand2_1 _16712_ (.Y(_06486_),
    .A(net2472),
    .B(net2293));
 sg13g2_a22oi_1 _16713_ (.Y(_06487_),
    .B1(_05484_),
    .B2(_05044_),
    .A2(_05363_),
    .A1(net2515));
 sg13g2_xnor2_1 _16714_ (.Y(_06488_),
    .A(net2698),
    .B(net2657));
 sg13g2_a21oi_1 _16715_ (.A1(_06486_),
    .A2(_06487_),
    .Y(_06489_),
    .B1(_06488_));
 sg13g2_xnor2_1 _16716_ (.Y(_06490_),
    .A(net2333),
    .B(net2227));
 sg13g2_nand3_1 _16717_ (.B(_06487_),
    .C(_06488_),
    .A(_06486_),
    .Y(_06491_));
 sg13g2_o21ai_1 _16718_ (.B1(_06491_),
    .Y(_06492_),
    .A1(_06489_),
    .A2(_06490_));
 sg13g2_xor2_1 _16719_ (.B(\net.in[208] ),
    .A(net2802),
    .X(_06493_));
 sg13g2_xor2_1 _16720_ (.B(net2760),
    .A(net2807),
    .X(_06494_));
 sg13g2_nor2_2 _16721_ (.A(_06493_),
    .B(_06494_),
    .Y(_06495_));
 sg13g2_nor2b_1 _16722_ (.A(net2430),
    .B_N(net2791),
    .Y(_06497_));
 sg13g2_xnor2_1 _16723_ (.Y(_06498_),
    .A(_00625_),
    .B(_06497_));
 sg13g2_nor2b_1 _16724_ (.A(_06498_),
    .B_N(_06495_),
    .Y(_06499_));
 sg13g2_xnor2_1 _16725_ (.Y(_06500_),
    .A(net2357),
    .B(\net.in[175] ));
 sg13g2_xnor2_1 _16726_ (.Y(_06501_),
    .A(_05088_),
    .B(_06500_));
 sg13g2_nand2b_1 _16727_ (.Y(_06502_),
    .B(_06498_),
    .A_N(_06495_));
 sg13g2_o21ai_1 _16728_ (.B1(_06502_),
    .Y(_06503_),
    .A1(_06499_),
    .A2(_06501_));
 sg13g2_nand2_1 _16729_ (.Y(_06504_),
    .A(_06492_),
    .B(_06503_));
 sg13g2_a22oi_1 _16730_ (.Y(_06505_),
    .B1(_05957_),
    .B2(net2376),
    .A2(net2784),
    .A1(_05792_));
 sg13g2_xor2_1 _16731_ (.B(net2293),
    .A(net2403),
    .X(_06506_));
 sg13g2_xnor2_1 _16732_ (.Y(_06508_),
    .A(net2598),
    .B(net2600));
 sg13g2_nand2_1 _16733_ (.Y(_06509_),
    .A(_06506_),
    .B(_06508_));
 sg13g2_o21ai_1 _16734_ (.B1(_00766_),
    .Y(_06510_),
    .A1(_05484_),
    .A2(net2200));
 sg13g2_nor2_1 _16735_ (.A(_06505_),
    .B(_06509_),
    .Y(_06511_));
 sg13g2_nor2_1 _16736_ (.A(_06510_),
    .B(_06511_),
    .Y(_06512_));
 sg13g2_a21oi_1 _16737_ (.A1(_06505_),
    .A2(_06509_),
    .Y(_06513_),
    .B1(_06512_));
 sg13g2_o21ai_1 _16738_ (.B1(_06513_),
    .Y(_06514_),
    .A1(_06492_),
    .A2(_06503_));
 sg13g2_nand2_2 _16739_ (.Y(_06515_),
    .A(_06504_),
    .B(_06514_));
 sg13g2_and2_1 _16740_ (.A(_06482_),
    .B(_06515_),
    .X(_06516_));
 sg13g2_or3_1 _16741_ (.A(_06409_),
    .B(_06484_),
    .C(_06516_),
    .X(_06517_));
 sg13g2_o21ai_1 _16742_ (.B1(_06409_),
    .Y(_06519_),
    .A1(_06484_),
    .A2(_06516_));
 sg13g2_inv_1 _16743_ (.Y(_06520_),
    .A(_06519_));
 sg13g2_xor2_1 _16744_ (.B(net2383),
    .A(net2290),
    .X(_06521_));
 sg13g2_nor2_1 _16745_ (.A(net2583),
    .B(net2706),
    .Y(_06522_));
 sg13g2_nor2b_1 _16746_ (.A(net2326),
    .B_N(net2366),
    .Y(_06523_));
 sg13g2_xnor2_1 _16747_ (.Y(_06524_),
    .A(_06522_),
    .B(_06523_));
 sg13g2_nand2b_1 _16748_ (.Y(_06525_),
    .B(_06524_),
    .A_N(_06521_));
 sg13g2_nand2_1 _16749_ (.Y(_06526_),
    .A(net2789),
    .B(_05726_));
 sg13g2_xnor2_1 _16750_ (.Y(_06527_),
    .A(\net.in[127] ),
    .B(\net.in[175] ));
 sg13g2_xnor2_1 _16751_ (.Y(_06528_),
    .A(_06526_),
    .B(_06527_));
 sg13g2_nand2b_1 _16752_ (.Y(_06530_),
    .B(_06521_),
    .A_N(_06524_));
 sg13g2_nand2_1 _16753_ (.Y(_06531_),
    .A(_06528_),
    .B(_06530_));
 sg13g2_xor2_1 _16754_ (.B(net2643),
    .A(net2598),
    .X(_06532_));
 sg13g2_nor2_1 _16755_ (.A(net2302),
    .B(net2589),
    .Y(_06533_));
 sg13g2_xor2_1 _16756_ (.B(net2206),
    .A(net2387),
    .X(_06534_));
 sg13g2_xnor2_1 _16757_ (.Y(_06535_),
    .A(_06533_),
    .B(_06534_));
 sg13g2_nand2_1 _16758_ (.Y(_06536_),
    .A(_06532_),
    .B(_06535_));
 sg13g2_xor2_1 _16759_ (.B(\net.in[175] ),
    .A(net2278),
    .X(_06537_));
 sg13g2_nand2_2 _16760_ (.Y(_06538_),
    .A(\net.in[237] ),
    .B(_06056_));
 sg13g2_xnor2_1 _16761_ (.Y(_06539_),
    .A(_06537_),
    .B(_06538_));
 sg13g2_or2_1 _16762_ (.X(_06541_),
    .B(_06535_),
    .A(_06532_));
 sg13g2_nand2b_1 _16763_ (.Y(_06542_),
    .B(_06541_),
    .A_N(_06539_));
 sg13g2_a22oi_1 _16764_ (.Y(_06543_),
    .B1(_06536_),
    .B2(_06542_),
    .A2(_06531_),
    .A1(_06525_));
 sg13g2_nand4_1 _16765_ (.B(_06531_),
    .C(_06536_),
    .A(_06525_),
    .Y(_06544_),
    .D(_06542_));
 sg13g2_xor2_1 _16766_ (.B(net2419),
    .A(net2508),
    .X(_06545_));
 sg13g2_nor2_1 _16767_ (.A(net2283),
    .B(net2321),
    .Y(_06546_));
 sg13g2_xnor2_1 _16768_ (.Y(_06547_),
    .A(net2219),
    .B(net2408));
 sg13g2_xnor2_1 _16769_ (.Y(_06548_),
    .A(_06546_),
    .B(_06547_));
 sg13g2_nor2_1 _16770_ (.A(_06545_),
    .B(_06548_),
    .Y(_06549_));
 sg13g2_nor2_1 _16771_ (.A(net2495),
    .B(net2208),
    .Y(_06550_));
 sg13g2_xnor2_1 _16772_ (.Y(_06552_),
    .A(_06166_),
    .B(_06550_));
 sg13g2_nand2_1 _16773_ (.Y(_06553_),
    .A(_06545_),
    .B(_06548_));
 sg13g2_o21ai_1 _16774_ (.B1(_06553_),
    .Y(_06554_),
    .A1(_06549_),
    .A2(_06552_));
 sg13g2_o21ai_1 _16775_ (.B1(_06544_),
    .Y(_06555_),
    .A1(_06543_),
    .A2(_06554_));
 sg13g2_xnor2_1 _16776_ (.Y(_06556_),
    .A(net2208),
    .B(_06401_));
 sg13g2_nor2_1 _16777_ (.A(net2317),
    .B(_02183_),
    .Y(_06557_));
 sg13g2_nor2b_1 _16778_ (.A(net2242),
    .B_N(net2316),
    .Y(_06558_));
 sg13g2_o21ai_1 _16779_ (.B1(_06556_),
    .Y(_06559_),
    .A1(_06557_),
    .A2(_06558_));
 sg13g2_xor2_1 _16780_ (.B(net2363),
    .A(\net.in[129] ),
    .X(_06560_));
 sg13g2_xor2_1 _16781_ (.B(net2247),
    .A(net2188),
    .X(_06561_));
 sg13g2_xnor2_1 _16782_ (.Y(_06563_),
    .A(_06560_),
    .B(_06561_));
 sg13g2_or3_1 _16783_ (.A(_06556_),
    .B(_06557_),
    .C(_06558_),
    .X(_06564_));
 sg13g2_nand2_1 _16784_ (.Y(_06565_),
    .A(_06559_),
    .B(_06563_));
 sg13g2_xor2_1 _16785_ (.B(net2203),
    .A(net2428),
    .X(_06566_));
 sg13g2_xnor2_1 _16786_ (.Y(_06567_),
    .A(net2470),
    .B(net2490));
 sg13g2_nor3_1 _16787_ (.A(net2527),
    .B(_06566_),
    .C(_06567_),
    .Y(_06568_));
 sg13g2_xnor2_1 _16788_ (.Y(_06569_),
    .A(net2601),
    .B(net2650));
 sg13g2_nand3b_1 _16789_ (.B(_06569_),
    .C(net2302),
    .Y(_06570_),
    .A_N(\net.in[110] ));
 sg13g2_o21ai_1 _16790_ (.B1(_06567_),
    .Y(_06571_),
    .A1(net2527),
    .A2(_06566_));
 sg13g2_o21ai_1 _16791_ (.B1(_06571_),
    .Y(_06572_),
    .A1(_06568_),
    .A2(_06570_));
 sg13g2_a21oi_1 _16792_ (.A1(_06564_),
    .A2(_06565_),
    .Y(_06574_),
    .B1(_06572_));
 sg13g2_nand3_1 _16793_ (.B(_06565_),
    .C(_06572_),
    .A(_06564_),
    .Y(_06575_));
 sg13g2_nor2b_1 _16794_ (.A(net2598),
    .B_N(net2795),
    .Y(_06576_));
 sg13g2_xnor2_1 _16795_ (.Y(_06577_),
    .A(_00003_),
    .B(_06576_));
 sg13g2_xnor2_1 _16796_ (.Y(_06578_),
    .A(net2628),
    .B(net2563));
 sg13g2_nor2_1 _16797_ (.A(_06577_),
    .B(_06578_),
    .Y(_06579_));
 sg13g2_xor2_1 _16798_ (.B(net2286),
    .A(net2417),
    .X(_06580_));
 sg13g2_xor2_1 _16799_ (.B(net2815),
    .A(net2233),
    .X(_06581_));
 sg13g2_nor2_2 _16800_ (.A(_06580_),
    .B(_06581_),
    .Y(_06582_));
 sg13g2_nor2_1 _16801_ (.A(_06579_),
    .B(_06582_),
    .Y(_06583_));
 sg13g2_a21oi_2 _16802_ (.B1(_06583_),
    .Y(_06585_),
    .A2(_06578_),
    .A1(_06577_));
 sg13g2_o21ai_1 _16803_ (.B1(_06575_),
    .Y(_06586_),
    .A1(_06574_),
    .A2(_06585_));
 sg13g2_nor2_1 _16804_ (.A(_06555_),
    .B(_06586_),
    .Y(_06587_));
 sg13g2_nand2_1 _16805_ (.Y(_06588_),
    .A(_06555_),
    .B(_06586_));
 sg13g2_xnor2_1 _16806_ (.Y(_06589_),
    .A(net2451),
    .B(net2288));
 sg13g2_xnor2_1 _16807_ (.Y(_06590_),
    .A(\net.in[145] ),
    .B(net2305));
 sg13g2_nand2_2 _16808_ (.Y(_06591_),
    .A(_06589_),
    .B(_06590_));
 sg13g2_a22oi_1 _16809_ (.Y(_06592_),
    .B1(_05704_),
    .B2(net2419),
    .A2(_05352_),
    .A1(_05099_));
 sg13g2_o21ai_1 _16810_ (.B1(_06592_),
    .Y(_06593_),
    .A1(_05099_),
    .A2(_05352_));
 sg13g2_or2_1 _16811_ (.X(_06594_),
    .B(_06593_),
    .A(_06591_));
 sg13g2_nor3_2 _16812_ (.A(net2593),
    .B(net2210),
    .C(_08410_),
    .Y(_06596_));
 sg13g2_and2_1 _16813_ (.A(_06591_),
    .B(_06593_),
    .X(_06597_));
 sg13g2_a21oi_2 _16814_ (.B1(_06597_),
    .Y(_06598_),
    .A2(_06596_),
    .A1(_06594_));
 sg13g2_nor2b_1 _16815_ (.A(net2636),
    .B_N(net2272),
    .Y(_06599_));
 sg13g2_nor3_1 _16816_ (.A(\net.in[4] ),
    .B(net2314),
    .C(_06599_),
    .Y(_06600_));
 sg13g2_nor2_2 _16817_ (.A(net2589),
    .B(net2593),
    .Y(_06601_));
 sg13g2_nor2_1 _16818_ (.A(net2486),
    .B(net2767),
    .Y(_06602_));
 sg13g2_xor2_1 _16819_ (.B(_06602_),
    .A(_06601_),
    .X(_06603_));
 sg13g2_or4_1 _16820_ (.A(\net.in[4] ),
    .B(net2314),
    .C(_06599_),
    .D(_06603_),
    .X(_06604_));
 sg13g2_a22oi_1 _16821_ (.Y(_06605_),
    .B1(_05979_),
    .B2(net2794),
    .A2(_05902_),
    .A1(\net.in[159] ));
 sg13g2_o21ai_1 _16822_ (.B1(_06605_),
    .Y(_06607_),
    .A1(net2404),
    .A2(_05902_));
 sg13g2_nor2b_1 _16823_ (.A(_06600_),
    .B_N(_06603_),
    .Y(_06608_));
 sg13g2_a21oi_2 _16824_ (.B1(_06608_),
    .Y(_06609_),
    .A2(_06607_),
    .A1(_06604_));
 sg13g2_nand2_1 _16825_ (.Y(_06610_),
    .A(_06598_),
    .B(_06609_));
 sg13g2_or2_1 _16826_ (.X(_06611_),
    .B(net2803),
    .A(net2593));
 sg13g2_a22oi_1 _16827_ (.Y(_06612_),
    .B1(net2593),
    .B2(net2803),
    .A2(net2462),
    .A1(net2419));
 sg13g2_xor2_1 _16828_ (.B(net2536),
    .A(net2617),
    .X(_06613_));
 sg13g2_xnor2_1 _16829_ (.Y(_06614_),
    .A(net2233),
    .B(net2379));
 sg13g2_nand4_1 _16830_ (.B(_06612_),
    .C(_06613_),
    .A(_06611_),
    .Y(_06615_),
    .D(_06614_));
 sg13g2_inv_1 _16831_ (.Y(_06616_),
    .A(_06615_));
 sg13g2_nor2_1 _16832_ (.A(net2242),
    .B(net2490),
    .Y(_06618_));
 sg13g2_xnor2_1 _16833_ (.Y(_06619_),
    .A(net2651),
    .B(_06618_));
 sg13g2_a22oi_1 _16834_ (.Y(_06620_),
    .B1(_06613_),
    .B2(_06614_),
    .A2(_06612_),
    .A1(_06611_));
 sg13g2_a21oi_2 _16835_ (.B1(_06620_),
    .Y(_06621_),
    .A2(_06619_),
    .A1(_06615_));
 sg13g2_o21ai_1 _16836_ (.B1(_06621_),
    .Y(_06622_),
    .A1(_06598_),
    .A2(_06609_));
 sg13g2_nand2_1 _16837_ (.Y(_06623_),
    .A(_06610_),
    .B(_06622_));
 sg13g2_o21ai_1 _16838_ (.B1(_06588_),
    .Y(_06624_),
    .A1(_06587_),
    .A2(_06623_));
 sg13g2_a21oi_2 _16839_ (.B1(_06520_),
    .Y(_06625_),
    .A2(_06624_),
    .A1(_06517_));
 sg13g2_inv_1 _16840_ (.Y(_06626_),
    .A(_06625_));
 sg13g2_xnor2_1 _16841_ (.Y(_06627_),
    .A(_06347_),
    .B(_06348_));
 sg13g2_xnor2_1 _16842_ (.Y(_06629_),
    .A(_06350_),
    .B(_06627_));
 sg13g2_xnor2_1 _16843_ (.Y(_06630_),
    .A(_06356_),
    .B(_06359_));
 sg13g2_xnor2_1 _16844_ (.Y(_06631_),
    .A(_06362_),
    .B(_06630_));
 sg13g2_nand2b_1 _16845_ (.Y(_06632_),
    .B(_06629_),
    .A_N(_06631_));
 sg13g2_nand2b_1 _16846_ (.Y(_06633_),
    .B(_06631_),
    .A_N(_06629_));
 sg13g2_xnor2_1 _16847_ (.Y(_06634_),
    .A(_06629_),
    .B(_06631_));
 sg13g2_xnor2_1 _16848_ (.Y(_06635_),
    .A(_06383_),
    .B(_06387_));
 sg13g2_xnor2_1 _16849_ (.Y(_06636_),
    .A(_06390_),
    .B(_06635_));
 sg13g2_xnor2_1 _16850_ (.Y(_06637_),
    .A(_06634_),
    .B(_06636_));
 sg13g2_xor2_1 _16851_ (.B(_06315_),
    .A(_06313_),
    .X(_06638_));
 sg13g2_xnor2_1 _16852_ (.Y(_06640_),
    .A(_06318_),
    .B(_06638_));
 sg13g2_or2_1 _16853_ (.X(_06641_),
    .B(_06329_),
    .A(_06328_));
 sg13g2_a22oi_1 _16854_ (.Y(_06642_),
    .B1(_06330_),
    .B2(_06641_),
    .A2(_06328_),
    .A1(_06325_));
 sg13g2_nor2_1 _16855_ (.A(_06640_),
    .B(_06642_),
    .Y(_06643_));
 sg13g2_nand2_1 _16856_ (.Y(_06644_),
    .A(_06640_),
    .B(_06642_));
 sg13g2_xor2_1 _16857_ (.B(_06642_),
    .A(_06640_),
    .X(_06645_));
 sg13g2_nand2_1 _16858_ (.Y(_06646_),
    .A(_06340_),
    .B(_06343_));
 sg13g2_xor2_1 _16859_ (.B(_06646_),
    .A(_06341_),
    .X(_06647_));
 sg13g2_xnor2_1 _16860_ (.Y(_06648_),
    .A(_06645_),
    .B(_06647_));
 sg13g2_inv_1 _16861_ (.Y(_06649_),
    .A(_06648_));
 sg13g2_nand2_1 _16862_ (.Y(_06651_),
    .A(_06637_),
    .B(_06649_));
 sg13g2_xnor2_1 _16863_ (.Y(_06652_),
    .A(_06445_),
    .B(_06447_));
 sg13g2_xnor2_1 _16864_ (.Y(_06653_),
    .A(_06448_),
    .B(_06652_));
 sg13g2_xor2_1 _16865_ (.B(_06374_),
    .A(_06371_),
    .X(_06654_));
 sg13g2_xnor2_1 _16866_ (.Y(_06655_),
    .A(_06380_),
    .B(_06654_));
 sg13g2_xnor2_1 _16867_ (.Y(_06656_),
    .A(_06395_),
    .B(_06399_));
 sg13g2_xnor2_1 _16868_ (.Y(_06657_),
    .A(_06403_),
    .B(_06656_));
 sg13g2_nor2_1 _16869_ (.A(_06655_),
    .B(_06657_),
    .Y(_06658_));
 sg13g2_and2_1 _16870_ (.A(_06655_),
    .B(_06657_),
    .X(_06659_));
 sg13g2_inv_1 _16871_ (.Y(_06660_),
    .A(_06659_));
 sg13g2_nor2_1 _16872_ (.A(_06658_),
    .B(_06659_),
    .Y(_06662_));
 sg13g2_a21oi_1 _16873_ (.A1(_06653_),
    .A2(_06660_),
    .Y(_06663_),
    .B1(_06658_));
 sg13g2_xnor2_1 _16874_ (.Y(_06664_),
    .A(_06653_),
    .B(_06662_));
 sg13g2_o21ai_1 _16875_ (.B1(_06664_),
    .Y(_06665_),
    .A1(_06637_),
    .A2(_06649_));
 sg13g2_xnor2_1 _16876_ (.Y(_06666_),
    .A(_06420_),
    .B(_06421_));
 sg13g2_xnor2_1 _16877_ (.Y(_06667_),
    .A(_06424_),
    .B(_06666_));
 sg13g2_xnor2_1 _16878_ (.Y(_06668_),
    .A(_06434_),
    .B(_06435_));
 sg13g2_xnor2_1 _16879_ (.Y(_06669_),
    .A(_06439_),
    .B(_06668_));
 sg13g2_or2_1 _16880_ (.X(_06670_),
    .B(_06669_),
    .A(_06667_));
 sg13g2_xor2_1 _16881_ (.B(_06669_),
    .A(_06667_),
    .X(_06671_));
 sg13g2_nand2b_1 _16882_ (.Y(_06673_),
    .B(_06491_),
    .A_N(_06489_));
 sg13g2_xor2_1 _16883_ (.B(_06673_),
    .A(_06490_),
    .X(_06674_));
 sg13g2_xnor2_1 _16884_ (.Y(_06675_),
    .A(_06671_),
    .B(_06674_));
 sg13g2_nand2_1 _16885_ (.Y(_06676_),
    .A(_06412_),
    .B(_06415_));
 sg13g2_nor2_1 _16886_ (.A(_06415_),
    .B(_06416_),
    .Y(_06677_));
 sg13g2_o21ai_1 _16887_ (.B1(_06676_),
    .Y(_06678_),
    .A1(_06417_),
    .A2(_06677_));
 sg13g2_xnor2_1 _16888_ (.Y(_06679_),
    .A(_06455_),
    .B(_06458_));
 sg13g2_xnor2_1 _16889_ (.Y(_06680_),
    .A(_06462_),
    .B(_06679_));
 sg13g2_nor2_1 _16890_ (.A(_06472_),
    .B(_06478_),
    .Y(_06681_));
 sg13g2_xnor2_1 _16891_ (.Y(_06682_),
    .A(_06477_),
    .B(_06681_));
 sg13g2_nor2b_1 _16892_ (.A(_06680_),
    .B_N(_06682_),
    .Y(_06684_));
 sg13g2_nand2b_1 _16893_ (.Y(_06685_),
    .B(_06680_),
    .A_N(_06682_));
 sg13g2_xor2_1 _16894_ (.B(_06682_),
    .A(_06680_),
    .X(_06686_));
 sg13g2_xnor2_1 _16895_ (.Y(_06687_),
    .A(_06678_),
    .B(_06686_));
 sg13g2_nand2_1 _16896_ (.Y(_06688_),
    .A(_06675_),
    .B(_06687_));
 sg13g2_xor2_1 _16897_ (.B(_06498_),
    .A(_06495_),
    .X(_06689_));
 sg13g2_xnor2_1 _16898_ (.Y(_06690_),
    .A(_06501_),
    .B(_06689_));
 sg13g2_xor2_1 _16899_ (.B(_06509_),
    .A(_06505_),
    .X(_06691_));
 sg13g2_xnor2_1 _16900_ (.Y(_06692_),
    .A(_06510_),
    .B(_06691_));
 sg13g2_nand2_1 _16901_ (.Y(_06693_),
    .A(_06690_),
    .B(_06692_));
 sg13g2_or2_1 _16902_ (.X(_06695_),
    .B(_06692_),
    .A(_06690_));
 sg13g2_nand2_1 _16903_ (.Y(_06696_),
    .A(_06693_),
    .B(_06695_));
 sg13g2_nand2_1 _16904_ (.Y(_06697_),
    .A(_06536_),
    .B(_06541_));
 sg13g2_xor2_1 _16905_ (.B(_06697_),
    .A(_06539_),
    .X(_06698_));
 sg13g2_xnor2_1 _16906_ (.Y(_06699_),
    .A(_06696_),
    .B(_06698_));
 sg13g2_o21ai_1 _16907_ (.B1(_06699_),
    .Y(_06700_),
    .A1(_06675_),
    .A2(_06687_));
 sg13g2_a22oi_1 _16908_ (.Y(_06701_),
    .B1(_06688_),
    .B2(_06700_),
    .A2(_06665_),
    .A1(_06651_));
 sg13g2_and4_1 _16909_ (.A(_06651_),
    .B(_06665_),
    .C(_06688_),
    .D(_06700_),
    .X(_06702_));
 sg13g2_xnor2_1 _16910_ (.Y(_06703_),
    .A(_06577_),
    .B(_06578_));
 sg13g2_xnor2_1 _16911_ (.Y(_06704_),
    .A(_06582_),
    .B(_06703_));
 sg13g2_nor2b_1 _16912_ (.A(_06568_),
    .B_N(_06571_),
    .Y(_06706_));
 sg13g2_xnor2_1 _16913_ (.Y(_06707_),
    .A(_06570_),
    .B(_06706_));
 sg13g2_inv_1 _16914_ (.Y(_06708_),
    .A(_06707_));
 sg13g2_nand2b_1 _16915_ (.Y(_06709_),
    .B(_06707_),
    .A_N(_06704_));
 sg13g2_nand2_1 _16916_ (.Y(_06710_),
    .A(_06704_),
    .B(_06708_));
 sg13g2_xnor2_1 _16917_ (.Y(_06711_),
    .A(_06704_),
    .B(_06707_));
 sg13g2_xnor2_1 _16918_ (.Y(_06712_),
    .A(_06591_),
    .B(_06593_));
 sg13g2_xnor2_1 _16919_ (.Y(_06713_),
    .A(_06596_),
    .B(_06712_));
 sg13g2_xnor2_1 _16920_ (.Y(_06714_),
    .A(_06711_),
    .B(_06713_));
 sg13g2_xor2_1 _16921_ (.B(_06524_),
    .A(_06521_),
    .X(_06715_));
 sg13g2_xnor2_1 _16922_ (.Y(_06717_),
    .A(_06528_),
    .B(_06715_));
 sg13g2_xor2_1 _16923_ (.B(_06548_),
    .A(_06545_),
    .X(_06718_));
 sg13g2_xnor2_1 _16924_ (.Y(_06719_),
    .A(_06552_),
    .B(_06718_));
 sg13g2_nand2_1 _16925_ (.Y(_06720_),
    .A(_06717_),
    .B(_06719_));
 sg13g2_nor2_1 _16926_ (.A(_06717_),
    .B(_06719_),
    .Y(_06721_));
 sg13g2_xor2_1 _16927_ (.B(_06719_),
    .A(_06717_),
    .X(_06722_));
 sg13g2_nand2_1 _16928_ (.Y(_06723_),
    .A(_06559_),
    .B(_06564_));
 sg13g2_xor2_1 _16929_ (.B(_06723_),
    .A(_06563_),
    .X(_06724_));
 sg13g2_xnor2_1 _16930_ (.Y(_06725_),
    .A(_06722_),
    .B(_06724_));
 sg13g2_nor2_1 _16931_ (.A(_06714_),
    .B(_06725_),
    .Y(_06726_));
 sg13g2_and2_1 _16932_ (.A(_06714_),
    .B(_06725_),
    .X(_06728_));
 sg13g2_inv_1 _16933_ (.Y(_06729_),
    .A(_06728_));
 sg13g2_xor2_1 _16934_ (.B(_06603_),
    .A(_06600_),
    .X(_06730_));
 sg13g2_xnor2_1 _16935_ (.Y(_06731_),
    .A(_06607_),
    .B(_06730_));
 sg13g2_nor2_1 _16936_ (.A(_06616_),
    .B(_06620_),
    .Y(_06732_));
 sg13g2_xor2_1 _16937_ (.B(_06732_),
    .A(_06619_),
    .X(_06733_));
 sg13g2_nand2_1 _16938_ (.Y(_06734_),
    .A(_06731_),
    .B(_06733_));
 sg13g2_or2_1 _16939_ (.X(_06735_),
    .B(_06733_),
    .A(_06731_));
 sg13g2_nand2_1 _16940_ (.Y(_06736_),
    .A(_06734_),
    .B(_06735_));
 sg13g2_xnor2_1 _16941_ (.Y(_06737_),
    .A(net2405),
    .B(net2251));
 sg13g2_xnor2_1 _16942_ (.Y(_06739_),
    .A(net2323),
    .B(net2217));
 sg13g2_nand2_2 _16943_ (.Y(_06740_),
    .A(_06737_),
    .B(_06739_));
 sg13g2_xor2_1 _16944_ (.B(net2486),
    .A(net2523),
    .X(_06741_));
 sg13g2_nor2b_1 _16945_ (.A(net2443),
    .B_N(net2657),
    .Y(_06742_));
 sg13g2_nor2_1 _16946_ (.A(_05297_),
    .B(net2657),
    .Y(_06743_));
 sg13g2_nor4_2 _16947_ (.A(net2817),
    .B(\net.in[49] ),
    .C(_06742_),
    .Y(_06744_),
    .D(_06743_));
 sg13g2_nand2_1 _16948_ (.Y(_06745_),
    .A(_06741_),
    .B(_06744_));
 sg13g2_or2_1 _16949_ (.X(_06746_),
    .B(_06744_),
    .A(_06741_));
 sg13g2_nand2_1 _16950_ (.Y(_06747_),
    .A(_06745_),
    .B(_06746_));
 sg13g2_xnor2_1 _16951_ (.Y(_06748_),
    .A(_06740_),
    .B(_06747_));
 sg13g2_xnor2_1 _16952_ (.Y(_06750_),
    .A(_06736_),
    .B(_06748_));
 sg13g2_a21oi_2 _16953_ (.B1(_06726_),
    .Y(_06751_),
    .A2(_06750_),
    .A1(_06729_));
 sg13g2_nor2b_1 _16954_ (.A(_06702_),
    .B_N(_06751_),
    .Y(_06752_));
 sg13g2_nor2b_1 _16955_ (.A(net2651),
    .B_N(net2302),
    .Y(_06753_));
 sg13g2_or3_2 _16956_ (.A(\net.in[145] ),
    .B(net2310),
    .C(_06753_),
    .X(_06754_));
 sg13g2_nor2b_1 _16957_ (.A(net2812),
    .B_N(net2802),
    .Y(_06755_));
 sg13g2_nor2b_1 _16958_ (.A(net2802),
    .B_N(net2812),
    .Y(_06756_));
 sg13g2_nor2b_1 _16959_ (.A(net2513),
    .B_N(net2266),
    .Y(_06757_));
 sg13g2_nor3_2 _16960_ (.A(_06755_),
    .B(_06756_),
    .C(_06757_),
    .Y(_06758_));
 sg13g2_nand2b_1 _16961_ (.Y(_06759_),
    .B(net2552),
    .A_N(net2209));
 sg13g2_xnor2_1 _16962_ (.Y(_06761_),
    .A(net2371),
    .B(net2365));
 sg13g2_xnor2_1 _16963_ (.Y(_06762_),
    .A(_06759_),
    .B(_06761_));
 sg13g2_nand2b_1 _16964_ (.Y(_06763_),
    .B(_06758_),
    .A_N(_06762_));
 sg13g2_nor2b_1 _16965_ (.A(_06758_),
    .B_N(_06762_),
    .Y(_06764_));
 sg13g2_xnor2_1 _16966_ (.Y(_06765_),
    .A(_06758_),
    .B(_06762_));
 sg13g2_xnor2_1 _16967_ (.Y(_06766_),
    .A(_06754_),
    .B(_06765_));
 sg13g2_nand2_1 _16968_ (.Y(_06767_),
    .A(net2683),
    .B(\net.in[191] ));
 sg13g2_o21ai_1 _16969_ (.B1(_06767_),
    .Y(_06768_),
    .A1(net2586),
    .A2(net2544));
 sg13g2_a21oi_2 _16970_ (.B1(_06768_),
    .Y(_06769_),
    .A2(net2544),
    .A1(net2586));
 sg13g2_nand2b_1 _16971_ (.Y(_06770_),
    .B(net2305),
    .A_N(net2488));
 sg13g2_nand2b_1 _16972_ (.Y(_06772_),
    .B(net2488),
    .A_N(net2304));
 sg13g2_nand4_1 _16973_ (.B(net2618),
    .C(_06770_),
    .A(_05253_),
    .Y(_06773_),
    .D(_06772_));
 sg13g2_nor2_1 _16974_ (.A(_02317_),
    .B(_06537_),
    .Y(_06774_));
 sg13g2_nor2b_1 _16975_ (.A(_06773_),
    .B_N(_06774_),
    .Y(_06775_));
 sg13g2_o21ai_1 _16976_ (.B1(_06773_),
    .Y(_06776_),
    .A1(_02317_),
    .A2(_06537_));
 sg13g2_xor2_1 _16977_ (.B(_06774_),
    .A(_06773_),
    .X(_06777_));
 sg13g2_o21ai_1 _16978_ (.B1(_06776_),
    .Y(_06778_),
    .A1(_06769_),
    .A2(_06775_));
 sg13g2_xnor2_1 _16979_ (.Y(_06779_),
    .A(_06769_),
    .B(_06777_));
 sg13g2_nand2_1 _16980_ (.Y(_06780_),
    .A(_06766_),
    .B(_06779_));
 sg13g2_xnor2_1 _16981_ (.Y(_06781_),
    .A(_06766_),
    .B(_06779_));
 sg13g2_nor2_1 _16982_ (.A(net2601),
    .B(net2208),
    .Y(_06783_));
 sg13g2_xor2_1 _16983_ (.B(_06783_),
    .A(_05874_),
    .X(_06784_));
 sg13g2_nor2_1 _16984_ (.A(net2412),
    .B(net2370),
    .Y(_06785_));
 sg13g2_xnor2_1 _16985_ (.Y(_06786_),
    .A(net2502),
    .B(_06785_));
 sg13g2_xnor2_1 _16986_ (.Y(_06787_),
    .A(net2283),
    .B(net2409));
 sg13g2_xnor2_1 _16987_ (.Y(_06788_),
    .A(net2218),
    .B(_06787_));
 sg13g2_inv_1 _16988_ (.Y(_06789_),
    .A(_06788_));
 sg13g2_nand2_1 _16989_ (.Y(_06790_),
    .A(_06786_),
    .B(_06789_));
 sg13g2_nor2_1 _16990_ (.A(_06786_),
    .B(_06789_),
    .Y(_06791_));
 sg13g2_xnor2_1 _16991_ (.Y(_06792_),
    .A(_06786_),
    .B(_06788_));
 sg13g2_xnor2_1 _16992_ (.Y(_06794_),
    .A(_06784_),
    .B(_06792_));
 sg13g2_xnor2_1 _16993_ (.Y(_06795_),
    .A(_06781_),
    .B(_06794_));
 sg13g2_xor2_1 _16994_ (.B(_06294_),
    .A(_06283_),
    .X(_06796_));
 sg13g2_xnor2_1 _16995_ (.Y(_06797_),
    .A(_06308_),
    .B(_06796_));
 sg13g2_nand2_1 _16996_ (.Y(_06798_),
    .A(_06795_),
    .B(_06797_));
 sg13g2_xnor2_1 _16997_ (.Y(_06799_),
    .A(net2283),
    .B(net2363));
 sg13g2_xnor2_1 _16998_ (.Y(_06800_),
    .A(net2218),
    .B(_06799_));
 sg13g2_or2_1 _16999_ (.X(_06801_),
    .B(_06797_),
    .A(_06795_));
 sg13g2_nand2_1 _17000_ (.Y(_06802_),
    .A(_06798_),
    .B(_06800_));
 sg13g2_xor2_1 _17001_ (.B(net2360),
    .A(net2405),
    .X(_06803_));
 sg13g2_xnor2_1 _17002_ (.Y(_06805_),
    .A(_02357_),
    .B(_06803_));
 sg13g2_nor2b_1 _17003_ (.A(net2473),
    .B_N(net2197),
    .Y(_06806_));
 sg13g2_nor3_2 _17004_ (.A(net2390),
    .B(net2342),
    .C(_06806_),
    .Y(_06807_));
 sg13g2_nor2_1 _17005_ (.A(net2382),
    .B(net2812),
    .Y(_06808_));
 sg13g2_xor2_1 _17006_ (.B(net2747),
    .A(net2414),
    .X(_06809_));
 sg13g2_xnor2_1 _17007_ (.Y(_06810_),
    .A(_06808_),
    .B(_06809_));
 sg13g2_nor2b_1 _17008_ (.A(_06810_),
    .B_N(_06807_),
    .Y(_06811_));
 sg13g2_nand2b_1 _17009_ (.Y(_06812_),
    .B(_06810_),
    .A_N(_06807_));
 sg13g2_xor2_1 _17010_ (.B(_06810_),
    .A(_06807_),
    .X(_06813_));
 sg13g2_xnor2_1 _17011_ (.Y(_06814_),
    .A(_06805_),
    .B(_06813_));
 sg13g2_nor2_1 _17012_ (.A(net2467),
    .B(net2361),
    .Y(_06816_));
 sg13g2_nor3_2 _17013_ (.A(net2336),
    .B(net2350),
    .C(_06816_),
    .Y(_06817_));
 sg13g2_xor2_1 _17014_ (.B(net2600),
    .A(net2646),
    .X(_06818_));
 sg13g2_xnor2_1 _17015_ (.Y(_06819_),
    .A(net2483),
    .B(net2397));
 sg13g2_xnor2_1 _17016_ (.Y(_06820_),
    .A(_00766_),
    .B(_06819_));
 sg13g2_inv_1 _17017_ (.Y(_06821_),
    .A(_06820_));
 sg13g2_nand2_1 _17018_ (.Y(_06822_),
    .A(_06818_),
    .B(_06821_));
 sg13g2_xnor2_1 _17019_ (.Y(_06823_),
    .A(_06818_),
    .B(_06820_));
 sg13g2_xnor2_1 _17020_ (.Y(_06824_),
    .A(_06817_),
    .B(_06823_));
 sg13g2_nand2b_1 _17021_ (.Y(_06825_),
    .B(_06814_),
    .A_N(_06824_));
 sg13g2_nand2b_1 _17022_ (.Y(_06827_),
    .B(_06824_),
    .A_N(_06814_));
 sg13g2_xnor2_1 _17023_ (.Y(_06828_),
    .A(_06814_),
    .B(_06824_));
 sg13g2_xor2_1 _17024_ (.B(net2291),
    .A(net2354),
    .X(_06829_));
 sg13g2_nand2b_1 _17025_ (.Y(_06830_),
    .B(net2222),
    .A_N(net2272));
 sg13g2_nor2_1 _17026_ (.A(net2526),
    .B(net2642),
    .Y(_06831_));
 sg13g2_xnor2_1 _17027_ (.Y(_06832_),
    .A(_06830_),
    .B(_06831_));
 sg13g2_nand2b_1 _17028_ (.Y(_06833_),
    .B(net2376),
    .A_N(net2359));
 sg13g2_nor2b_1 _17029_ (.A(net2381),
    .B_N(net2506),
    .Y(_06834_));
 sg13g2_xnor2_1 _17030_ (.Y(_06835_),
    .A(_06833_),
    .B(_06834_));
 sg13g2_nand2_1 _17031_ (.Y(_06836_),
    .A(_06832_),
    .B(_06835_));
 sg13g2_or2_1 _17032_ (.X(_06838_),
    .B(_06835_),
    .A(_06832_));
 sg13g2_nand2_1 _17033_ (.Y(_06839_),
    .A(_06836_),
    .B(_06838_));
 sg13g2_xor2_1 _17034_ (.B(_06839_),
    .A(_06829_),
    .X(_06840_));
 sg13g2_xnor2_1 _17035_ (.Y(_06841_),
    .A(_06828_),
    .B(_06840_));
 sg13g2_nor2_1 _17036_ (.A(net2357),
    .B(net2403),
    .Y(_06842_));
 sg13g2_o21ai_1 _17037_ (.B1(_06842_),
    .Y(_06843_),
    .A1(net2480),
    .A2(net2395));
 sg13g2_a21oi_2 _17038_ (.B1(_06843_),
    .Y(_06844_),
    .A2(net2395),
    .A1(net2480));
 sg13g2_xnor2_1 _17039_ (.Y(_06845_),
    .A(net2660),
    .B(net2544));
 sg13g2_nand2_1 _17040_ (.Y(_06846_),
    .A(net2247),
    .B(\net.in[188] ));
 sg13g2_o21ai_1 _17041_ (.B1(_06846_),
    .Y(_06847_),
    .A1(\net.in[188] ),
    .A2(_02057_));
 sg13g2_nand2b_1 _17042_ (.Y(_06849_),
    .B(_06847_),
    .A_N(_06845_));
 sg13g2_nand2b_1 _17043_ (.Y(_06850_),
    .B(_06845_),
    .A_N(_06847_));
 sg13g2_xnor2_1 _17044_ (.Y(_06851_),
    .A(_06845_),
    .B(_06847_));
 sg13g2_xnor2_1 _17045_ (.Y(_06852_),
    .A(_06844_),
    .B(_06851_));
 sg13g2_xnor2_1 _17046_ (.Y(_06853_),
    .A(net2390),
    .B(net2188));
 sg13g2_mux2_2 _17047_ (.A0(net2241),
    .A1(_06317_),
    .S(_05253_),
    .X(_06854_));
 sg13g2_nor2b_1 _17048_ (.A(net2521),
    .B_N(net2592),
    .Y(_06855_));
 sg13g2_xnor2_1 _17049_ (.Y(_06856_),
    .A(net2200),
    .B(net2600));
 sg13g2_xnor2_1 _17050_ (.Y(_06857_),
    .A(_06855_),
    .B(_06856_));
 sg13g2_nand2_1 _17051_ (.Y(_06858_),
    .A(_06854_),
    .B(_06857_));
 sg13g2_xor2_1 _17052_ (.B(_06857_),
    .A(_06854_),
    .X(_06860_));
 sg13g2_xnor2_1 _17053_ (.Y(_06861_),
    .A(_06853_),
    .B(_06860_));
 sg13g2_nand2_1 _17054_ (.Y(_06862_),
    .A(_06852_),
    .B(_06861_));
 sg13g2_xnor2_1 _17055_ (.Y(_06863_),
    .A(net2376),
    .B(net2254));
 sg13g2_xor2_1 _17056_ (.B(net2281),
    .A(net2217),
    .X(_06864_));
 sg13g2_nor2_1 _17057_ (.A(net2687),
    .B(net2630),
    .Y(_06865_));
 sg13g2_xnor2_1 _17058_ (.Y(_06866_),
    .A(net2696),
    .B(net2812));
 sg13g2_xnor2_1 _17059_ (.Y(_06867_),
    .A(_06865_),
    .B(_06866_));
 sg13g2_o21ai_1 _17060_ (.B1(_06867_),
    .Y(_06868_),
    .A1(_07486_),
    .A2(_06864_));
 sg13g2_or3_1 _17061_ (.A(_07486_),
    .B(_06864_),
    .C(_06867_),
    .X(_06869_));
 sg13g2_nand2_1 _17062_ (.Y(_06871_),
    .A(_06868_),
    .B(_06869_));
 sg13g2_xor2_1 _17063_ (.B(_06871_),
    .A(_06863_),
    .X(_06872_));
 sg13g2_o21ai_1 _17064_ (.B1(_06872_),
    .Y(_06873_),
    .A1(_06852_),
    .A2(_06861_));
 sg13g2_xnor2_1 _17065_ (.Y(_06874_),
    .A(_06852_),
    .B(_06861_));
 sg13g2_xnor2_1 _17066_ (.Y(_06875_),
    .A(_06872_),
    .B(_06874_));
 sg13g2_nand2_1 _17067_ (.Y(_06876_),
    .A(_06841_),
    .B(_06875_));
 sg13g2_or2_1 _17068_ (.X(_06877_),
    .B(_06875_),
    .A(_06841_));
 sg13g2_nor2_1 _17069_ (.A(net2280),
    .B(net2316),
    .Y(_06878_));
 sg13g2_nor2_2 _17070_ (.A(net2452),
    .B(net2213),
    .Y(_06879_));
 sg13g2_xnor2_1 _17071_ (.Y(_06880_),
    .A(_06878_),
    .B(_06879_));
 sg13g2_xnor2_1 _17072_ (.Y(_06882_),
    .A(net2236),
    .B(net2197));
 sg13g2_xnor2_1 _17073_ (.Y(_06883_),
    .A(net2426),
    .B(_06882_));
 sg13g2_xnor2_1 _17074_ (.Y(_06884_),
    .A(_06437_),
    .B(_06601_));
 sg13g2_nor2_1 _17075_ (.A(_06883_),
    .B(_06884_),
    .Y(_06885_));
 sg13g2_nand2_1 _17076_ (.Y(_06886_),
    .A(_06883_),
    .B(_06884_));
 sg13g2_nor2b_1 _17077_ (.A(_06885_),
    .B_N(_06886_),
    .Y(_06887_));
 sg13g2_xnor2_1 _17078_ (.Y(_06888_),
    .A(_06880_),
    .B(_06887_));
 sg13g2_nor2_1 _17079_ (.A(net2781),
    .B(\net.in[191] ),
    .Y(_06889_));
 sg13g2_xnor2_1 _17080_ (.Y(_06890_),
    .A(_06297_),
    .B(_06889_));
 sg13g2_nor2_1 _17081_ (.A(net2596),
    .B(net2639),
    .Y(_06891_));
 sg13g2_nor2_1 _17082_ (.A(net2586),
    .B(net2209),
    .Y(_06893_));
 sg13g2_xor2_1 _17083_ (.B(_06893_),
    .A(_06891_),
    .X(_06894_));
 sg13g2_nor2_1 _17084_ (.A(net2809),
    .B(net2370),
    .Y(_06895_));
 sg13g2_nand2b_1 _17085_ (.Y(_06896_),
    .B(net2467),
    .A_N(net2409));
 sg13g2_xnor2_1 _17086_ (.Y(_06897_),
    .A(_06895_),
    .B(_06896_));
 sg13g2_nand2_1 _17087_ (.Y(_06898_),
    .A(_06894_),
    .B(_06897_));
 sg13g2_or2_1 _17088_ (.X(_06899_),
    .B(_06897_),
    .A(_06894_));
 sg13g2_nand2_1 _17089_ (.Y(_06900_),
    .A(_06898_),
    .B(_06899_));
 sg13g2_xor2_1 _17090_ (.B(_06900_),
    .A(_06890_),
    .X(_06901_));
 sg13g2_or2_1 _17091_ (.X(_06902_),
    .B(_06901_),
    .A(_06888_));
 sg13g2_nand2_1 _17092_ (.Y(_06904_),
    .A(_06888_),
    .B(_06901_));
 sg13g2_nand2_1 _17093_ (.Y(_06905_),
    .A(_06902_),
    .B(_06904_));
 sg13g2_nand2b_1 _17094_ (.Y(_06906_),
    .B(\net.in[222] ),
    .A_N(net2704));
 sg13g2_o21ai_1 _17095_ (.B1(_06906_),
    .Y(_06907_),
    .A1(_05121_),
    .A2(net2207));
 sg13g2_a21oi_2 _17096_ (.B1(_06907_),
    .Y(_06908_),
    .A2(net2704),
    .A1(_06067_));
 sg13g2_nor2_2 _17097_ (.A(net2277),
    .B(_05968_),
    .Y(_06909_));
 sg13g2_xnor2_1 _17098_ (.Y(_06910_),
    .A(net2405),
    .B(_06909_));
 sg13g2_xor2_1 _17099_ (.B(net2221),
    .A(net2371),
    .X(_06911_));
 sg13g2_nor2_1 _17100_ (.A(_06910_),
    .B(_06911_),
    .Y(_06912_));
 sg13g2_nand2_1 _17101_ (.Y(_06913_),
    .A(_06910_),
    .B(_06911_));
 sg13g2_nand2b_1 _17102_ (.Y(_06915_),
    .B(_06913_),
    .A_N(_06912_));
 sg13g2_xnor2_1 _17103_ (.Y(_06916_),
    .A(_06908_),
    .B(_06915_));
 sg13g2_xor2_1 _17104_ (.B(_06916_),
    .A(_06905_),
    .X(_06917_));
 sg13g2_nand2_1 _17105_ (.Y(_06918_),
    .A(_06877_),
    .B(_06917_));
 sg13g2_and4_1 _17106_ (.A(_06801_),
    .B(_06802_),
    .C(_06876_),
    .D(_06918_),
    .X(_06919_));
 sg13g2_inv_1 _17107_ (.Y(_06920_),
    .A(_06919_));
 sg13g2_a22oi_1 _17108_ (.Y(_06921_),
    .B1(_06876_),
    .B2(_06918_),
    .A2(_06802_),
    .A1(_06801_));
 sg13g2_o21ai_1 _17109_ (.B1(_06644_),
    .Y(_06922_),
    .A1(_06643_),
    .A2(_06647_));
 sg13g2_a21oi_2 _17110_ (.B1(_06921_),
    .Y(_06923_),
    .A2(_06922_),
    .A1(_06920_));
 sg13g2_o21ai_1 _17111_ (.B1(_06923_),
    .Y(_06924_),
    .A1(_06701_),
    .A2(_06752_));
 sg13g2_nand2_1 _17112_ (.Y(_06926_),
    .A(_06633_),
    .B(_06636_));
 sg13g2_a21oi_1 _17113_ (.A1(_06632_),
    .A2(_06926_),
    .Y(_06927_),
    .B1(_06663_));
 sg13g2_a21o_1 _17114_ (.A2(_06685_),
    .A1(_06678_),
    .B1(_06684_),
    .X(_06928_));
 sg13g2_and3_1 _17115_ (.X(_06929_),
    .A(_06632_),
    .B(_06663_),
    .C(_06926_));
 sg13g2_nor2_1 _17116_ (.A(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sg13g2_nor2_1 _17117_ (.A(_06927_),
    .B(_06930_),
    .Y(_06931_));
 sg13g2_inv_1 _17118_ (.Y(_06932_),
    .A(_06931_));
 sg13g2_or3_1 _17119_ (.A(_06701_),
    .B(_06752_),
    .C(_06923_),
    .X(_06933_));
 sg13g2_nand2_1 _17120_ (.Y(_06934_),
    .A(_06924_),
    .B(_06932_));
 sg13g2_nand2_2 _17121_ (.Y(_06935_),
    .A(_06933_),
    .B(_06934_));
 sg13g2_o21ai_1 _17122_ (.B1(_06886_),
    .Y(_06937_),
    .A1(_06880_),
    .A2(_06885_));
 sg13g2_nand2_1 _17123_ (.Y(_06938_),
    .A(_06829_),
    .B(_06836_));
 sg13g2_nand2b_1 _17124_ (.Y(_06939_),
    .B(_06898_),
    .A_N(_06890_));
 sg13g2_and4_1 _17125_ (.A(_06838_),
    .B(_06899_),
    .C(_06938_),
    .D(_06939_),
    .X(_06940_));
 sg13g2_inv_1 _17126_ (.Y(_06941_),
    .A(_06940_));
 sg13g2_a22oi_1 _17127_ (.Y(_06942_),
    .B1(_06939_),
    .B2(_06899_),
    .A2(_06938_),
    .A1(_06838_));
 sg13g2_nor2_1 _17128_ (.A(_06940_),
    .B(_06942_),
    .Y(_06943_));
 sg13g2_xnor2_1 _17129_ (.Y(_06944_),
    .A(_06937_),
    .B(_06943_));
 sg13g2_o21ai_1 _17130_ (.B1(_06913_),
    .Y(_06945_),
    .A1(_06908_),
    .A2(_06912_));
 sg13g2_a21o_1 _17131_ (.A2(_06763_),
    .A1(_06754_),
    .B1(_06764_),
    .X(_06946_));
 sg13g2_xor2_1 _17132_ (.B(_06946_),
    .A(_06945_),
    .X(_06948_));
 sg13g2_xnor2_1 _17133_ (.Y(_06949_),
    .A(_06778_),
    .B(_06948_));
 sg13g2_nand2_1 _17134_ (.Y(_06950_),
    .A(_06944_),
    .B(_06949_));
 sg13g2_nor2_1 _17135_ (.A(_06944_),
    .B(_06949_),
    .Y(_06951_));
 sg13g2_a21oi_2 _17136_ (.B1(_06281_),
    .Y(_06952_),
    .A2(_06280_),
    .A1(_06272_));
 sg13g2_o21ai_1 _17137_ (.B1(_06790_),
    .Y(_06953_),
    .A1(_06784_),
    .A2(_06791_));
 sg13g2_a21oi_2 _17138_ (.B1(_06292_),
    .Y(_06954_),
    .A2(_06291_),
    .A1(_06284_));
 sg13g2_xor2_1 _17139_ (.B(_06954_),
    .A(_06953_),
    .X(_06955_));
 sg13g2_a21o_1 _17140_ (.A2(_06954_),
    .A1(_06953_),
    .B1(_06952_),
    .X(_06956_));
 sg13g2_o21ai_1 _17141_ (.B1(_06956_),
    .Y(_06957_),
    .A1(_06953_),
    .A2(_06954_));
 sg13g2_xnor2_1 _17142_ (.Y(_06959_),
    .A(_06952_),
    .B(_06955_));
 sg13g2_a21oi_1 _17143_ (.A1(_06950_),
    .A2(_06959_),
    .Y(_06960_),
    .B1(_06951_));
 sg13g2_xor2_1 _17144_ (.B(_06609_),
    .A(_06598_),
    .X(_06961_));
 sg13g2_xnor2_1 _17145_ (.Y(_06962_),
    .A(_06621_),
    .B(_06961_));
 sg13g2_o21ai_1 _17146_ (.B1(_06853_),
    .Y(_06963_),
    .A1(_06854_),
    .A2(_06857_));
 sg13g2_nand2_1 _17147_ (.Y(_06964_),
    .A(_06858_),
    .B(_06963_));
 sg13g2_nand2_1 _17148_ (.Y(_06965_),
    .A(_06740_),
    .B(_06745_));
 sg13g2_nand2b_1 _17149_ (.Y(_06966_),
    .B(_06849_),
    .A_N(_06844_));
 sg13g2_and4_1 _17150_ (.A(_06746_),
    .B(_06850_),
    .C(_06965_),
    .D(_06966_),
    .X(_06967_));
 sg13g2_a22oi_1 _17151_ (.Y(_06968_),
    .B1(_06966_),
    .B2(_06850_),
    .A2(_06965_),
    .A1(_06746_));
 sg13g2_inv_1 _17152_ (.Y(_06970_),
    .A(_06968_));
 sg13g2_o21ai_1 _17153_ (.B1(_06970_),
    .Y(_06971_),
    .A1(_06964_),
    .A2(_06967_));
 sg13g2_a21o_1 _17154_ (.A2(_06967_),
    .A1(_06964_),
    .B1(_06971_),
    .X(_06972_));
 sg13g2_o21ai_1 _17155_ (.B1(_06972_),
    .Y(_06973_),
    .A1(_06964_),
    .A2(_06970_));
 sg13g2_nor2_1 _17156_ (.A(_06962_),
    .B(_06973_),
    .Y(_06974_));
 sg13g2_and2_1 _17157_ (.A(_06962_),
    .B(_06973_),
    .X(_06975_));
 sg13g2_o21ai_1 _17158_ (.B1(_06812_),
    .Y(_06976_),
    .A1(_06805_),
    .A2(_06811_));
 sg13g2_nand2_1 _17159_ (.Y(_06977_),
    .A(_06863_),
    .B(_06868_));
 sg13g2_o21ai_1 _17160_ (.B1(_06817_),
    .Y(_06978_),
    .A1(_06818_),
    .A2(_06821_));
 sg13g2_and4_1 _17161_ (.A(_06822_),
    .B(_06869_),
    .C(_06977_),
    .D(_06978_),
    .X(_06979_));
 sg13g2_a22oi_1 _17162_ (.Y(_06981_),
    .B1(_06978_),
    .B2(_06822_),
    .A2(_06977_),
    .A1(_06869_));
 sg13g2_nor2_1 _17163_ (.A(_06979_),
    .B(_06981_),
    .Y(_06982_));
 sg13g2_xnor2_1 _17164_ (.Y(_06983_),
    .A(_06976_),
    .B(_06982_));
 sg13g2_nor2_1 _17165_ (.A(_06974_),
    .B(_06983_),
    .Y(_06984_));
 sg13g2_nor2_1 _17166_ (.A(_06975_),
    .B(_06984_),
    .Y(_06985_));
 sg13g2_nand2_1 _17167_ (.Y(_06986_),
    .A(_06960_),
    .B(_06985_));
 sg13g2_nand2_1 _17168_ (.Y(_06987_),
    .A(_06798_),
    .B(_06801_));
 sg13g2_xor2_1 _17169_ (.B(_06987_),
    .A(_06800_),
    .X(_06988_));
 sg13g2_nand2_1 _17170_ (.Y(_06989_),
    .A(_06876_),
    .B(_06877_));
 sg13g2_xor2_1 _17171_ (.B(_06989_),
    .A(_06917_),
    .X(_06990_));
 sg13g2_nor2_1 _17172_ (.A(_06988_),
    .B(_06990_),
    .Y(_06992_));
 sg13g2_nand2_1 _17173_ (.Y(_06993_),
    .A(_06988_),
    .B(_06990_));
 sg13g2_nand2b_1 _17174_ (.Y(_06994_),
    .B(_06993_),
    .A_N(_06992_));
 sg13g2_xnor2_1 _17175_ (.Y(_06995_),
    .A(_06637_),
    .B(_06648_));
 sg13g2_xnor2_1 _17176_ (.Y(_06996_),
    .A(_06664_),
    .B(_06995_));
 sg13g2_xor2_1 _17177_ (.B(_06687_),
    .A(_06675_),
    .X(_06997_));
 sg13g2_xnor2_1 _17178_ (.Y(_06998_),
    .A(_06699_),
    .B(_06997_));
 sg13g2_nand2_1 _17179_ (.Y(_06999_),
    .A(_06996_),
    .B(_06998_));
 sg13g2_nor2_1 _17180_ (.A(_06996_),
    .B(_06998_),
    .Y(_07000_));
 sg13g2_xor2_1 _17181_ (.B(_06998_),
    .A(_06996_),
    .X(_07001_));
 sg13g2_nor2_1 _17182_ (.A(_06726_),
    .B(_06728_),
    .Y(_07003_));
 sg13g2_xnor2_1 _17183_ (.Y(_07004_),
    .A(_06750_),
    .B(_07003_));
 sg13g2_xnor2_1 _17184_ (.Y(_07005_),
    .A(_07001_),
    .B(_07004_));
 sg13g2_a21oi_1 _17185_ (.A1(_06993_),
    .A2(_07005_),
    .Y(_07006_),
    .B1(_06992_));
 sg13g2_a21oi_2 _17186_ (.B1(_07000_),
    .Y(_07007_),
    .A2(_07004_),
    .A1(_06999_));
 sg13g2_nand2b_1 _17187_ (.Y(_07008_),
    .B(_07007_),
    .A_N(_07006_));
 sg13g2_or2_1 _17188_ (.X(_07009_),
    .B(_06985_),
    .A(_06960_));
 sg13g2_nand2_1 _17189_ (.Y(_07010_),
    .A(_07008_),
    .B(_07009_));
 sg13g2_and2_1 _17190_ (.A(_06986_),
    .B(_07010_),
    .X(_07011_));
 sg13g2_or2_1 _17191_ (.X(_07012_),
    .B(_07011_),
    .A(_06935_));
 sg13g2_and2_1 _17192_ (.A(_06935_),
    .B(_07011_),
    .X(_07014_));
 sg13g2_a21o_1 _17193_ (.A2(_06669_),
    .A1(_06667_),
    .B1(_06674_),
    .X(_07015_));
 sg13g2_nand2_1 _17194_ (.Y(_07016_),
    .A(_06695_),
    .B(_06698_));
 sg13g2_a22oi_1 _17195_ (.Y(_07017_),
    .B1(_07016_),
    .B2(_06693_),
    .A2(_07015_),
    .A1(_06670_));
 sg13g2_nand4_1 _17196_ (.B(_06693_),
    .C(_07015_),
    .A(_06670_),
    .Y(_07018_),
    .D(_07016_));
 sg13g2_o21ai_1 _17197_ (.B1(_06720_),
    .Y(_07019_),
    .A1(_06721_),
    .A2(_06724_));
 sg13g2_nand2_1 _17198_ (.Y(_07020_),
    .A(_07018_),
    .B(_07019_));
 sg13g2_nand2b_1 _17199_ (.Y(_07021_),
    .B(_07020_),
    .A_N(_07017_));
 sg13g2_nand2_1 _17200_ (.Y(_07022_),
    .A(_06735_),
    .B(_06748_));
 sg13g2_nand2_1 _17201_ (.Y(_07023_),
    .A(_06710_),
    .B(_06713_));
 sg13g2_and2_1 _17202_ (.A(_06709_),
    .B(_07023_),
    .X(_07025_));
 sg13g2_nand3_1 _17203_ (.B(_07022_),
    .C(_07025_),
    .A(_06734_),
    .Y(_07026_));
 sg13g2_nand2_2 _17204_ (.Y(_07027_),
    .A(_06862_),
    .B(_06873_));
 sg13g2_a21o_1 _17205_ (.A2(_07022_),
    .A1(_06734_),
    .B1(_07025_),
    .X(_07028_));
 sg13g2_nand2_1 _17206_ (.Y(_07029_),
    .A(_07026_),
    .B(_07027_));
 sg13g2_nand3_1 _17207_ (.B(_07028_),
    .C(_07029_),
    .A(_07021_),
    .Y(_07030_));
 sg13g2_inv_1 _17208_ (.Y(_07031_),
    .A(_07030_));
 sg13g2_a21o_1 _17209_ (.A2(_07029_),
    .A1(_07028_),
    .B1(_07021_),
    .X(_07032_));
 sg13g2_nand2_1 _17210_ (.Y(_07033_),
    .A(_06827_),
    .B(_06840_));
 sg13g2_nand2_1 _17211_ (.Y(_07034_),
    .A(_06904_),
    .B(_06916_));
 sg13g2_a22oi_1 _17212_ (.Y(_07036_),
    .B1(_07034_),
    .B2(_06902_),
    .A2(_07033_),
    .A1(_06825_));
 sg13g2_o21ai_1 _17213_ (.B1(_06794_),
    .Y(_07037_),
    .A1(_06766_),
    .A2(_06779_));
 sg13g2_nand2_1 _17214_ (.Y(_07038_),
    .A(_06780_),
    .B(_07037_));
 sg13g2_and4_1 _17215_ (.A(_06825_),
    .B(_06902_),
    .C(_07033_),
    .D(_07034_),
    .X(_07039_));
 sg13g2_nor2_1 _17216_ (.A(_07036_),
    .B(_07038_),
    .Y(_07040_));
 sg13g2_nor2_2 _17217_ (.A(_07039_),
    .B(_07040_),
    .Y(_07041_));
 sg13g2_o21ai_1 _17218_ (.B1(_07032_),
    .Y(_07042_),
    .A1(_07031_),
    .A2(_07041_));
 sg13g2_a21oi_2 _17219_ (.B1(_07014_),
    .Y(_07043_),
    .A2(_07042_),
    .A1(_07012_));
 sg13g2_xor2_1 _17220_ (.B(_07007_),
    .A(_07006_),
    .X(_07044_));
 sg13g2_nor2_1 _17221_ (.A(_06701_),
    .B(_06702_),
    .Y(_07045_));
 sg13g2_xnor2_1 _17222_ (.Y(_07047_),
    .A(_06751_),
    .B(_07045_));
 sg13g2_inv_1 _17223_ (.Y(_07048_),
    .A(_07047_));
 sg13g2_nand2b_1 _17224_ (.Y(_07049_),
    .B(_07047_),
    .A_N(_07044_));
 sg13g2_xnor2_1 _17225_ (.Y(_07050_),
    .A(_07044_),
    .B(_07048_));
 sg13g2_nor2_1 _17226_ (.A(_06919_),
    .B(_06921_),
    .Y(_07051_));
 sg13g2_xnor2_1 _17227_ (.Y(_07052_),
    .A(_06922_),
    .B(_07051_));
 sg13g2_xnor2_1 _17228_ (.Y(_07053_),
    .A(_07050_),
    .B(_07052_));
 sg13g2_nand2_1 _17229_ (.Y(_07054_),
    .A(_07026_),
    .B(_07028_));
 sg13g2_xor2_1 _17230_ (.B(_07054_),
    .A(_07027_),
    .X(_07055_));
 sg13g2_nor2b_1 _17231_ (.A(_07017_),
    .B_N(_07018_),
    .Y(_07056_));
 sg13g2_xnor2_1 _17232_ (.Y(_07058_),
    .A(_07019_),
    .B(_07056_));
 sg13g2_nor2_1 _17233_ (.A(_06927_),
    .B(_06929_),
    .Y(_07059_));
 sg13g2_xnor2_1 _17234_ (.Y(_07060_),
    .A(_06928_),
    .B(_07059_));
 sg13g2_nand2_1 _17235_ (.Y(_07061_),
    .A(_07058_),
    .B(_07060_));
 sg13g2_or2_1 _17236_ (.X(_07062_),
    .B(_07060_),
    .A(_07058_));
 sg13g2_nand2_1 _17237_ (.Y(_07063_),
    .A(_07061_),
    .B(_07062_));
 sg13g2_nand2_1 _17238_ (.Y(_07064_),
    .A(_07055_),
    .B(_07061_));
 sg13g2_nand2_1 _17239_ (.Y(_07065_),
    .A(_07062_),
    .B(_07064_));
 sg13g2_inv_1 _17240_ (.Y(_07066_),
    .A(_07065_));
 sg13g2_xor2_1 _17241_ (.B(_07063_),
    .A(_07055_),
    .X(_07067_));
 sg13g2_nand2b_1 _17242_ (.Y(_07069_),
    .B(_07067_),
    .A_N(_07053_));
 sg13g2_nor2b_1 _17243_ (.A(_07067_),
    .B_N(_07053_),
    .Y(_07070_));
 sg13g2_xnor2_1 _17244_ (.Y(_07071_),
    .A(_07053_),
    .B(_07067_));
 sg13g2_nor2_1 _17245_ (.A(_06323_),
    .B(_06332_),
    .Y(_07072_));
 sg13g2_xnor2_1 _17246_ (.Y(_07073_),
    .A(_06330_),
    .B(_07072_));
 sg13g2_nor2_1 _17247_ (.A(_07036_),
    .B(_07039_),
    .Y(_07074_));
 sg13g2_xnor2_1 _17248_ (.Y(_07075_),
    .A(_07038_),
    .B(_07074_));
 sg13g2_nand2b_1 _17249_ (.Y(_07076_),
    .B(_07073_),
    .A_N(_07075_));
 sg13g2_nor2b_1 _17250_ (.A(_07073_),
    .B_N(_07075_),
    .Y(_07077_));
 sg13g2_xnor2_1 _17251_ (.Y(_07078_),
    .A(_07073_),
    .B(_07075_));
 sg13g2_xnor2_1 _17252_ (.Y(_07080_),
    .A(_06345_),
    .B(_06352_));
 sg13g2_xnor2_1 _17253_ (.Y(_07081_),
    .A(_06365_),
    .B(_07080_));
 sg13g2_xnor2_1 _17254_ (.Y(_07082_),
    .A(_07078_),
    .B(_07081_));
 sg13g2_xnor2_1 _17255_ (.Y(_07083_),
    .A(_07071_),
    .B(_07082_));
 sg13g2_nand2b_1 _17256_ (.Y(_07084_),
    .B(_06575_),
    .A_N(_06574_));
 sg13g2_xnor2_1 _17257_ (.Y(_07085_),
    .A(_06585_),
    .B(_07084_));
 sg13g2_xnor2_1 _17258_ (.Y(_07086_),
    .A(_06492_),
    .B(_06503_));
 sg13g2_xnor2_1 _17259_ (.Y(_07087_),
    .A(_06513_),
    .B(_07086_));
 sg13g2_nor2b_1 _17260_ (.A(_06543_),
    .B_N(_06544_),
    .Y(_07088_));
 sg13g2_xnor2_1 _17261_ (.Y(_07089_),
    .A(_06554_),
    .B(_07088_));
 sg13g2_nand2_1 _17262_ (.Y(_07091_),
    .A(_07087_),
    .B(_07089_));
 sg13g2_nor2_1 _17263_ (.A(_07087_),
    .B(_07089_),
    .Y(_07092_));
 sg13g2_o21ai_1 _17264_ (.B1(_07091_),
    .Y(_07093_),
    .A1(_07085_),
    .A2(_07092_));
 sg13g2_a21o_1 _17265_ (.A2(_07092_),
    .A1(_07085_),
    .B1(_07093_),
    .X(_07094_));
 sg13g2_o21ai_1 _17266_ (.B1(_07094_),
    .Y(_07095_),
    .A1(_07085_),
    .A2(_07091_));
 sg13g2_xor2_1 _17267_ (.B(_06392_),
    .A(_06382_),
    .X(_07096_));
 sg13g2_xnor2_1 _17268_ (.Y(_07097_),
    .A(_06405_),
    .B(_07096_));
 sg13g2_nor2_1 _17269_ (.A(_06467_),
    .B(_06468_),
    .Y(_07098_));
 sg13g2_xor2_1 _17270_ (.B(_07098_),
    .A(_06480_),
    .X(_07099_));
 sg13g2_inv_1 _17271_ (.Y(_07100_),
    .A(_07099_));
 sg13g2_nand2_1 _17272_ (.Y(_07102_),
    .A(_07097_),
    .B(_07100_));
 sg13g2_nand2b_1 _17273_ (.Y(_07103_),
    .B(_07099_),
    .A_N(_07097_));
 sg13g2_nand2_1 _17274_ (.Y(_07104_),
    .A(_07102_),
    .B(_07103_));
 sg13g2_nor2_1 _17275_ (.A(_06428_),
    .B(_06429_),
    .Y(_07105_));
 sg13g2_xnor2_1 _17276_ (.Y(_07106_),
    .A(_06442_),
    .B(_07105_));
 sg13g2_xor2_1 _17277_ (.B(_07106_),
    .A(_07104_),
    .X(_07107_));
 sg13g2_nand2_1 _17278_ (.Y(_07108_),
    .A(_07095_),
    .B(_07107_));
 sg13g2_or2_1 _17279_ (.X(_07109_),
    .B(_07107_),
    .A(_07095_));
 sg13g2_nand2_1 _17280_ (.Y(_07110_),
    .A(_07108_),
    .B(_07109_));
 sg13g2_nor2_1 _17281_ (.A(_06974_),
    .B(_06975_),
    .Y(_07111_));
 sg13g2_xnor2_1 _17282_ (.Y(_07113_),
    .A(_06983_),
    .B(_07111_));
 sg13g2_xnor2_1 _17283_ (.Y(_07114_),
    .A(_07110_),
    .B(_07113_));
 sg13g2_nand2_1 _17284_ (.Y(_07115_),
    .A(_07083_),
    .B(_07114_));
 sg13g2_nor2_1 _17285_ (.A(_07083_),
    .B(_07114_),
    .Y(_07116_));
 sg13g2_xor2_1 _17286_ (.B(_07114_),
    .A(_07083_),
    .X(_07117_));
 sg13g2_or2_1 _17287_ (.X(_07118_),
    .B(_06959_),
    .A(_06950_));
 sg13g2_a22oi_1 _17288_ (.Y(_07119_),
    .B1(_06960_),
    .B2(_07118_),
    .A2(_06959_),
    .A1(_06951_));
 sg13g2_xnor2_1 _17289_ (.Y(_07120_),
    .A(_07117_),
    .B(_07119_));
 sg13g2_a21o_2 _17290_ (.A2(_06307_),
    .A1(_06302_),
    .B1(_06303_),
    .X(_07121_));
 sg13g2_inv_1 _17291_ (.Y(_07122_),
    .A(_07121_));
 sg13g2_o21ai_1 _17292_ (.B1(_07115_),
    .Y(_07124_),
    .A1(_07116_),
    .A2(_07119_));
 sg13g2_nor3_1 _17293_ (.A(_07115_),
    .B(_07119_),
    .C(_07121_),
    .Y(_07125_));
 sg13g2_a21oi_2 _17294_ (.B1(_07124_),
    .Y(_07126_),
    .A2(_07122_),
    .A1(_07120_));
 sg13g2_o21ai_1 _17295_ (.B1(_07069_),
    .Y(_07127_),
    .A1(_07070_),
    .A2(_07082_));
 sg13g2_o21ai_1 _17296_ (.B1(_07127_),
    .Y(_07128_),
    .A1(_07125_),
    .A2(_07126_));
 sg13g2_or3_1 _17297_ (.A(_07125_),
    .B(_07126_),
    .C(_07127_),
    .X(_07129_));
 sg13g2_a21o_1 _17298_ (.A2(_07048_),
    .A1(_07044_),
    .B1(_07052_),
    .X(_07130_));
 sg13g2_nand2_1 _17299_ (.Y(_07131_),
    .A(_07109_),
    .B(_07113_));
 sg13g2_a22oi_1 _17300_ (.Y(_07132_),
    .B1(_07131_),
    .B2(_07108_),
    .A2(_07130_),
    .A1(_07049_));
 sg13g2_nand4_1 _17301_ (.B(_07108_),
    .C(_07130_),
    .A(_07049_),
    .Y(_07133_),
    .D(_07131_));
 sg13g2_nor2b_1 _17302_ (.A(_07132_),
    .B_N(_07133_),
    .Y(_07135_));
 sg13g2_xnor2_1 _17303_ (.Y(_07136_),
    .A(_07065_),
    .B(_07135_));
 sg13g2_inv_1 _17304_ (.Y(_07137_),
    .A(_07136_));
 sg13g2_a21oi_1 _17305_ (.A1(_07128_),
    .A2(_07129_),
    .Y(_07138_),
    .B1(_07137_));
 sg13g2_and3_1 _17306_ (.X(_07139_),
    .A(_07128_),
    .B(_07129_),
    .C(_07137_));
 sg13g2_nand2_1 _17307_ (.Y(_07140_),
    .A(_07103_),
    .B(_07106_));
 sg13g2_and2_1 _17308_ (.A(_07102_),
    .B(_07140_),
    .X(_07141_));
 sg13g2_a21o_1 _17309_ (.A2(_07081_),
    .A1(_07076_),
    .B1(_07077_),
    .X(_07142_));
 sg13g2_xnor2_1 _17310_ (.Y(_07143_),
    .A(_07141_),
    .B(_07142_));
 sg13g2_xor2_1 _17311_ (.B(_07143_),
    .A(_07093_),
    .X(_07144_));
 sg13g2_or3_1 _17312_ (.A(_07138_),
    .B(_07139_),
    .C(_07144_),
    .X(_07146_));
 sg13g2_o21ai_1 _17313_ (.B1(_07144_),
    .Y(_07147_),
    .A1(_07138_),
    .A2(_07139_));
 sg13g2_nand2_1 _17314_ (.Y(_07148_),
    .A(_06986_),
    .B(_07009_));
 sg13g2_xor2_1 _17315_ (.B(_07148_),
    .A(_07008_),
    .X(_07149_));
 sg13g2_nand2_1 _17316_ (.Y(_07150_),
    .A(_06924_),
    .B(_06933_));
 sg13g2_xnor2_1 _17317_ (.Y(_07151_),
    .A(_06932_),
    .B(_07150_));
 sg13g2_xnor2_1 _17318_ (.Y(_07152_),
    .A(_07149_),
    .B(_07151_));
 sg13g2_nand2_1 _17319_ (.Y(_07153_),
    .A(_07030_),
    .B(_07032_));
 sg13g2_xor2_1 _17320_ (.B(_07153_),
    .A(_07041_),
    .X(_07154_));
 sg13g2_xnor2_1 _17321_ (.Y(_07155_),
    .A(_07152_),
    .B(_07154_));
 sg13g2_a21oi_1 _17322_ (.A1(_07146_),
    .A2(_07147_),
    .Y(_07157_),
    .B1(_07155_));
 sg13g2_nand3_1 _17323_ (.B(_07147_),
    .C(_07155_),
    .A(_07146_),
    .Y(_07158_));
 sg13g2_nor2_1 _17324_ (.A(_06588_),
    .B(_06623_),
    .Y(_07159_));
 sg13g2_a21oi_1 _17325_ (.A1(_06587_),
    .A2(_06623_),
    .Y(_07160_),
    .B1(_06624_));
 sg13g2_nor2_2 _17326_ (.A(_07159_),
    .B(_07160_),
    .Y(_07161_));
 sg13g2_nor2_1 _17327_ (.A(_06367_),
    .B(_06407_),
    .Y(_07162_));
 sg13g2_nor2_1 _17328_ (.A(_06409_),
    .B(_07162_),
    .Y(_07163_));
 sg13g2_a21oi_1 _17329_ (.A1(_06368_),
    .A2(_06407_),
    .Y(_07164_),
    .B1(_07163_));
 sg13g2_nor2_1 _17330_ (.A(_06483_),
    .B(_06484_),
    .Y(_07165_));
 sg13g2_xnor2_1 _17331_ (.Y(_07166_),
    .A(_06515_),
    .B(_07165_));
 sg13g2_nand2_1 _17332_ (.Y(_07168_),
    .A(_07164_),
    .B(_07166_));
 sg13g2_or2_1 _17333_ (.X(_07169_),
    .B(_07166_),
    .A(_07164_));
 sg13g2_nand2_1 _17334_ (.Y(_07170_),
    .A(_07161_),
    .B(_07169_));
 sg13g2_nand2_1 _17335_ (.Y(_07171_),
    .A(_07168_),
    .B(_07170_));
 sg13g2_nand2_1 _17336_ (.Y(_07172_),
    .A(_07168_),
    .B(_07169_));
 sg13g2_xnor2_1 _17337_ (.Y(_07173_),
    .A(_07161_),
    .B(_07172_));
 sg13g2_o21ai_1 _17338_ (.B1(_07158_),
    .Y(_07174_),
    .A1(_07157_),
    .A2(_07173_));
 sg13g2_a21o_1 _17339_ (.A2(_06946_),
    .A1(_06945_),
    .B1(_06778_),
    .X(_07175_));
 sg13g2_o21ai_1 _17340_ (.B1(_07175_),
    .Y(_07176_),
    .A1(_06945_),
    .A2(_06946_));
 sg13g2_nor2_1 _17341_ (.A(_06976_),
    .B(_06979_),
    .Y(_07177_));
 sg13g2_nor2_2 _17342_ (.A(_06981_),
    .B(_07177_),
    .Y(_07179_));
 sg13g2_nand2_1 _17343_ (.Y(_07180_),
    .A(_06971_),
    .B(_07179_));
 sg13g2_xor2_1 _17344_ (.B(_07179_),
    .A(_06971_),
    .X(_07181_));
 sg13g2_a21oi_1 _17345_ (.A1(_06937_),
    .A2(_06941_),
    .Y(_07182_),
    .B1(_06942_));
 sg13g2_xnor2_1 _17346_ (.Y(_07183_),
    .A(_07181_),
    .B(_07182_));
 sg13g2_nand2b_1 _17347_ (.Y(_07184_),
    .B(_07183_),
    .A_N(_07176_));
 sg13g2_inv_1 _17348_ (.Y(_07185_),
    .A(_07184_));
 sg13g2_nand2b_1 _17349_ (.Y(_07186_),
    .B(_07176_),
    .A_N(_07183_));
 sg13g2_a21oi_2 _17350_ (.B1(_07185_),
    .Y(_07187_),
    .A2(_07186_),
    .A1(_06957_));
 sg13g2_or2_1 _17351_ (.X(_07188_),
    .B(_07186_),
    .A(_06957_));
 sg13g2_a22oi_1 _17352_ (.Y(_07190_),
    .B1(_07187_),
    .B2(_07188_),
    .A2(_07185_),
    .A1(_06957_));
 sg13g2_inv_1 _17353_ (.Y(_07191_),
    .A(_07190_));
 sg13g2_and2_1 _17354_ (.A(_07157_),
    .B(_07173_),
    .X(_07192_));
 sg13g2_or2_1 _17355_ (.X(_07193_),
    .B(_07173_),
    .A(_07158_));
 sg13g2_o21ai_1 _17356_ (.B1(_07193_),
    .Y(_07194_),
    .A1(_07174_),
    .A2(_07192_));
 sg13g2_a21oi_1 _17357_ (.A1(_07191_),
    .A2(_07194_),
    .Y(_07195_),
    .B1(_07174_));
 sg13g2_nor2_1 _17358_ (.A(_07190_),
    .B(_07193_),
    .Y(_07196_));
 sg13g2_nor2_1 _17359_ (.A(_07139_),
    .B(_07144_),
    .Y(_07197_));
 sg13g2_or2_1 _17360_ (.X(_07198_),
    .B(_07197_),
    .A(_07138_));
 sg13g2_nor2_1 _17361_ (.A(_07196_),
    .B(_07198_),
    .Y(_07199_));
 sg13g2_or2_1 _17362_ (.X(_07201_),
    .B(_07199_),
    .A(_07195_));
 sg13g2_a21o_1 _17363_ (.A2(_07151_),
    .A1(_07149_),
    .B1(_07154_),
    .X(_07202_));
 sg13g2_o21ai_1 _17364_ (.B1(_07202_),
    .Y(_07203_),
    .A1(_07149_),
    .A2(_07151_));
 sg13g2_nand2_1 _17365_ (.Y(_07204_),
    .A(_07171_),
    .B(_07203_));
 sg13g2_or2_1 _17366_ (.X(_07205_),
    .B(_07203_),
    .A(_07171_));
 sg13g2_nand2_1 _17367_ (.Y(_07206_),
    .A(_07187_),
    .B(_07205_));
 sg13g2_nand2_1 _17368_ (.Y(_07207_),
    .A(_07204_),
    .B(_07206_));
 sg13g2_nand2_1 _17369_ (.Y(_07208_),
    .A(_07201_),
    .B(_07207_));
 sg13g2_nor2_1 _17370_ (.A(_07201_),
    .B(_07207_),
    .Y(_07209_));
 sg13g2_inv_1 _17371_ (.Y(_07210_),
    .A(_07209_));
 sg13g2_nand2_1 _17372_ (.Y(_07212_),
    .A(_07208_),
    .B(_07210_));
 sg13g2_nor2_1 _17373_ (.A(_07125_),
    .B(_07127_),
    .Y(_07213_));
 sg13g2_nor2_1 _17374_ (.A(_07126_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_a21oi_2 _17375_ (.B1(_07132_),
    .Y(_07215_),
    .A2(_07133_),
    .A1(_07066_));
 sg13g2_or3_1 _17376_ (.A(_07126_),
    .B(_07213_),
    .C(_07215_),
    .X(_07216_));
 sg13g2_nor2b_1 _17377_ (.A(_07214_),
    .B_N(_07215_),
    .Y(_07217_));
 sg13g2_a21o_1 _17378_ (.A2(_07142_),
    .A1(_07141_),
    .B1(_07093_),
    .X(_07218_));
 sg13g2_o21ai_1 _17379_ (.B1(_07218_),
    .Y(_07219_),
    .A1(_07141_),
    .A2(_07142_));
 sg13g2_a21oi_2 _17380_ (.B1(_07217_),
    .Y(_07220_),
    .A2(_07219_),
    .A1(_07216_));
 sg13g2_xnor2_1 _17381_ (.Y(_07221_),
    .A(_07212_),
    .B(_07220_));
 sg13g2_or2_1 _17382_ (.X(_07223_),
    .B(_06624_),
    .A(_06517_));
 sg13g2_a22oi_1 _17383_ (.Y(_07224_),
    .B1(_06625_),
    .B2(_07223_),
    .A2(_06624_),
    .A1(_06520_));
 sg13g2_xor2_1 _17384_ (.B(_07011_),
    .A(_06935_),
    .X(_07225_));
 sg13g2_xnor2_1 _17385_ (.Y(_07226_),
    .A(_07042_),
    .B(_07225_));
 sg13g2_xor2_1 _17386_ (.B(_07226_),
    .A(_07224_),
    .X(_07227_));
 sg13g2_nand2_1 _17387_ (.Y(_07228_),
    .A(_07180_),
    .B(_07182_));
 sg13g2_o21ai_1 _17388_ (.B1(_07228_),
    .Y(_07229_),
    .A1(_06971_),
    .A2(_07179_));
 sg13g2_xnor2_1 _17389_ (.Y(_07230_),
    .A(_07227_),
    .B(_07229_));
 sg13g2_nand2_1 _17390_ (.Y(_07231_),
    .A(_07204_),
    .B(_07205_));
 sg13g2_xor2_1 _17391_ (.B(_07231_),
    .A(_07187_),
    .X(_07232_));
 sg13g2_inv_1 _17392_ (.Y(_07234_),
    .A(_07232_));
 sg13g2_or3_1 _17393_ (.A(_07195_),
    .B(_07196_),
    .C(_07198_),
    .X(_07235_));
 sg13g2_o21ai_1 _17394_ (.B1(_07198_),
    .Y(_07236_),
    .A1(_07195_),
    .A2(_07196_));
 sg13g2_a21oi_1 _17395_ (.A1(_07235_),
    .A2(_07236_),
    .Y(_07237_),
    .B1(_07234_));
 sg13g2_a21o_1 _17396_ (.A2(_07236_),
    .A1(_07235_),
    .B1(_07234_),
    .X(_07238_));
 sg13g2_nand3_1 _17397_ (.B(_07235_),
    .C(_07236_),
    .A(_07234_),
    .Y(_07239_));
 sg13g2_xnor2_1 _17398_ (.Y(_07240_),
    .A(_07214_),
    .B(_07215_));
 sg13g2_xnor2_1 _17399_ (.Y(_07241_),
    .A(_07219_),
    .B(_07240_));
 sg13g2_a21o_1 _17400_ (.A2(_07239_),
    .A1(_07238_),
    .B1(_07241_),
    .X(_07242_));
 sg13g2_nand3_1 _17401_ (.B(_07239_),
    .C(_07241_),
    .A(_07238_),
    .Y(_07243_));
 sg13g2_and3_1 _17402_ (.X(_07245_),
    .A(_07230_),
    .B(_07242_),
    .C(_07243_));
 sg13g2_o21ai_1 _17403_ (.B1(_07239_),
    .Y(_07246_),
    .A1(_07237_),
    .A2(_07241_));
 sg13g2_nand2b_1 _17404_ (.Y(_07247_),
    .B(_07246_),
    .A_N(_07245_));
 sg13g2_nor2b_1 _17405_ (.A(_07246_),
    .B_N(_07245_),
    .Y(_07248_));
 sg13g2_xor2_1 _17406_ (.B(_07246_),
    .A(_07245_),
    .X(_07249_));
 sg13g2_a21o_1 _17407_ (.A2(_07226_),
    .A1(_07224_),
    .B1(_07229_),
    .X(_07250_));
 sg13g2_o21ai_1 _17408_ (.B1(_07250_),
    .Y(_07251_),
    .A1(_07224_),
    .A2(_07226_));
 sg13g2_xnor2_1 _17409_ (.Y(_07252_),
    .A(_07249_),
    .B(_07251_));
 sg13g2_nand2_1 _17410_ (.Y(_07253_),
    .A(_07221_),
    .B(_07252_));
 sg13g2_nor2_1 _17411_ (.A(_07221_),
    .B(_07252_),
    .Y(_07254_));
 sg13g2_xor2_1 _17412_ (.B(_07252_),
    .A(_07221_),
    .X(_07256_));
 sg13g2_xnor2_1 _17413_ (.Y(_07257_),
    .A(_07043_),
    .B(_07256_));
 sg13g2_o21ai_1 _17414_ (.B1(_07253_),
    .Y(_07258_),
    .A1(_07043_),
    .A2(_07254_));
 sg13g2_nor3_1 _17415_ (.A(_06625_),
    .B(_07043_),
    .C(_07253_),
    .Y(_07259_));
 sg13g2_inv_1 _17416_ (.Y(_07260_),
    .A(_07259_));
 sg13g2_a21o_1 _17417_ (.A2(_07257_),
    .A1(_06626_),
    .B1(_07258_),
    .X(_07261_));
 sg13g2_a21o_1 _17418_ (.A2(_07251_),
    .A1(_07247_),
    .B1(_07248_),
    .X(_07262_));
 sg13g2_inv_1 _17419_ (.Y(_07263_),
    .A(_07262_));
 sg13g2_a21oi_1 _17420_ (.A1(_07260_),
    .A2(_07261_),
    .Y(_07264_),
    .B1(_07263_));
 sg13g2_and3_1 _17421_ (.X(_07265_),
    .A(_07260_),
    .B(_07261_),
    .C(_07263_));
 sg13g2_a21oi_1 _17422_ (.A1(_07208_),
    .A2(_07220_),
    .Y(_07267_),
    .B1(_07209_));
 sg13g2_inv_1 _17423_ (.Y(_07268_),
    .A(_07267_));
 sg13g2_o21ai_1 _17424_ (.B1(_07268_),
    .Y(_07269_),
    .A1(_07264_),
    .A2(_07265_));
 sg13g2_o21ai_1 _17425_ (.B1(_07261_),
    .Y(_07270_),
    .A1(_07259_),
    .A2(_07262_));
 sg13g2_and2_1 _17426_ (.A(_07269_),
    .B(_07270_),
    .X(_07271_));
 sg13g2_nand2_2 _17427_ (.Y(_07272_),
    .A(_07269_),
    .B(_07270_));
 sg13g2_nand2b_1 _17428_ (.Y(_07273_),
    .B(_05846_),
    .A_N(_05842_));
 sg13g2_o21ai_1 _17429_ (.B1(_05826_),
    .Y(_07274_),
    .A1(_05828_),
    .A2(_05831_));
 sg13g2_a22oi_1 _17430_ (.Y(_07275_),
    .B1(_07274_),
    .B2(_05832_),
    .A2(_07273_),
    .A1(_05845_));
 sg13g2_nand4_1 _17431_ (.B(_05845_),
    .C(_07273_),
    .A(_05832_),
    .Y(_07276_),
    .D(_07274_));
 sg13g2_nand2b_1 _17432_ (.Y(_07278_),
    .B(_07276_),
    .A_N(_07275_));
 sg13g2_a21oi_2 _17433_ (.B1(_07275_),
    .Y(_07279_),
    .A2(_07276_),
    .A1(_05823_));
 sg13g2_xnor2_1 _17434_ (.Y(_07280_),
    .A(_05823_),
    .B(_07278_));
 sg13g2_a21o_2 _17435_ (.A2(_05764_),
    .A1(_05760_),
    .B1(_05763_),
    .X(_07281_));
 sg13g2_o21ai_1 _17436_ (.B1(_05808_),
    .Y(_07282_),
    .A1(_05802_),
    .A2(_05809_));
 sg13g2_nor2b_1 _17437_ (.A(_07281_),
    .B_N(_07282_),
    .Y(_07283_));
 sg13g2_nand2b_1 _17438_ (.Y(_07284_),
    .B(_07281_),
    .A_N(_07282_));
 sg13g2_nor2b_1 _17439_ (.A(_07283_),
    .B_N(_07284_),
    .Y(_07285_));
 sg13g2_a21oi_2 _17440_ (.B1(_07283_),
    .Y(_07286_),
    .A2(_07284_),
    .A1(_05779_));
 sg13g2_xnor2_1 _17441_ (.Y(_07287_),
    .A(_05778_),
    .B(_07285_));
 sg13g2_nor2_1 _17442_ (.A(_07280_),
    .B(_07287_),
    .Y(_07289_));
 sg13g2_nand2_1 _17443_ (.Y(_07290_),
    .A(_07280_),
    .B(_07287_));
 sg13g2_a21oi_1 _17444_ (.A1(_05727_),
    .A2(_05730_),
    .Y(_07291_),
    .B1(_05729_));
 sg13g2_a21oi_1 _17445_ (.A1(_05736_),
    .A2(_05738_),
    .Y(_07292_),
    .B1(_05733_));
 sg13g2_nor2_1 _17446_ (.A(_05739_),
    .B(_07292_),
    .Y(_07293_));
 sg13g2_nor2b_1 _17447_ (.A(_05786_),
    .B_N(_05790_),
    .Y(_07294_));
 sg13g2_nor2_2 _17448_ (.A(_05791_),
    .B(_07294_),
    .Y(_07295_));
 sg13g2_and2_1 _17449_ (.A(_07293_),
    .B(_07295_),
    .X(_07296_));
 sg13g2_xor2_1 _17450_ (.B(_07295_),
    .A(_07293_),
    .X(_07297_));
 sg13g2_xnor2_1 _17451_ (.Y(_07298_),
    .A(_07291_),
    .B(_07297_));
 sg13g2_o21ai_1 _17452_ (.B1(_07290_),
    .Y(_07300_),
    .A1(_07289_),
    .A2(_07298_));
 sg13g2_o21ai_1 _17453_ (.B1(_06244_),
    .Y(_07301_),
    .A1(_06242_),
    .A2(_06246_));
 sg13g2_o21ai_1 _17454_ (.B1(_06183_),
    .Y(_07302_),
    .A1(_06176_),
    .A2(_06182_));
 sg13g2_nand2b_1 _17455_ (.Y(_07303_),
    .B(_07301_),
    .A_N(_07302_));
 sg13g2_nor2b_1 _17456_ (.A(_07301_),
    .B_N(_07302_),
    .Y(_07304_));
 sg13g2_xnor2_1 _17457_ (.Y(_07305_),
    .A(_07301_),
    .B(_07302_));
 sg13g2_a21o_1 _17458_ (.A2(_06236_),
    .A1(_06231_),
    .B1(_06233_),
    .X(_07306_));
 sg13g2_xnor2_1 _17459_ (.Y(_07307_),
    .A(_07305_),
    .B(_07306_));
 sg13g2_o21ai_1 _17460_ (.B1(_05905_),
    .Y(_07308_),
    .A1(_05899_),
    .A2(_05906_));
 sg13g2_a21oi_1 _17461_ (.A1(_05892_),
    .A2(_05895_),
    .Y(_07309_),
    .B1(_05890_));
 sg13g2_o21ai_1 _17462_ (.B1(_06260_),
    .Y(_07311_),
    .A1(_05896_),
    .A2(_07309_));
 sg13g2_nor3_1 _17463_ (.A(_05896_),
    .B(_06260_),
    .C(_07309_),
    .Y(_07312_));
 sg13g2_inv_1 _17464_ (.Y(_07313_),
    .A(_07312_));
 sg13g2_nand2_1 _17465_ (.Y(_07314_),
    .A(_07311_),
    .B(_07313_));
 sg13g2_xnor2_1 _17466_ (.Y(_07315_),
    .A(_07308_),
    .B(_07314_));
 sg13g2_inv_1 _17467_ (.Y(_07316_),
    .A(_07315_));
 sg13g2_nand2_1 _17468_ (.Y(_07317_),
    .A(_07307_),
    .B(_07316_));
 sg13g2_nand2b_1 _17469_ (.Y(_07318_),
    .B(_07315_),
    .A_N(_07307_));
 sg13g2_o21ai_1 _17470_ (.B1(_05862_),
    .Y(_07319_),
    .A1(_05863_),
    .A2(_05864_));
 sg13g2_nand2_2 _17471_ (.Y(_07320_),
    .A(_05865_),
    .B(_07319_));
 sg13g2_o21ai_1 _17472_ (.B1(_05884_),
    .Y(_07322_),
    .A1(_05875_),
    .A2(_05885_));
 sg13g2_a21oi_2 _17473_ (.B1(_05857_),
    .Y(_07323_),
    .A2(_05859_),
    .A1(_05850_));
 sg13g2_nor2_1 _17474_ (.A(_07322_),
    .B(_07323_),
    .Y(_07324_));
 sg13g2_nand2_1 _17475_ (.Y(_07325_),
    .A(_07322_),
    .B(_07323_));
 sg13g2_nor2b_1 _17476_ (.A(_07324_),
    .B_N(_07325_),
    .Y(_07326_));
 sg13g2_xnor2_1 _17477_ (.Y(_07327_),
    .A(_07320_),
    .B(_07326_));
 sg13g2_nand2_1 _17478_ (.Y(_07328_),
    .A(_07318_),
    .B(_07327_));
 sg13g2_a21oi_1 _17479_ (.A1(_07317_),
    .A2(_07328_),
    .Y(_07329_),
    .B1(_07300_));
 sg13g2_a21oi_2 _17480_ (.B1(_05919_),
    .Y(_07330_),
    .A2(_06268_),
    .A1(_05920_));
 sg13g2_o21ai_1 _17481_ (.B1(_06151_),
    .Y(_07331_),
    .A1(_06150_),
    .A2(_06267_));
 sg13g2_nor2b_1 _17482_ (.A(_07330_),
    .B_N(_07331_),
    .Y(_07333_));
 sg13g2_and3_1 _17483_ (.X(_07334_),
    .A(_07300_),
    .B(_07317_),
    .C(_07328_));
 sg13g2_nor2_1 _17484_ (.A(_07333_),
    .B(_07334_),
    .Y(_07335_));
 sg13g2_nor2_1 _17485_ (.A(_07329_),
    .B(_07335_),
    .Y(_07336_));
 sg13g2_or2_1 _17486_ (.X(_07337_),
    .B(_06146_),
    .A(_06069_));
 sg13g2_nand2_1 _17487_ (.Y(_07338_),
    .A(_05956_),
    .B(_06031_));
 sg13g2_a22oi_1 _17488_ (.Y(_07339_),
    .B1(_07338_),
    .B2(_06032_),
    .A2(_07337_),
    .A1(_06147_));
 sg13g2_and4_1 _17489_ (.A(_06032_),
    .B(_06147_),
    .C(_07337_),
    .D(_07338_),
    .X(_07340_));
 sg13g2_nand2_1 _17490_ (.Y(_07341_),
    .A(_06226_),
    .B(_06264_));
 sg13g2_nor2_1 _17491_ (.A(_07340_),
    .B(_07341_),
    .Y(_07342_));
 sg13g2_o21ai_1 _17492_ (.B1(_05723_),
    .Y(_07344_),
    .A1(_05756_),
    .A2(_05796_));
 sg13g2_nand2_1 _17493_ (.Y(_07345_),
    .A(_05839_),
    .B(_05916_));
 sg13g2_and4_1 _17494_ (.A(_05797_),
    .B(_05915_),
    .C(_07344_),
    .D(_07345_),
    .X(_07346_));
 sg13g2_inv_1 _17495_ (.Y(_07347_),
    .A(_07346_));
 sg13g2_a22oi_1 _17496_ (.Y(_07348_),
    .B1(_07345_),
    .B2(_05915_),
    .A2(_07344_),
    .A1(_05797_));
 sg13g2_a21oi_2 _17497_ (.B1(_07348_),
    .Y(_07349_),
    .A2(_07347_),
    .A1(_05989_));
 sg13g2_o21ai_1 _17498_ (.B1(_07349_),
    .Y(_07350_),
    .A1(_07339_),
    .A2(_07342_));
 sg13g2_o21ai_1 _17499_ (.B1(_06003_),
    .Y(_07351_),
    .A1(_06017_),
    .A2(_06027_));
 sg13g2_and3_1 _17500_ (.X(_07352_),
    .A(_05954_),
    .B(_06028_),
    .C(_07351_));
 sg13g2_a21oi_1 _17501_ (.A1(_06028_),
    .A2(_07351_),
    .Y(_07353_),
    .B1(_05954_));
 sg13g2_o21ai_1 _17502_ (.B1(_06103_),
    .Y(_07355_),
    .A1(_06080_),
    .A2(_06104_));
 sg13g2_nor2_1 _17503_ (.A(_07353_),
    .B(_07355_),
    .Y(_07356_));
 sg13g2_nor2_1 _17504_ (.A(_07352_),
    .B(_07356_),
    .Y(_07357_));
 sg13g2_or3_1 _17505_ (.A(_07339_),
    .B(_07342_),
    .C(_07349_),
    .X(_07358_));
 sg13g2_nand2b_1 _17506_ (.Y(_07359_),
    .B(_07358_),
    .A_N(_07357_));
 sg13g2_a21oi_1 _17507_ (.A1(_07350_),
    .A2(_07359_),
    .Y(_07360_),
    .B1(_07336_));
 sg13g2_inv_1 _17508_ (.Y(_07361_),
    .A(_07360_));
 sg13g2_a21oi_1 _17509_ (.A1(_06116_),
    .A2(_06127_),
    .Y(_07362_),
    .B1(_06143_));
 sg13g2_nor2_1 _17510_ (.A(_06128_),
    .B(_07362_),
    .Y(_07363_));
 sg13g2_nand2_1 _17511_ (.Y(_07364_),
    .A(_06054_),
    .B(_06068_));
 sg13g2_nand3_1 _17512_ (.B(_07363_),
    .C(_07364_),
    .A(_06053_),
    .Y(_07366_));
 sg13g2_a21o_1 _17513_ (.A2(_07364_),
    .A1(_06053_),
    .B1(_07363_),
    .X(_07367_));
 sg13g2_nand2_1 _17514_ (.Y(_07368_),
    .A(_06224_),
    .B(_07367_));
 sg13g2_nand2_1 _17515_ (.Y(_07369_),
    .A(_07366_),
    .B(_07368_));
 sg13g2_inv_1 _17516_ (.Y(_07370_),
    .A(_07369_));
 sg13g2_o21ai_1 _17517_ (.B1(_06172_),
    .Y(_07371_),
    .A1(_06173_),
    .A2(_06185_));
 sg13g2_nand2_1 _17518_ (.Y(_07372_),
    .A(_06249_),
    .B(_06262_));
 sg13g2_and3_1 _17519_ (.X(_07373_),
    .A(_06248_),
    .B(_07371_),
    .C(_07372_));
 sg13g2_a21oi_1 _17520_ (.A1(_06248_),
    .A2(_07372_),
    .Y(_07374_),
    .B1(_07371_));
 sg13g2_nor2_1 _17521_ (.A(_05911_),
    .B(_07374_),
    .Y(_07375_));
 sg13g2_nor2_1 _17522_ (.A(_07373_),
    .B(_07375_),
    .Y(_07377_));
 sg13g2_nor2_1 _17523_ (.A(_07370_),
    .B(_07377_),
    .Y(_07378_));
 sg13g2_a21oi_2 _17524_ (.B1(_05835_),
    .Y(_07379_),
    .A2(_05837_),
    .A1(_05811_));
 sg13g2_nand2_1 _17525_ (.Y(_07380_),
    .A(_05872_),
    .B(_07379_));
 sg13g2_nor2_1 _17526_ (.A(_05872_),
    .B(_07379_),
    .Y(_07381_));
 sg13g2_o21ai_1 _17527_ (.B1(_05783_),
    .Y(_07382_),
    .A1(_05784_),
    .A2(_05794_));
 sg13g2_a21oi_2 _17528_ (.B1(_07381_),
    .Y(_07383_),
    .A2(_07382_),
    .A1(_07380_));
 sg13g2_nand2_1 _17529_ (.Y(_07384_),
    .A(_07370_),
    .B(_07377_));
 sg13g2_o21ai_1 _17530_ (.B1(_07384_),
    .Y(_07385_),
    .A1(_07378_),
    .A2(_07383_));
 sg13g2_and3_1 _17531_ (.X(_07386_),
    .A(_07336_),
    .B(_07350_),
    .C(_07359_));
 sg13g2_a21oi_2 _17532_ (.B1(_07386_),
    .Y(_07388_),
    .A2(_07385_),
    .A1(_07361_));
 sg13g2_inv_1 _17533_ (.Y(_07389_),
    .A(_07388_));
 sg13g2_o21ai_1 _17534_ (.B1(_07311_),
    .Y(_07390_),
    .A1(_07308_),
    .A2(_07312_));
 sg13g2_a21oi_2 _17535_ (.B1(_07324_),
    .Y(_07391_),
    .A2(_07325_),
    .A1(_07320_));
 sg13g2_a21o_1 _17536_ (.A2(_07391_),
    .A1(_07390_),
    .B1(_07279_),
    .X(_07392_));
 sg13g2_o21ai_1 _17537_ (.B1(_07392_),
    .Y(_07393_),
    .A1(_07390_),
    .A2(_07391_));
 sg13g2_xnor2_1 _17538_ (.Y(_07394_),
    .A(_07390_),
    .B(_07391_));
 sg13g2_xnor2_1 _17539_ (.Y(_07395_),
    .A(_07279_),
    .B(_07394_));
 sg13g2_nand2_1 _17540_ (.Y(_07396_),
    .A(_07286_),
    .B(_07395_));
 sg13g2_xor2_1 _17541_ (.B(_07395_),
    .A(_07286_),
    .X(_07397_));
 sg13g2_o21ai_1 _17542_ (.B1(_07291_),
    .Y(_07399_),
    .A1(_07293_),
    .A2(_07295_));
 sg13g2_nor2b_2 _17543_ (.A(_07296_),
    .B_N(_07399_),
    .Y(_07400_));
 sg13g2_xnor2_1 _17544_ (.Y(_07401_),
    .A(_07397_),
    .B(_07400_));
 sg13g2_nand2_1 _17545_ (.Y(_07402_),
    .A(_07350_),
    .B(_07358_));
 sg13g2_xor2_1 _17546_ (.B(_07402_),
    .A(_07357_),
    .X(_07403_));
 sg13g2_nor2_1 _17547_ (.A(_07329_),
    .B(_07334_),
    .Y(_07404_));
 sg13g2_xnor2_1 _17548_ (.Y(_07405_),
    .A(_07333_),
    .B(_07404_));
 sg13g2_nor2_1 _17549_ (.A(_07403_),
    .B(_07405_),
    .Y(_07406_));
 sg13g2_nand2_1 _17550_ (.Y(_07407_),
    .A(_07403_),
    .B(_07405_));
 sg13g2_nand2b_1 _17551_ (.Y(_07408_),
    .B(_07407_),
    .A_N(_07406_));
 sg13g2_nor2b_1 _17552_ (.A(_07378_),
    .B_N(_07384_),
    .Y(_07410_));
 sg13g2_xnor2_1 _17553_ (.Y(_07411_),
    .A(_07383_),
    .B(_07410_));
 sg13g2_xnor2_1 _17554_ (.Y(_07412_),
    .A(_07408_),
    .B(_07411_));
 sg13g2_and2_1 _17555_ (.A(_07317_),
    .B(_07318_),
    .X(_07413_));
 sg13g2_xnor2_1 _17556_ (.Y(_07414_),
    .A(_07327_),
    .B(_07413_));
 sg13g2_o21ai_1 _17557_ (.B1(_05944_),
    .Y(_07415_),
    .A1(_05945_),
    .A2(_05949_));
 sg13g2_nand2_1 _17558_ (.Y(_07416_),
    .A(_05950_),
    .B(_07415_));
 sg13g2_a21oi_2 _17559_ (.B1(_06095_),
    .Y(_07417_),
    .A2(_06101_),
    .A1(_06094_));
 sg13g2_and2_1 _17560_ (.A(_07416_),
    .B(_07417_),
    .X(_07418_));
 sg13g2_nor2_1 _17561_ (.A(_07416_),
    .B(_07417_),
    .Y(_07419_));
 sg13g2_nor2_1 _17562_ (.A(_07418_),
    .B(_07419_),
    .Y(_07421_));
 sg13g2_nor2b_1 _17563_ (.A(_07418_),
    .B_N(_06090_),
    .Y(_07422_));
 sg13g2_xnor2_1 _17564_ (.Y(_07423_),
    .A(_06090_),
    .B(_07421_));
 sg13g2_o21ai_1 _17565_ (.B1(_05930_),
    .Y(_07424_),
    .A1(_05923_),
    .A2(_05931_));
 sg13g2_o21ai_1 _17566_ (.B1(_05997_),
    .Y(_07425_),
    .A1(_05996_),
    .A2(_06002_));
 sg13g2_nor2_1 _17567_ (.A(_07424_),
    .B(_07425_),
    .Y(_07426_));
 sg13g2_nand2_1 _17568_ (.Y(_07427_),
    .A(_07424_),
    .B(_07425_));
 sg13g2_nand2b_1 _17569_ (.Y(_07428_),
    .B(_07427_),
    .A_N(_07426_));
 sg13g2_a21oi_1 _17570_ (.A1(_05938_),
    .A2(_05941_),
    .Y(_07429_),
    .B1(_05937_));
 sg13g2_xnor2_1 _17571_ (.Y(_07430_),
    .A(_07428_),
    .B(_07429_));
 sg13g2_and2_1 _17572_ (.A(_07423_),
    .B(_07430_),
    .X(_07432_));
 sg13g2_nor2_1 _17573_ (.A(_07423_),
    .B(_07430_),
    .Y(_07433_));
 sg13g2_nor2_1 _17574_ (.A(_07432_),
    .B(_07433_),
    .Y(_07434_));
 sg13g2_nand2_1 _17575_ (.Y(_07435_),
    .A(_06123_),
    .B(_06126_));
 sg13g2_o21ai_1 _17576_ (.B1(_06075_),
    .Y(_07436_),
    .A1(_06074_),
    .A2(_06079_));
 sg13g2_nand3_1 _17577_ (.B(_07435_),
    .C(_07436_),
    .A(_06124_),
    .Y(_07437_));
 sg13g2_a21oi_1 _17578_ (.A1(_06124_),
    .A2(_07435_),
    .Y(_07438_),
    .B1(_07436_));
 sg13g2_inv_1 _17579_ (.Y(_07439_),
    .A(_07438_));
 sg13g2_nand2_1 _17580_ (.Y(_07440_),
    .A(_07437_),
    .B(_07439_));
 sg13g2_a21oi_2 _17581_ (.B1(_06114_),
    .Y(_07441_),
    .A2(_06113_),
    .A1(_06108_));
 sg13g2_xnor2_1 _17582_ (.Y(_07443_),
    .A(_07440_),
    .B(_07441_));
 sg13g2_xor2_1 _17583_ (.B(_07443_),
    .A(_07434_),
    .X(_07444_));
 sg13g2_a21o_1 _17584_ (.A2(_06156_),
    .A1(_06154_),
    .B1(_06153_),
    .X(_07445_));
 sg13g2_o21ai_1 _17585_ (.B1(_07445_),
    .Y(_07446_),
    .A1(_06154_),
    .A2(_06156_));
 sg13g2_a21o_1 _17586_ (.A2(_06193_),
    .A1(_06189_),
    .B1(_06194_),
    .X(_07447_));
 sg13g2_xnor2_1 _17587_ (.Y(_07448_),
    .A(_06170_),
    .B(_07447_));
 sg13g2_xnor2_1 _17588_ (.Y(_07449_),
    .A(_07446_),
    .B(_07448_));
 sg13g2_nor2_1 _17589_ (.A(_06132_),
    .B(_06140_),
    .Y(_07450_));
 sg13g2_a21oi_1 _17590_ (.A1(_06036_),
    .A2(_06039_),
    .Y(_07451_),
    .B1(_06040_));
 sg13g2_o21ai_1 _17591_ (.B1(_07451_),
    .Y(_07452_),
    .A1(_06141_),
    .A2(_07450_));
 sg13g2_or3_1 _17592_ (.A(_06141_),
    .B(_07450_),
    .C(_07451_),
    .X(_07454_));
 sg13g2_nand2_1 _17593_ (.Y(_07455_),
    .A(_07452_),
    .B(_07454_));
 sg13g2_a21o_1 _17594_ (.A2(_06049_),
    .A1(_06047_),
    .B1(_06044_),
    .X(_07456_));
 sg13g2_o21ai_1 _17595_ (.B1(_07456_),
    .Y(_07457_),
    .A1(_06047_),
    .A2(_06049_));
 sg13g2_xnor2_1 _17596_ (.Y(_07458_),
    .A(_07455_),
    .B(_07457_));
 sg13g2_a21o_1 _17597_ (.A2(_06063_),
    .A1(_06059_),
    .B1(_06066_),
    .X(_07459_));
 sg13g2_a21o_1 _17598_ (.A2(_07459_),
    .A1(_06064_),
    .B1(_06205_),
    .X(_07460_));
 sg13g2_nand3_1 _17599_ (.B(_06205_),
    .C(_07459_),
    .A(_06064_),
    .Y(_07461_));
 sg13g2_nand2_1 _17600_ (.Y(_07462_),
    .A(_07460_),
    .B(_07461_));
 sg13g2_a21oi_1 _17601_ (.A1(_06209_),
    .A2(_06216_),
    .Y(_07463_),
    .B1(_06217_));
 sg13g2_xnor2_1 _17602_ (.Y(_07465_),
    .A(_07462_),
    .B(_07463_));
 sg13g2_nand2_1 _17603_ (.Y(_07466_),
    .A(_07458_),
    .B(_07465_));
 sg13g2_nor2_1 _17604_ (.A(_07458_),
    .B(_07465_),
    .Y(_07467_));
 sg13g2_xnor2_1 _17605_ (.Y(_07468_),
    .A(_07458_),
    .B(_07465_));
 sg13g2_xnor2_1 _17606_ (.Y(_07469_),
    .A(_07449_),
    .B(_07468_));
 sg13g2_nand2b_1 _17607_ (.Y(_07470_),
    .B(_07469_),
    .A_N(_07444_));
 sg13g2_nand2b_1 _17608_ (.Y(_07471_),
    .B(_07444_),
    .A_N(_07469_));
 sg13g2_and2_1 _17609_ (.A(_07470_),
    .B(_07471_),
    .X(_07472_));
 sg13g2_xnor2_1 _17610_ (.Y(_07473_),
    .A(_07414_),
    .B(_07472_));
 sg13g2_xnor2_1 _17611_ (.Y(_07474_),
    .A(_07330_),
    .B(_07331_));
 sg13g2_nor2_1 _17612_ (.A(_07339_),
    .B(_07340_),
    .Y(_07476_));
 sg13g2_xnor2_1 _17613_ (.Y(_07477_),
    .A(_07341_),
    .B(_07476_));
 sg13g2_nor2b_1 _17614_ (.A(_07477_),
    .B_N(_07474_),
    .Y(_07478_));
 sg13g2_nand2b_1 _17615_ (.Y(_07479_),
    .B(_07477_),
    .A_N(_07474_));
 sg13g2_xor2_1 _17616_ (.B(_07477_),
    .A(_07474_),
    .X(_07480_));
 sg13g2_nor2_1 _17617_ (.A(_07346_),
    .B(_07348_),
    .Y(_07481_));
 sg13g2_xor2_1 _17618_ (.B(_07481_),
    .A(_05989_),
    .X(_07482_));
 sg13g2_xnor2_1 _17619_ (.Y(_07483_),
    .A(_07480_),
    .B(_07482_));
 sg13g2_nor2_1 _17620_ (.A(_07352_),
    .B(_07353_),
    .Y(_07484_));
 sg13g2_xor2_1 _17621_ (.B(_07484_),
    .A(_07355_),
    .X(_07485_));
 sg13g2_nand2_1 _17622_ (.Y(_07487_),
    .A(_07366_),
    .B(_07367_));
 sg13g2_xor2_1 _17623_ (.B(_07487_),
    .A(_06224_),
    .X(_07488_));
 sg13g2_nand2_1 _17624_ (.Y(_07489_),
    .A(_07485_),
    .B(_07488_));
 sg13g2_xnor2_1 _17625_ (.Y(_07490_),
    .A(_07485_),
    .B(_07488_));
 sg13g2_nor2_1 _17626_ (.A(_07373_),
    .B(_07374_),
    .Y(_07491_));
 sg13g2_xnor2_1 _17627_ (.Y(_07492_),
    .A(_05911_),
    .B(_07491_));
 sg13g2_xnor2_1 _17628_ (.Y(_07493_),
    .A(_07490_),
    .B(_07492_));
 sg13g2_inv_1 _17629_ (.Y(_07494_),
    .A(_07493_));
 sg13g2_nor2_1 _17630_ (.A(_07483_),
    .B(_07494_),
    .Y(_07495_));
 sg13g2_xnor2_1 _17631_ (.Y(_07496_),
    .A(_07483_),
    .B(_07494_));
 sg13g2_nand2_1 _17632_ (.Y(_07498_),
    .A(_05959_),
    .B(_05964_));
 sg13g2_a21oi_1 _17633_ (.A1(_05965_),
    .A2(_07498_),
    .Y(_07499_),
    .B1(_06016_));
 sg13g2_nand3_1 _17634_ (.B(_06016_),
    .C(_07498_),
    .A(_05965_),
    .Y(_07500_));
 sg13g2_nand2b_1 _17635_ (.Y(_07501_),
    .B(_07500_),
    .A_N(_07499_));
 sg13g2_o21ai_1 _17636_ (.B1(_06025_),
    .Y(_07502_),
    .A1(_06019_),
    .A2(_06020_));
 sg13g2_nand2_1 _17637_ (.Y(_07503_),
    .A(_06021_),
    .B(_07502_));
 sg13g2_and2_1 _17638_ (.A(_07500_),
    .B(_07503_),
    .X(_07504_));
 sg13g2_xnor2_1 _17639_ (.Y(_07505_),
    .A(_07501_),
    .B(_07503_));
 sg13g2_xor2_1 _17640_ (.B(_07379_),
    .A(_05872_),
    .X(_07506_));
 sg13g2_xnor2_1 _17641_ (.Y(_07507_),
    .A(_07382_),
    .B(_07506_));
 sg13g2_o21ai_1 _17642_ (.B1(_05983_),
    .Y(_07509_),
    .A1(_05976_),
    .A2(_05981_));
 sg13g2_o21ai_1 _17643_ (.B1(_05973_),
    .Y(_07510_),
    .A1(_04750_),
    .A2(_05970_));
 sg13g2_nand2_2 _17644_ (.Y(_07511_),
    .A(_05971_),
    .B(_07510_));
 sg13g2_o21ai_1 _17645_ (.B1(_05755_),
    .Y(_07512_),
    .A1(_05732_),
    .A2(_05741_));
 sg13g2_nand2_1 _17646_ (.Y(_07513_),
    .A(_05742_),
    .B(_07512_));
 sg13g2_nor2_1 _17647_ (.A(_07511_),
    .B(_07513_),
    .Y(_07514_));
 sg13g2_xor2_1 _17648_ (.B(_07513_),
    .A(_07511_),
    .X(_07515_));
 sg13g2_xnor2_1 _17649_ (.Y(_07516_),
    .A(_07509_),
    .B(_07515_));
 sg13g2_nand2_1 _17650_ (.Y(_07517_),
    .A(_07507_),
    .B(_07516_));
 sg13g2_xor2_1 _17651_ (.B(_07516_),
    .A(_07507_),
    .X(_07518_));
 sg13g2_nand2_1 _17652_ (.Y(_07520_),
    .A(_07505_),
    .B(_07517_));
 sg13g2_o21ai_1 _17653_ (.B1(_07520_),
    .Y(_07521_),
    .A1(_07507_),
    .A2(_07516_));
 sg13g2_xnor2_1 _17654_ (.Y(_07522_),
    .A(_07505_),
    .B(_07518_));
 sg13g2_xnor2_1 _17655_ (.Y(_07523_),
    .A(_07496_),
    .B(_07522_));
 sg13g2_nor2_1 _17656_ (.A(_07473_),
    .B(_07523_),
    .Y(_07524_));
 sg13g2_xnor2_1 _17657_ (.Y(_07525_),
    .A(_07473_),
    .B(_07523_));
 sg13g2_nand2b_1 _17658_ (.Y(_07526_),
    .B(_07290_),
    .A_N(_07289_));
 sg13g2_xnor2_1 _17659_ (.Y(_07527_),
    .A(_07298_),
    .B(_07526_));
 sg13g2_xnor2_1 _17660_ (.Y(_07528_),
    .A(_07525_),
    .B(_07527_));
 sg13g2_a21oi_2 _17661_ (.B1(_05752_),
    .Y(_07529_),
    .A2(_05754_),
    .A1(_05751_));
 sg13g2_a21oi_1 _17662_ (.A1(_07473_),
    .A2(_07523_),
    .Y(_07531_),
    .B1(_07527_));
 sg13g2_nor2_1 _17663_ (.A(_07524_),
    .B(_07531_),
    .Y(_07532_));
 sg13g2_o21ai_1 _17664_ (.B1(_07532_),
    .Y(_07533_),
    .A1(_07528_),
    .A2(_07529_));
 sg13g2_or3_1 _17665_ (.A(_07528_),
    .B(_07529_),
    .C(_07532_),
    .X(_07534_));
 sg13g2_nor2_1 _17666_ (.A(_07495_),
    .B(_07522_),
    .Y(_07535_));
 sg13g2_a21oi_1 _17667_ (.A1(_07483_),
    .A2(_07494_),
    .Y(_07536_),
    .B1(_07535_));
 sg13g2_and3_1 _17668_ (.X(_07537_),
    .A(_07533_),
    .B(_07534_),
    .C(_07536_));
 sg13g2_a21oi_1 _17669_ (.A1(_07533_),
    .A2(_07534_),
    .Y(_07538_),
    .B1(_07536_));
 sg13g2_nand2_1 _17670_ (.Y(_07539_),
    .A(_07414_),
    .B(_07471_));
 sg13g2_o21ai_1 _17671_ (.B1(_07479_),
    .Y(_07540_),
    .A1(_07478_),
    .A2(_07482_));
 sg13g2_nand3_1 _17672_ (.B(_07539_),
    .C(_07540_),
    .A(_07470_),
    .Y(_07542_));
 sg13g2_a21o_1 _17673_ (.A2(_07539_),
    .A1(_07470_),
    .B1(_07540_),
    .X(_07543_));
 sg13g2_nand2_1 _17674_ (.Y(_07544_),
    .A(_07542_),
    .B(_07543_));
 sg13g2_nand2_1 _17675_ (.Y(_07545_),
    .A(_07489_),
    .B(_07492_));
 sg13g2_o21ai_1 _17676_ (.B1(_07545_),
    .Y(_07546_),
    .A1(_07485_),
    .A2(_07488_));
 sg13g2_nand2_1 _17677_ (.Y(_07547_),
    .A(_07543_),
    .B(_07546_));
 sg13g2_xor2_1 _17678_ (.B(_07546_),
    .A(_07544_),
    .X(_07548_));
 sg13g2_or3_1 _17679_ (.A(_07537_),
    .B(_07538_),
    .C(_07548_),
    .X(_07549_));
 sg13g2_o21ai_1 _17680_ (.B1(_07548_),
    .Y(_07550_),
    .A1(_07537_),
    .A2(_07538_));
 sg13g2_nor2_1 _17681_ (.A(_07432_),
    .B(_07443_),
    .Y(_07551_));
 sg13g2_nor3_1 _17682_ (.A(_07433_),
    .B(_07521_),
    .C(_07551_),
    .Y(_07553_));
 sg13g2_o21ai_1 _17683_ (.B1(_07521_),
    .Y(_07554_),
    .A1(_07433_),
    .A2(_07551_));
 sg13g2_nand2b_1 _17684_ (.Y(_07555_),
    .B(_07554_),
    .A_N(_07553_));
 sg13g2_o21ai_1 _17685_ (.B1(_07466_),
    .Y(_07556_),
    .A1(_07449_),
    .A2(_07467_));
 sg13g2_xnor2_1 _17686_ (.Y(_07557_),
    .A(_07555_),
    .B(_07556_));
 sg13g2_and3_1 _17687_ (.X(_07558_),
    .A(_07549_),
    .B(_07550_),
    .C(_07557_));
 sg13g2_a21oi_1 _17688_ (.A1(_07549_),
    .A2(_07550_),
    .Y(_07559_),
    .B1(_07557_));
 sg13g2_or3_1 _17689_ (.A(_07412_),
    .B(_07558_),
    .C(_07559_),
    .X(_07560_));
 sg13g2_o21ai_1 _17690_ (.B1(_07412_),
    .Y(_07561_),
    .A1(_07558_),
    .A2(_07559_));
 sg13g2_a21oi_1 _17691_ (.A1(_07511_),
    .A2(_07513_),
    .Y(_07562_),
    .B1(_07509_));
 sg13g2_nor2_2 _17692_ (.A(_07514_),
    .B(_07562_),
    .Y(_07564_));
 sg13g2_or3_1 _17693_ (.A(_07499_),
    .B(_07504_),
    .C(_07564_),
    .X(_07565_));
 sg13g2_o21ai_1 _17694_ (.B1(_07564_),
    .Y(_07566_),
    .A1(_07499_),
    .A2(_07504_));
 sg13g2_nand2_1 _17695_ (.Y(_07567_),
    .A(_07565_),
    .B(_07566_));
 sg13g2_o21ai_1 _17696_ (.B1(_07427_),
    .Y(_07568_),
    .A1(_07426_),
    .A2(_07429_));
 sg13g2_xnor2_1 _17697_ (.Y(_07569_),
    .A(_07567_),
    .B(_07568_));
 sg13g2_a21oi_2 _17698_ (.B1(_07438_),
    .Y(_07570_),
    .A2(_07441_),
    .A1(_07437_));
 sg13g2_nor3_1 _17699_ (.A(_07419_),
    .B(_07422_),
    .C(_07570_),
    .Y(_07571_));
 sg13g2_o21ai_1 _17700_ (.B1(_07570_),
    .Y(_07572_),
    .A1(_07419_),
    .A2(_07422_));
 sg13g2_nor2b_1 _17701_ (.A(_07571_),
    .B_N(_07572_),
    .Y(_07573_));
 sg13g2_nand2_1 _17702_ (.Y(_07575_),
    .A(_07454_),
    .B(_07457_));
 sg13g2_nand2_1 _17703_ (.Y(_07576_),
    .A(_07452_),
    .B(_07575_));
 sg13g2_xnor2_1 _17704_ (.Y(_07577_),
    .A(_07573_),
    .B(_07576_));
 sg13g2_nor2_1 _17705_ (.A(_07569_),
    .B(_07577_),
    .Y(_07578_));
 sg13g2_nand2_1 _17706_ (.Y(_07579_),
    .A(_07569_),
    .B(_07577_));
 sg13g2_nand2b_1 _17707_ (.Y(_07580_),
    .B(_07579_),
    .A_N(_07578_));
 sg13g2_a21o_1 _17708_ (.A2(_07447_),
    .A1(_06170_),
    .B1(_07446_),
    .X(_07581_));
 sg13g2_o21ai_1 _17709_ (.B1(_07581_),
    .Y(_07582_),
    .A1(_06170_),
    .A2(_07447_));
 sg13g2_nand2_1 _17710_ (.Y(_07583_),
    .A(_07461_),
    .B(_07463_));
 sg13g2_nand2_1 _17711_ (.Y(_07584_),
    .A(_07460_),
    .B(_07583_));
 sg13g2_nor2_1 _17712_ (.A(_07582_),
    .B(_07584_),
    .Y(_07586_));
 sg13g2_xor2_1 _17713_ (.B(_07584_),
    .A(_07582_),
    .X(_07587_));
 sg13g2_a21o_1 _17714_ (.A2(_07306_),
    .A1(_07303_),
    .B1(_07304_),
    .X(_07588_));
 sg13g2_xnor2_1 _17715_ (.Y(_07589_),
    .A(_07587_),
    .B(_07588_));
 sg13g2_xnor2_1 _17716_ (.Y(_07590_),
    .A(_07580_),
    .B(_07589_));
 sg13g2_and3_1 _17717_ (.X(_07591_),
    .A(_07560_),
    .B(_07561_),
    .C(_07590_));
 sg13g2_a21oi_1 _17718_ (.A1(_07560_),
    .A2(_07561_),
    .Y(_07592_),
    .B1(_07590_));
 sg13g2_or2_1 _17719_ (.X(_07593_),
    .B(_07592_),
    .A(_07591_));
 sg13g2_o21ai_1 _17720_ (.B1(_07401_),
    .Y(_07594_),
    .A1(_07591_),
    .A2(_07592_));
 sg13g2_nand2_1 _17721_ (.Y(_07595_),
    .A(_07561_),
    .B(_07590_));
 sg13g2_and2_1 _17722_ (.A(_07560_),
    .B(_07595_),
    .X(_07597_));
 sg13g2_a21o_1 _17723_ (.A2(_07593_),
    .A1(_07401_),
    .B1(_07597_),
    .X(_07598_));
 sg13g2_nor2b_1 _17724_ (.A(_07594_),
    .B_N(_07597_),
    .Y(_07599_));
 sg13g2_xnor2_1 _17725_ (.Y(_07600_),
    .A(_07594_),
    .B(_07597_));
 sg13g2_nand2_1 _17726_ (.Y(_07601_),
    .A(_07550_),
    .B(_07557_));
 sg13g2_and2_1 _17727_ (.A(_07549_),
    .B(_07601_),
    .X(_07602_));
 sg13g2_xnor2_1 _17728_ (.Y(_07603_),
    .A(_07600_),
    .B(_07602_));
 sg13g2_a21oi_1 _17729_ (.A1(_07407_),
    .A2(_07411_),
    .Y(_07604_),
    .B1(_07406_));
 sg13g2_o21ai_1 _17730_ (.B1(_07579_),
    .Y(_07605_),
    .A1(_07578_),
    .A2(_07589_));
 sg13g2_nand2b_1 _17731_ (.Y(_07606_),
    .B(_07604_),
    .A_N(_07605_));
 sg13g2_nand2b_1 _17732_ (.Y(_07608_),
    .B(_07605_),
    .A_N(_07604_));
 sg13g2_nand2_1 _17733_ (.Y(_07609_),
    .A(_07606_),
    .B(_07608_));
 sg13g2_o21ai_1 _17734_ (.B1(_07400_),
    .Y(_07610_),
    .A1(_07286_),
    .A2(_07395_));
 sg13g2_nand2_2 _17735_ (.Y(_07611_),
    .A(_07396_),
    .B(_07610_));
 sg13g2_xnor2_1 _17736_ (.Y(_07612_),
    .A(_07609_),
    .B(_07611_));
 sg13g2_and2_1 _17737_ (.A(_07603_),
    .B(_07612_),
    .X(_07613_));
 sg13g2_or2_1 _17738_ (.X(_07614_),
    .B(_07612_),
    .A(_07603_));
 sg13g2_xor2_1 _17739_ (.B(_07612_),
    .A(_07603_),
    .X(_07615_));
 sg13g2_o21ai_1 _17740_ (.B1(_07554_),
    .Y(_07616_),
    .A1(_07553_),
    .A2(_07556_));
 sg13g2_nand2_1 _17741_ (.Y(_07617_),
    .A(_07542_),
    .B(_07547_));
 sg13g2_nand2_1 _17742_ (.Y(_07619_),
    .A(_07534_),
    .B(_07536_));
 sg13g2_nand2_1 _17743_ (.Y(_07620_),
    .A(_07533_),
    .B(_07619_));
 sg13g2_nand2_1 _17744_ (.Y(_07621_),
    .A(_07617_),
    .B(_07620_));
 sg13g2_inv_1 _17745_ (.Y(_07622_),
    .A(_07621_));
 sg13g2_nor2_1 _17746_ (.A(_07617_),
    .B(_07620_),
    .Y(_07623_));
 sg13g2_nor2_1 _17747_ (.A(_07622_),
    .B(_07623_),
    .Y(_07624_));
 sg13g2_xnor2_1 _17748_ (.Y(_07625_),
    .A(_07616_),
    .B(_07624_));
 sg13g2_xnor2_1 _17749_ (.Y(_07626_),
    .A(_07615_),
    .B(_07625_));
 sg13g2_or2_1 _17750_ (.X(_07627_),
    .B(_07576_),
    .A(_07571_));
 sg13g2_nand2_1 _17751_ (.Y(_07628_),
    .A(_07565_),
    .B(_07568_));
 sg13g2_and2_1 _17752_ (.A(_07566_),
    .B(_07628_),
    .X(_07630_));
 sg13g2_and3_1 _17753_ (.X(_07631_),
    .A(_07572_),
    .B(_07627_),
    .C(_07630_));
 sg13g2_a21o_1 _17754_ (.A2(_07627_),
    .A1(_07572_),
    .B1(_07630_),
    .X(_07632_));
 sg13g2_nand2b_1 _17755_ (.Y(_07633_),
    .B(_07632_),
    .A_N(_07631_));
 sg13g2_nor2_1 _17756_ (.A(_07586_),
    .B(_07588_),
    .Y(_07634_));
 sg13g2_a21o_1 _17757_ (.A2(_07584_),
    .A1(_07582_),
    .B1(_07634_),
    .X(_07635_));
 sg13g2_xnor2_1 _17758_ (.Y(_07636_),
    .A(_07633_),
    .B(_07635_));
 sg13g2_nand2b_1 _17759_ (.Y(_07637_),
    .B(_07360_),
    .A_N(_07385_));
 sg13g2_a22oi_1 _17760_ (.Y(_07638_),
    .B1(_07388_),
    .B2(_07637_),
    .A2(_07386_),
    .A1(_07385_));
 sg13g2_or2_1 _17761_ (.X(_07639_),
    .B(_07638_),
    .A(_07636_));
 sg13g2_nand2_1 _17762_ (.Y(_07641_),
    .A(_07636_),
    .B(_07638_));
 sg13g2_nand2_1 _17763_ (.Y(_07642_),
    .A(_07639_),
    .B(_07641_));
 sg13g2_xor2_1 _17764_ (.B(_07642_),
    .A(_07393_),
    .X(_07643_));
 sg13g2_inv_1 _17765_ (.Y(_07644_),
    .A(_07643_));
 sg13g2_o21ai_1 _17766_ (.B1(_07614_),
    .Y(_07645_),
    .A1(_07613_),
    .A2(_07625_));
 sg13g2_a21o_1 _17767_ (.A2(_07644_),
    .A1(_07626_),
    .B1(_07645_),
    .X(_07646_));
 sg13g2_nor3_1 _17768_ (.A(_07614_),
    .B(_07625_),
    .C(_07643_),
    .Y(_07647_));
 sg13g2_inv_1 _17769_ (.Y(_07648_),
    .A(_07647_));
 sg13g2_nand2_1 _17770_ (.Y(_07649_),
    .A(_07393_),
    .B(_07641_));
 sg13g2_nand2_1 _17771_ (.Y(_07650_),
    .A(_07639_),
    .B(_07649_));
 sg13g2_and4_1 _17772_ (.A(_07639_),
    .B(_07646_),
    .C(_07648_),
    .D(_07649_),
    .X(_07652_));
 sg13g2_a22oi_1 _17773_ (.Y(_07653_),
    .B1(_07649_),
    .B2(_07639_),
    .A2(_07648_),
    .A1(_07646_));
 sg13g2_a21oi_2 _17774_ (.B1(_07623_),
    .Y(_07654_),
    .A2(_07621_),
    .A1(_07616_));
 sg13g2_nand2_1 _17775_ (.Y(_07655_),
    .A(_07608_),
    .B(_07611_));
 sg13g2_nand2_1 _17776_ (.Y(_07656_),
    .A(_07606_),
    .B(_07655_));
 sg13g2_a21oi_2 _17777_ (.B1(_07599_),
    .Y(_07657_),
    .A2(_07602_),
    .A1(_07598_));
 sg13g2_nor2_1 _17778_ (.A(_07656_),
    .B(_07657_),
    .Y(_07658_));
 sg13g2_xor2_1 _17779_ (.B(_07657_),
    .A(_07656_),
    .X(_07659_));
 sg13g2_xnor2_1 _17780_ (.Y(_07660_),
    .A(_07654_),
    .B(_07659_));
 sg13g2_o21ai_1 _17781_ (.B1(_07660_),
    .Y(_07661_),
    .A1(_07652_),
    .A2(_07653_));
 sg13g2_or3_1 _17782_ (.A(_07652_),
    .B(_07653_),
    .C(_07660_),
    .X(_07663_));
 sg13g2_nand2_1 _17783_ (.Y(_07664_),
    .A(_07389_),
    .B(_07663_));
 sg13g2_and3_1 _17784_ (.X(_07665_),
    .A(_07389_),
    .B(_07661_),
    .C(_07663_));
 sg13g2_a21oi_1 _17785_ (.A1(_07661_),
    .A2(_07663_),
    .Y(_07666_),
    .B1(_07389_));
 sg13g2_nor2_1 _17786_ (.A(_07665_),
    .B(_07666_),
    .Y(_07667_));
 sg13g2_o21ai_1 _17787_ (.B1(_07632_),
    .Y(_07668_),
    .A1(_07631_),
    .A2(_07635_));
 sg13g2_inv_1 _17788_ (.Y(_07669_),
    .A(_07668_));
 sg13g2_nor3_1 _17789_ (.A(_07665_),
    .B(_07666_),
    .C(_07669_),
    .Y(_07670_));
 sg13g2_nand2_1 _17790_ (.Y(_07671_),
    .A(_07661_),
    .B(_07664_));
 sg13g2_nor3_1 _17791_ (.A(_07388_),
    .B(_07661_),
    .C(_07669_),
    .Y(_07672_));
 sg13g2_xnor2_1 _17792_ (.Y(_07674_),
    .A(_07670_),
    .B(_07671_));
 sg13g2_a21oi_2 _17793_ (.B1(_07647_),
    .Y(_07675_),
    .A2(_07650_),
    .A1(_07646_));
 sg13g2_xnor2_1 _17794_ (.Y(_07676_),
    .A(_07674_),
    .B(_07675_));
 sg13g2_a21oi_1 _17795_ (.A1(_07656_),
    .A2(_07657_),
    .Y(_07677_),
    .B1(_07654_));
 sg13g2_nor2_2 _17796_ (.A(_07658_),
    .B(_07677_),
    .Y(_07678_));
 sg13g2_nand2b_1 _17797_ (.Y(_07679_),
    .B(_07675_),
    .A_N(_07672_));
 sg13g2_o21ai_1 _17798_ (.B1(_07679_),
    .Y(_07680_),
    .A1(_07670_),
    .A2(_07671_));
 sg13g2_o21ai_1 _17799_ (.B1(_07680_),
    .Y(_07681_),
    .A1(_07676_),
    .A2(_07678_));
 sg13g2_nor2_1 _17800_ (.A(_07271_),
    .B(net9),
    .Y(_07682_));
 sg13g2_nand2b_1 _17801_ (.Y(_07683_),
    .B(_07272_),
    .A_N(net9));
 sg13g2_or3_2 _17802_ (.A(_07264_),
    .B(_07265_),
    .C(_07268_),
    .X(_07685_));
 sg13g2_nand2_1 _17803_ (.Y(_07686_),
    .A(_07269_),
    .B(_07685_));
 sg13g2_xnor2_1 _17804_ (.Y(_07687_),
    .A(_06625_),
    .B(_07257_));
 sg13g2_xnor2_1 _17805_ (.Y(_07688_),
    .A(_07667_),
    .B(_07668_));
 sg13g2_xnor2_1 _17806_ (.Y(_07689_),
    .A(_07626_),
    .B(_07644_));
 sg13g2_a21oi_1 _17807_ (.A1(_07242_),
    .A2(_07243_),
    .Y(_07690_),
    .B1(_07230_));
 sg13g2_nor2_2 _17808_ (.A(_07245_),
    .B(_07690_),
    .Y(_07691_));
 sg13g2_xnor2_1 _17809_ (.Y(_07692_),
    .A(_07401_),
    .B(_07593_));
 sg13g2_inv_8 _17810_ (.Y(_07693_),
    .A(_07692_));
 sg13g2_xnor2_1 _17811_ (.Y(_07694_),
    .A(_07120_),
    .B(_07122_));
 sg13g2_inv_1 _17812_ (.Y(_07696_),
    .A(_07694_));
 sg13g2_xnor2_1 _17813_ (.Y(_07697_),
    .A(_07528_),
    .B(_07529_));
 sg13g2_inv_1 _17814_ (.Y(_07698_),
    .A(_07697_));
 sg13g2_xnor2_1 _17815_ (.Y(_07699_),
    .A(_06994_),
    .B(_07005_));
 sg13g2_nand2_1 _17816_ (.Y(_07700_),
    .A(_06269_),
    .B(_07699_));
 sg13g2_o21ai_1 _17817_ (.B1(_07700_),
    .Y(_07701_),
    .A1(_07694_),
    .A2(_07698_));
 sg13g2_o21ai_1 _17818_ (.B1(_07701_),
    .Y(_07702_),
    .A1(_07696_),
    .A2(_07697_));
 sg13g2_xnor2_1 _17819_ (.Y(_07703_),
    .A(_07191_),
    .B(_07194_));
 sg13g2_o21ai_1 _17820_ (.B1(_07703_),
    .Y(_07704_),
    .A1(_07693_),
    .A2(_07702_));
 sg13g2_o21ai_1 _17821_ (.B1(_07704_),
    .Y(_07705_),
    .A1(_07689_),
    .A2(_07691_));
 sg13g2_a21oi_1 _17822_ (.A1(_07693_),
    .A2(_07702_),
    .Y(_07707_),
    .B1(_07705_));
 sg13g2_a221oi_1 _17823_ (.B2(_07691_),
    .C1(_07707_),
    .B1(_07689_),
    .A1(_07687_),
    .Y(_07708_),
    .A2(_07688_));
 sg13g2_nor2_1 _17824_ (.A(_07687_),
    .B(_07688_),
    .Y(_07709_));
 sg13g2_nor2_2 _17825_ (.A(_07708_),
    .B(_07709_),
    .Y(_07710_));
 sg13g2_xnor2_1 _17826_ (.Y(_07711_),
    .A(_07676_),
    .B(_07678_));
 sg13g2_nand2_1 _17827_ (.Y(_07712_),
    .A(_07710_),
    .B(_07711_));
 sg13g2_a22oi_1 _17828_ (.Y(_07713_),
    .B1(_07710_),
    .B2(_07711_),
    .A2(_07685_),
    .A1(_07269_));
 sg13g2_nand3_1 _17829_ (.B(_07270_),
    .C(net9),
    .A(_07269_),
    .Y(_07714_));
 sg13g2_nor2_1 _17830_ (.A(_07710_),
    .B(_07711_),
    .Y(_07715_));
 sg13g2_or2_1 _17831_ (.X(_07716_),
    .B(_07711_),
    .A(_07710_));
 sg13g2_a221oi_1 _17832_ (.B2(_07712_),
    .C1(_07715_),
    .B1(_07686_),
    .A1(_07271_),
    .Y(_07718_),
    .A2(net9));
 sg13g2_nand3b_1 _17833_ (.B(_07714_),
    .C(_07716_),
    .Y(_07719_),
    .A_N(_07713_));
 sg13g2_nor2_1 _17834_ (.A(_07682_),
    .B(_07718_),
    .Y(_07720_));
 sg13g2_a21o_1 _17835_ (.A2(net2170),
    .A1(net2171),
    .B1(_07699_),
    .X(_07721_));
 sg13g2_nand3_1 _17836_ (.B(net2171),
    .C(net2169),
    .A(_06269_),
    .Y(_07722_));
 sg13g2_nand2_1 _17837_ (.Y(_07723_),
    .A(_07721_),
    .B(_07722_));
 sg13g2_xor2_1 _17838_ (.B(net2279),
    .A(net2215),
    .X(_07724_));
 sg13g2_nor2_1 _17839_ (.A(net2728),
    .B(net2249),
    .Y(_07725_));
 sg13g2_nor2_1 _17840_ (.A(net2553),
    .B(net2328),
    .Y(_07726_));
 sg13g2_xnor2_1 _17841_ (.Y(_07727_),
    .A(_07725_),
    .B(_07726_));
 sg13g2_nand2_1 _17842_ (.Y(_07729_),
    .A(_07724_),
    .B(_07727_));
 sg13g2_nor2_1 _17843_ (.A(_07724_),
    .B(_07727_),
    .Y(_07730_));
 sg13g2_xnor2_1 _17844_ (.Y(_07731_),
    .A(net2276),
    .B(net2776));
 sg13g2_nand2_1 _17845_ (.Y(_07732_),
    .A(_07729_),
    .B(_07731_));
 sg13g2_inv_1 _17846_ (.Y(_07733_),
    .A(_07732_));
 sg13g2_xnor2_1 _17847_ (.Y(_07734_),
    .A(net2673),
    .B(net2790));
 sg13g2_xnor2_1 _17848_ (.Y(_07735_),
    .A(net2300),
    .B(net2220));
 sg13g2_xnor2_1 _17849_ (.Y(_07736_),
    .A(net2482),
    .B(net2292));
 sg13g2_o21ai_1 _17850_ (.B1(_07736_),
    .Y(_07737_),
    .A1(_07734_),
    .A2(_07735_));
 sg13g2_or3_1 _17851_ (.A(_07734_),
    .B(_07735_),
    .C(_07736_),
    .X(_07738_));
 sg13g2_nor2_1 _17852_ (.A(net2587),
    .B(net2270),
    .Y(_07740_));
 sg13g2_xnor2_1 _17853_ (.Y(_07741_),
    .A(_01204_),
    .B(_07740_));
 sg13g2_nand2_1 _17854_ (.Y(_07742_),
    .A(_07737_),
    .B(_07741_));
 sg13g2_and2_1 _17855_ (.A(_07738_),
    .B(_07742_),
    .X(_07743_));
 sg13g2_o21ai_1 _17856_ (.B1(_07743_),
    .Y(_07744_),
    .A1(_07730_),
    .A2(_07733_));
 sg13g2_or3_1 _17857_ (.A(_07730_),
    .B(_07733_),
    .C(_07743_),
    .X(_07745_));
 sg13g2_inv_1 _17858_ (.Y(_07746_),
    .A(_07745_));
 sg13g2_nor2_1 _17859_ (.A(net2792),
    .B(net2466),
    .Y(_07747_));
 sg13g2_xnor2_1 _17860_ (.Y(_07748_),
    .A(net2756),
    .B(_07747_));
 sg13g2_nor2_1 _17861_ (.A(net2562),
    .B(net2245),
    .Y(_07749_));
 sg13g2_nor2b_1 _17862_ (.A(net2655),
    .B_N(net2421),
    .Y(_07751_));
 sg13g2_xnor2_1 _17863_ (.Y(_07752_),
    .A(_07749_),
    .B(_07751_));
 sg13g2_nor2b_1 _17864_ (.A(_07748_),
    .B_N(_07752_),
    .Y(_07753_));
 sg13g2_nand2b_1 _17865_ (.Y(_07754_),
    .B(_07748_),
    .A_N(_07752_));
 sg13g2_xnor2_1 _17866_ (.Y(_07755_),
    .A(net2764),
    .B(net2309));
 sg13g2_xor2_1 _17867_ (.B(net2461),
    .A(net2677),
    .X(_07756_));
 sg13g2_nand2_1 _17868_ (.Y(_07757_),
    .A(_07755_),
    .B(_07756_));
 sg13g2_o21ai_1 _17869_ (.B1(_07754_),
    .Y(_07758_),
    .A1(_07753_),
    .A2(_07757_));
 sg13g2_a21oi_1 _17870_ (.A1(_07744_),
    .A2(_07758_),
    .Y(_07759_),
    .B1(_07746_));
 sg13g2_nor2b_2 _17871_ (.A(net2642),
    .B_N(net2382),
    .Y(_07760_));
 sg13g2_or3_1 _17872_ (.A(net2215),
    .B(net2244),
    .C(_07760_),
    .X(_07762_));
 sg13g2_xor2_1 _17873_ (.B(net2734),
    .A(net2816),
    .X(_07763_));
 sg13g2_xor2_1 _17874_ (.B(net2746),
    .A(net2609),
    .X(_07764_));
 sg13g2_nor2_2 _17875_ (.A(_07763_),
    .B(_07764_),
    .Y(_07765_));
 sg13g2_nor2b_1 _17876_ (.A(net2244),
    .B_N(net2215),
    .Y(_07766_));
 sg13g2_mux2_1 _17877_ (.A0(net2244),
    .A1(_07766_),
    .S(_07760_),
    .X(_07767_));
 sg13g2_o21ai_1 _17878_ (.B1(_07762_),
    .Y(_07768_),
    .A1(_07765_),
    .A2(_07767_));
 sg13g2_o21ai_1 _17879_ (.B1(net2471),
    .Y(_07769_),
    .A1(net2332),
    .A2(net2265));
 sg13g2_xor2_1 _17880_ (.B(net2618),
    .A(net2751),
    .X(_07770_));
 sg13g2_nor3_1 _17881_ (.A(net2413),
    .B(_07769_),
    .C(_07770_),
    .Y(_07771_));
 sg13g2_o21ai_1 _17882_ (.B1(_07770_),
    .Y(_07773_),
    .A1(net2413),
    .A2(_07769_));
 sg13g2_xnor2_1 _17883_ (.Y(_07774_),
    .A(net2255),
    .B(net2746));
 sg13g2_nand3_1 _17884_ (.B(_05924_),
    .C(_07774_),
    .A(_05154_),
    .Y(_07775_));
 sg13g2_o21ai_1 _17885_ (.B1(_07773_),
    .Y(_07776_),
    .A1(_07771_),
    .A2(_07775_));
 sg13g2_nand2_1 _17886_ (.Y(_07777_),
    .A(_07768_),
    .B(_07776_));
 sg13g2_or2_1 _17887_ (.X(_07778_),
    .B(_07776_),
    .A(_07768_));
 sg13g2_nor2_1 _17888_ (.A(net2484),
    .B(net2609),
    .Y(_07779_));
 sg13g2_nor2b_1 _17889_ (.A(net2394),
    .B_N(net2292),
    .Y(_07780_));
 sg13g2_nor2_1 _17890_ (.A(net2397),
    .B(net2799),
    .Y(_07781_));
 sg13g2_xor2_1 _17891_ (.B(net2790),
    .A(net2235),
    .X(_07782_));
 sg13g2_a22oi_1 _17892_ (.Y(_07784_),
    .B1(_07781_),
    .B2(_07782_),
    .A2(_07780_),
    .A1(_07779_));
 sg13g2_nand4_1 _17893_ (.B(_07780_),
    .C(_07781_),
    .A(_07779_),
    .Y(_07785_),
    .D(_07782_));
 sg13g2_xor2_1 _17894_ (.B(net2277),
    .A(net2215),
    .X(_07786_));
 sg13g2_nor2_1 _17895_ (.A(_06573_),
    .B(_07786_),
    .Y(_07787_));
 sg13g2_o21ai_1 _17896_ (.B1(_07785_),
    .Y(_07788_),
    .A1(_07784_),
    .A2(_07787_));
 sg13g2_nand2_1 _17897_ (.Y(_07789_),
    .A(_07777_),
    .B(_07788_));
 sg13g2_nand3_1 _17898_ (.B(_07778_),
    .C(_07789_),
    .A(_07759_),
    .Y(_07790_));
 sg13g2_a21o_2 _17899_ (.A2(_07789_),
    .A1(_07778_),
    .B1(_07759_),
    .X(_07791_));
 sg13g2_xor2_1 _17900_ (.B(net2748),
    .A(net2786),
    .X(_07792_));
 sg13g2_xor2_1 _17901_ (.B(net2255),
    .A(net2349),
    .X(_07793_));
 sg13g2_nand2_1 _17902_ (.Y(_07795_),
    .A(_07792_),
    .B(_07793_));
 sg13g2_or2_1 _17903_ (.X(_07796_),
    .B(_07793_),
    .A(_07792_));
 sg13g2_nor2_1 _17904_ (.A(_05187_),
    .B(net2461),
    .Y(_07797_));
 sg13g2_nor2_1 _17905_ (.A(net2289),
    .B(net2713),
    .Y(_07798_));
 sg13g2_xnor2_1 _17906_ (.Y(_07799_),
    .A(_07797_),
    .B(_07798_));
 sg13g2_nand2_1 _17907_ (.Y(_07800_),
    .A(_07795_),
    .B(_07799_));
 sg13g2_nand2_1 _17908_ (.Y(_07801_),
    .A(_07796_),
    .B(_07800_));
 sg13g2_xor2_1 _17909_ (.B(net2624),
    .A(net2793),
    .X(_07802_));
 sg13g2_nor2_2 _17910_ (.A(net2230),
    .B(net2458),
    .Y(_07803_));
 sg13g2_xor2_1 _17911_ (.B(_07803_),
    .A(_00846_),
    .X(_07804_));
 sg13g2_nand2b_1 _17912_ (.Y(_07806_),
    .B(_07802_),
    .A_N(_07804_));
 sg13g2_nor2b_1 _17913_ (.A(_07802_),
    .B_N(_07804_),
    .Y(_07807_));
 sg13g2_nor2_1 _17914_ (.A(net2786),
    .B(net2790),
    .Y(_07808_));
 sg13g2_nor2_1 _17915_ (.A(net2277),
    .B(net2682),
    .Y(_07809_));
 sg13g2_xor2_1 _17916_ (.B(_07809_),
    .A(_07808_),
    .X(_07810_));
 sg13g2_a21o_1 _17917_ (.A2(_07810_),
    .A1(_07806_),
    .B1(_07807_),
    .X(_07811_));
 sg13g2_or2_1 _17918_ (.X(_07812_),
    .B(_07811_),
    .A(_07801_));
 sg13g2_and2_1 _17919_ (.A(_07801_),
    .B(_07811_),
    .X(_07813_));
 sg13g2_nor2_1 _17920_ (.A(net2415),
    .B(net2799),
    .Y(_07814_));
 sg13g2_xnor2_1 _17921_ (.Y(_07815_),
    .A(net2618),
    .B(_07814_));
 sg13g2_nor2_1 _17922_ (.A(net2214),
    .B(net2731),
    .Y(_07817_));
 sg13g2_xnor2_1 _17923_ (.Y(_07818_),
    .A(_00022_),
    .B(_07817_));
 sg13g2_nand2_1 _17924_ (.Y(_07819_),
    .A(_07815_),
    .B(_07818_));
 sg13g2_nor2_1 _17925_ (.A(_07815_),
    .B(_07818_),
    .Y(_07820_));
 sg13g2_xnor2_1 _17926_ (.Y(_07821_),
    .A(net2576),
    .B(net2271));
 sg13g2_xor2_1 _17927_ (.B(net2368),
    .A(net2614),
    .X(_07822_));
 sg13g2_nor2_2 _17928_ (.A(_07821_),
    .B(_07822_),
    .Y(_07823_));
 sg13g2_a21oi_2 _17929_ (.B1(_07820_),
    .Y(_07824_),
    .A2(_07823_),
    .A1(_07819_));
 sg13g2_a21oi_2 _17930_ (.B1(_07813_),
    .Y(_07825_),
    .A2(_07824_),
    .A1(_07812_));
 sg13g2_nand2_1 _17931_ (.Y(_07826_),
    .A(_07790_),
    .B(_07825_));
 sg13g2_nor2_1 _17932_ (.A(net2634),
    .B(net2274),
    .Y(_07828_));
 sg13g2_xor2_1 _17933_ (.B(net2274),
    .A(net2634),
    .X(_07829_));
 sg13g2_nor2_1 _17934_ (.A(net2482),
    .B(net2394),
    .Y(_07830_));
 sg13g2_xnor2_1 _17935_ (.Y(_07831_),
    .A(net2232),
    .B(net2740));
 sg13g2_nand2_1 _17936_ (.Y(_07832_),
    .A(_07830_),
    .B(_07831_));
 sg13g2_nor2_1 _17937_ (.A(net2587),
    .B(net2249),
    .Y(_07833_));
 sg13g2_nor2_1 _17938_ (.A(net2447),
    .B(net2287),
    .Y(_07834_));
 sg13g2_xnor2_1 _17939_ (.Y(_07835_),
    .A(_07833_),
    .B(_07834_));
 sg13g2_a21o_1 _17940_ (.A2(_07831_),
    .A1(_07830_),
    .B1(_07835_),
    .X(_07836_));
 sg13g2_nor2b_1 _17941_ (.A(_07832_),
    .B_N(_07835_),
    .Y(_07837_));
 sg13g2_xor2_1 _17942_ (.B(_07835_),
    .A(_07832_),
    .X(_07839_));
 sg13g2_xnor2_1 _17943_ (.Y(_07840_),
    .A(_07829_),
    .B(_07839_));
 sg13g2_or2_1 _17944_ (.X(_07841_),
    .B(net2597),
    .A(net2415));
 sg13g2_xnor2_1 _17945_ (.Y(_07842_),
    .A(net2245),
    .B(net2319));
 sg13g2_nor2_1 _17946_ (.A(_07841_),
    .B(_07842_),
    .Y(_07843_));
 sg13g2_xnor2_1 _17947_ (.Y(_07844_),
    .A(_07841_),
    .B(_07842_));
 sg13g2_xnor2_1 _17948_ (.Y(_07845_),
    .A(net2716),
    .B(net2690));
 sg13g2_xnor2_1 _17949_ (.Y(_07846_),
    .A(_07844_),
    .B(_07845_));
 sg13g2_inv_1 _17950_ (.Y(_07847_),
    .A(_07846_));
 sg13g2_nor2_1 _17951_ (.A(_07840_),
    .B(_07847_),
    .Y(_07848_));
 sg13g2_nor2_1 _17952_ (.A(net2413),
    .B(net2360),
    .Y(_07850_));
 sg13g2_xnor2_1 _17953_ (.Y(_07851_),
    .A(_00000_),
    .B(_07850_));
 sg13g2_xnor2_1 _17954_ (.Y(_07852_),
    .A(net2332),
    .B(net2222));
 sg13g2_nand2_1 _17955_ (.Y(_07853_),
    .A(_07851_),
    .B(_07852_));
 sg13g2_nor2_1 _17956_ (.A(_07851_),
    .B(_07852_),
    .Y(_07854_));
 sg13g2_xor2_1 _17957_ (.B(_07852_),
    .A(_07851_),
    .X(_07855_));
 sg13g2_nor2_2 _17958_ (.A(net2482),
    .B(net2673),
    .Y(_07856_));
 sg13g2_xor2_1 _17959_ (.B(net2203),
    .A(\net.in[96] ),
    .X(_07857_));
 sg13g2_xnor2_1 _17960_ (.Y(_07858_),
    .A(_07856_),
    .B(_07857_));
 sg13g2_xnor2_1 _17961_ (.Y(_07859_),
    .A(_07855_),
    .B(_07858_));
 sg13g2_a21oi_1 _17962_ (.A1(_07840_),
    .A2(_07847_),
    .Y(_07861_),
    .B1(_07859_));
 sg13g2_xnor2_1 _17963_ (.Y(_07862_),
    .A(net2764),
    .B(net2731));
 sg13g2_inv_1 _17964_ (.Y(_07863_),
    .A(_07862_));
 sg13g2_nand2b_1 _17965_ (.Y(_07864_),
    .B(net2799),
    .A_N(net2282));
 sg13g2_xnor2_1 _17966_ (.Y(_07865_),
    .A(net2694),
    .B(net2629));
 sg13g2_xnor2_1 _17967_ (.Y(_07866_),
    .A(_07864_),
    .B(_07865_));
 sg13g2_nand2_1 _17968_ (.Y(_07867_),
    .A(_07863_),
    .B(_07866_));
 sg13g2_nor2_1 _17969_ (.A(_07863_),
    .B(_07866_),
    .Y(_07868_));
 sg13g2_a22oi_1 _17970_ (.Y(_07869_),
    .B1(_05737_),
    .B2(net2237),
    .A2(net2809),
    .A1(net2180));
 sg13g2_o21ai_1 _17971_ (.B1(_07869_),
    .Y(_07870_),
    .A1(_05737_),
    .A2(net2237));
 sg13g2_a21oi_1 _17972_ (.A1(_07867_),
    .A2(_07870_),
    .Y(_07872_),
    .B1(_07868_));
 sg13g2_o21ai_1 _17973_ (.B1(_07872_),
    .Y(_07873_),
    .A1(_07848_),
    .A2(_07861_));
 sg13g2_or3_1 _17974_ (.A(_07848_),
    .B(_07861_),
    .C(_07872_),
    .X(_07874_));
 sg13g2_nor2_2 _17975_ (.A(net2662),
    .B(net2461),
    .Y(_07875_));
 sg13g2_or2_1 _17976_ (.X(_07876_),
    .B(net2235),
    .A(net2634));
 sg13g2_nand2_1 _17977_ (.Y(_07877_),
    .A(_07875_),
    .B(_07876_));
 sg13g2_nor2_1 _17978_ (.A(net2792),
    .B(net2245),
    .Y(_07878_));
 sg13g2_xnor2_1 _17979_ (.Y(_07879_),
    .A(net2792),
    .B(net2244));
 sg13g2_nor2b_1 _17980_ (.A(net2691),
    .B_N(net2623),
    .Y(_07880_));
 sg13g2_xnor2_1 _17981_ (.Y(_07881_),
    .A(_07879_),
    .B(_07880_));
 sg13g2_a21oi_1 _17982_ (.A1(_07875_),
    .A2(_07876_),
    .Y(_07883_),
    .B1(_07881_));
 sg13g2_nand2b_1 _17983_ (.Y(_07884_),
    .B(_07881_),
    .A_N(_07877_));
 sg13g2_or3_2 _17984_ (.A(net2372),
    .B(net2587),
    .C(net2800),
    .X(_07885_));
 sg13g2_o21ai_1 _17985_ (.B1(_07884_),
    .Y(_07886_),
    .A1(_07883_),
    .A2(_07885_));
 sg13g2_nand2_1 _17986_ (.Y(_07887_),
    .A(_07873_),
    .B(_07886_));
 sg13g2_nor2_2 _17987_ (.A(net2243),
    .B(net2193),
    .Y(_07888_));
 sg13g2_and2_1 _17988_ (.A(net2243),
    .B(net2190),
    .X(_07889_));
 sg13g2_xnor2_1 _17989_ (.Y(_07890_),
    .A(net2345),
    .B(net2252));
 sg13g2_o21ai_1 _17990_ (.B1(_07890_),
    .Y(_07891_),
    .A1(_07888_),
    .A2(_07889_));
 sg13g2_or3_1 _17991_ (.A(_07888_),
    .B(_07889_),
    .C(_07890_),
    .X(_07892_));
 sg13g2_nor2_1 _17992_ (.A(net2178),
    .B(net2690),
    .Y(_07894_));
 sg13g2_xnor2_1 _17993_ (.Y(_07895_),
    .A(_07878_),
    .B(_07894_));
 sg13g2_nand2_1 _17994_ (.Y(_07896_),
    .A(_07891_),
    .B(_07895_));
 sg13g2_and2_1 _17995_ (.A(_07892_),
    .B(_07896_),
    .X(_07897_));
 sg13g2_xor2_1 _17996_ (.B(net2289),
    .A(net2306),
    .X(_07898_));
 sg13g2_inv_1 _17997_ (.Y(_07899_),
    .A(_07898_));
 sg13g2_nor2_1 _17998_ (.A(net2193),
    .B(net2194),
    .Y(_07900_));
 sg13g2_nor2b_1 _17999_ (.A(net2699),
    .B_N(net2466),
    .Y(_07901_));
 sg13g2_xnor2_1 _18000_ (.Y(_07902_),
    .A(_07900_),
    .B(_07901_));
 sg13g2_nand2_1 _18001_ (.Y(_07903_),
    .A(_07899_),
    .B(_07902_));
 sg13g2_nor2_1 _18002_ (.A(_07899_),
    .B(_07902_),
    .Y(_07905_));
 sg13g2_nor2_1 _18003_ (.A(_05209_),
    .B(net2647),
    .Y(_07906_));
 sg13g2_xnor2_1 _18004_ (.Y(_07907_),
    .A(_00019_),
    .B(_07906_));
 sg13g2_a21oi_1 _18005_ (.A1(_07903_),
    .A2(_07907_),
    .Y(_07908_),
    .B1(_07905_));
 sg13g2_and2_1 _18006_ (.A(_07897_),
    .B(_07908_),
    .X(_07909_));
 sg13g2_nor2_1 _18007_ (.A(_07897_),
    .B(_07908_),
    .Y(_07910_));
 sg13g2_nor2_1 _18008_ (.A(net2178),
    .B(net2587),
    .Y(_07911_));
 sg13g2_xor2_1 _18009_ (.B(net2766),
    .A(net2329),
    .X(_07912_));
 sg13g2_o21ai_1 _18010_ (.B1(_07912_),
    .Y(_07913_),
    .A1(net2178),
    .A2(net2587));
 sg13g2_nor3_1 _18011_ (.A(net2178),
    .B(net2587),
    .C(_07912_),
    .Y(_07914_));
 sg13g2_nor2_1 _18012_ (.A(net2807),
    .B(net2805),
    .Y(_07916_));
 sg13g2_xnor2_1 _18013_ (.Y(_07917_),
    .A(\net.in[209] ),
    .B(_07916_));
 sg13g2_a21oi_1 _18014_ (.A1(_07913_),
    .A2(_07917_),
    .Y(_07918_),
    .B1(_07914_));
 sg13g2_nor2_1 _18015_ (.A(_07909_),
    .B(_07918_),
    .Y(_07919_));
 sg13g2_nor2_2 _18016_ (.A(_07910_),
    .B(_07919_),
    .Y(_07920_));
 sg13g2_and3_1 _18017_ (.X(_07921_),
    .A(_07874_),
    .B(_07887_),
    .C(_07920_));
 sg13g2_a21o_1 _18018_ (.A2(_07887_),
    .A1(_07874_),
    .B1(_07920_),
    .X(_07922_));
 sg13g2_nor2b_1 _18019_ (.A(net2726),
    .B_N(net2746),
    .Y(_07923_));
 sg13g2_xnor2_1 _18020_ (.Y(_07924_),
    .A(net2226),
    .B(net2328));
 sg13g2_xnor2_1 _18021_ (.Y(_07925_),
    .A(_07923_),
    .B(_07924_));
 sg13g2_nand2b_1 _18022_ (.Y(_07927_),
    .B(net2800),
    .A_N(net2655));
 sg13g2_xnor2_1 _18023_ (.Y(_07928_),
    .A(net2437),
    .B(net2372));
 sg13g2_xnor2_1 _18024_ (.Y(_07929_),
    .A(_07927_),
    .B(_07928_));
 sg13g2_nor2_1 _18025_ (.A(_07925_),
    .B(_07929_),
    .Y(_07930_));
 sg13g2_nand2_1 _18026_ (.Y(_07931_),
    .A(_07925_),
    .B(_07929_));
 sg13g2_xor2_1 _18027_ (.B(net2731),
    .A(net2567),
    .X(_07932_));
 sg13g2_xnor2_1 _18028_ (.Y(_07933_),
    .A(net2796),
    .B(net2237));
 sg13g2_nand2_2 _18029_ (.Y(_07934_),
    .A(_07932_),
    .B(_07933_));
 sg13g2_o21ai_1 _18030_ (.B1(_07931_),
    .Y(_07935_),
    .A1(_07930_),
    .A2(_07934_));
 sg13g2_nor2_1 _18031_ (.A(net2805),
    .B(net2276),
    .Y(_07936_));
 sg13g2_xnor2_1 _18032_ (.Y(_07938_),
    .A(net2239),
    .B(\net.in[13] ));
 sg13g2_nand2_1 _18033_ (.Y(_07939_),
    .A(_07936_),
    .B(_07938_));
 sg13g2_nor2_1 _18034_ (.A(net2222),
    .B(net2782),
    .Y(_07940_));
 sg13g2_nor2_1 _18035_ (.A(net2322),
    .B(net2614),
    .Y(_07941_));
 sg13g2_xnor2_1 _18036_ (.Y(_07942_),
    .A(_07940_),
    .B(_07941_));
 sg13g2_nand2b_1 _18037_ (.Y(_07943_),
    .B(_07942_),
    .A_N(_07939_));
 sg13g2_a21oi_1 _18038_ (.A1(_07936_),
    .A2(_07938_),
    .Y(_07944_),
    .B1(_07942_));
 sg13g2_xor2_1 _18039_ (.B(net2248),
    .A(net2289),
    .X(_07945_));
 sg13g2_xor2_1 _18040_ (.B(net2324),
    .A(net2415),
    .X(_07946_));
 sg13g2_nor2_1 _18041_ (.A(_07945_),
    .B(_07946_),
    .Y(_07947_));
 sg13g2_a21oi_2 _18042_ (.B1(_07944_),
    .Y(_07949_),
    .A2(_07947_),
    .A1(_07943_));
 sg13g2_inv_1 _18043_ (.Y(_07950_),
    .A(_07949_));
 sg13g2_nor2_1 _18044_ (.A(_07935_),
    .B(_07950_),
    .Y(_07951_));
 sg13g2_nor3_1 _18045_ (.A(net2214),
    .B(net2776),
    .C(_07856_),
    .Y(_07952_));
 sg13g2_nand2_1 _18046_ (.Y(_07953_),
    .A(net2415),
    .B(net2770));
 sg13g2_or2_1 _18047_ (.X(_07954_),
    .B(net2770),
    .A(net2415));
 sg13g2_nand2b_1 _18048_ (.Y(_07955_),
    .B(net2248),
    .A_N(net2368));
 sg13g2_nand3_1 _18049_ (.B(_07954_),
    .C(_07955_),
    .A(_07953_),
    .Y(_07956_));
 sg13g2_nor4_2 _18050_ (.A(net2214),
    .B(net2776),
    .C(_07856_),
    .Y(_07957_),
    .D(_07956_));
 sg13g2_nand2b_1 _18051_ (.Y(_07958_),
    .B(_07956_),
    .A_N(_07952_));
 sg13g2_o21ai_1 _18052_ (.B1(net2422),
    .Y(_07960_),
    .A1(_05627_),
    .A2(net2646));
 sg13g2_a21oi_1 _18053_ (.A1(_05627_),
    .A2(net2646),
    .Y(_07961_),
    .B1(net2597));
 sg13g2_nand2b_2 _18054_ (.Y(_07962_),
    .B(_07961_),
    .A_N(_07960_));
 sg13g2_o21ai_1 _18055_ (.B1(_07958_),
    .Y(_07963_),
    .A1(_07957_),
    .A2(_07962_));
 sg13g2_a21oi_1 _18056_ (.A1(_07935_),
    .A2(_07950_),
    .Y(_07964_),
    .B1(_07963_));
 sg13g2_nor2_2 _18057_ (.A(_07951_),
    .B(_07964_),
    .Y(_07965_));
 sg13g2_nand2b_1 _18058_ (.Y(_07966_),
    .B(_07965_),
    .A_N(_07921_));
 sg13g2_and2_2 _18059_ (.A(_07922_),
    .B(_07966_),
    .X(_07967_));
 sg13g2_nand3_1 _18060_ (.B(_07826_),
    .C(_07967_),
    .A(_07791_),
    .Y(_07968_));
 sg13g2_a21oi_1 _18061_ (.A1(_07791_),
    .A2(_07826_),
    .Y(_07969_),
    .B1(_07967_));
 sg13g2_nand2_2 _18062_ (.Y(_07971_),
    .A(_05220_),
    .B(_05957_));
 sg13g2_nand2_1 _18063_ (.Y(_07972_),
    .A(_05451_),
    .B(_05693_));
 sg13g2_nand2b_1 _18064_ (.Y(_07973_),
    .B(net2576),
    .A_N(net2673));
 sg13g2_xnor2_1 _18065_ (.Y(_07974_),
    .A(net2728),
    .B(net2562));
 sg13g2_a22oi_1 _18066_ (.Y(_07975_),
    .B1(_07973_),
    .B2(_07974_),
    .A2(_07972_),
    .A1(_07971_));
 sg13g2_nand4_1 _18067_ (.B(_07972_),
    .C(_07973_),
    .A(_07971_),
    .Y(_07976_),
    .D(_07974_));
 sg13g2_nor2b_1 _18068_ (.A(net2322),
    .B_N(net2686),
    .Y(_07977_));
 sg13g2_nor2_1 _18069_ (.A(net2558),
    .B(net2265),
    .Y(_07978_));
 sg13g2_xnor2_1 _18070_ (.Y(_07979_),
    .A(_07977_),
    .B(_07978_));
 sg13g2_o21ai_1 _18071_ (.B1(_07976_),
    .Y(_07980_),
    .A1(_07975_),
    .A2(_07979_));
 sg13g2_nor2_1 _18072_ (.A(net2695),
    .B(net2642),
    .Y(_07982_));
 sg13g2_xnor2_1 _18073_ (.Y(_07983_),
    .A(net2623),
    .B(_07982_));
 sg13g2_xnor2_1 _18074_ (.Y(_07984_),
    .A(net2467),
    .B(net2566));
 sg13g2_o21ai_1 _18075_ (.B1(_07984_),
    .Y(_07985_),
    .A1(net2292),
    .A2(net2235));
 sg13g2_nor2b_1 _18076_ (.A(_07983_),
    .B_N(_07985_),
    .Y(_07986_));
 sg13g2_nand2b_1 _18077_ (.Y(_07987_),
    .B(_07983_),
    .A_N(_07985_));
 sg13g2_or4_2 _18078_ (.A(net2492),
    .B(net2614),
    .C(net2503),
    .D(net2410),
    .X(_07988_));
 sg13g2_o21ai_1 _18079_ (.B1(_07987_),
    .Y(_07989_),
    .A1(_07986_),
    .A2(_07988_));
 sg13g2_nand2b_1 _18080_ (.Y(_07990_),
    .B(_07980_),
    .A_N(_07989_));
 sg13g2_nor2b_1 _18081_ (.A(_07980_),
    .B_N(_07989_),
    .Y(_07991_));
 sg13g2_nor2b_1 _18082_ (.A(net2509),
    .B_N(net2675),
    .Y(_07993_));
 sg13g2_nor2b_1 _18083_ (.A(net2675),
    .B_N(net2509),
    .Y(_07994_));
 sg13g2_nor2_1 _18084_ (.A(net2329),
    .B(net2235),
    .Y(_07995_));
 sg13g2_nor3_2 _18085_ (.A(_07993_),
    .B(_07994_),
    .C(_07995_),
    .Y(_07996_));
 sg13g2_nor2_1 _18086_ (.A(net2412),
    .B(net2814),
    .Y(_07997_));
 sg13g2_xnor2_1 _18087_ (.Y(_07998_),
    .A(_07755_),
    .B(_07997_));
 sg13g2_nor2_1 _18088_ (.A(_07996_),
    .B(_07998_),
    .Y(_07999_));
 sg13g2_nand2_1 _18089_ (.Y(_08000_),
    .A(_07996_),
    .B(_07998_));
 sg13g2_xor2_1 _18090_ (.B(net2786),
    .A(net2372),
    .X(_08001_));
 sg13g2_xor2_1 _18091_ (.B(net2682),
    .A(net2740),
    .X(_08002_));
 sg13g2_nand2_1 _18092_ (.Y(_08004_),
    .A(_08001_),
    .B(_08002_));
 sg13g2_o21ai_1 _18093_ (.B1(_08000_),
    .Y(_08005_),
    .A1(_07999_),
    .A2(_08004_));
 sg13g2_a21oi_2 _18094_ (.B1(_07991_),
    .Y(_08006_),
    .A2(_08005_),
    .A1(_07990_));
 sg13g2_nor2_1 _18095_ (.A(net2397),
    .B(net2597),
    .Y(_08007_));
 sg13g2_nor2_1 _18096_ (.A(net2244),
    .B(net2394),
    .Y(_08008_));
 sg13g2_nand2b_1 _18097_ (.Y(_08009_),
    .B(net2336),
    .A_N(net2781));
 sg13g2_xnor2_1 _18098_ (.Y(_08010_),
    .A(_08008_),
    .B(_08009_));
 sg13g2_nor2b_1 _18099_ (.A(_08007_),
    .B_N(_08010_),
    .Y(_08011_));
 sg13g2_nand2b_1 _18100_ (.Y(_08012_),
    .B(_08007_),
    .A_N(_08010_));
 sg13g2_nor2b_1 _18101_ (.A(net2348),
    .B_N(net2597),
    .Y(_08013_));
 sg13g2_nor3_1 _18102_ (.A(net2669),
    .B(net2503),
    .C(_08013_),
    .Y(_08015_));
 sg13g2_o21ai_1 _18103_ (.B1(_08015_),
    .Y(_08016_),
    .A1(_05121_),
    .A2(net2596));
 sg13g2_o21ai_1 _18104_ (.B1(_08012_),
    .Y(_08017_),
    .A1(_08011_),
    .A2(_08016_));
 sg13g2_nor2_1 _18105_ (.A(net2306),
    .B(net2731),
    .Y(_08018_));
 sg13g2_nor3_2 _18106_ (.A(net2187),
    .B(net2274),
    .C(_08018_),
    .Y(_08019_));
 sg13g2_nor2_1 _18107_ (.A(net2437),
    .B(net2740),
    .Y(_08020_));
 sg13g2_xnor2_1 _18108_ (.Y(_08021_),
    .A(net2805),
    .B(net2716));
 sg13g2_xnor2_1 _18109_ (.Y(_08022_),
    .A(_08020_),
    .B(_08021_));
 sg13g2_nor2b_1 _18110_ (.A(_08022_),
    .B_N(_08019_),
    .Y(_08023_));
 sg13g2_nand2b_1 _18111_ (.Y(_08024_),
    .B(_08022_),
    .A_N(_08019_));
 sg13g2_nand2_1 _18112_ (.Y(_08026_),
    .A(_05715_),
    .B(net2790));
 sg13g2_xnor2_1 _18113_ (.Y(_08027_),
    .A(_00023_),
    .B(_08026_));
 sg13g2_o21ai_1 _18114_ (.B1(_08024_),
    .Y(_08028_),
    .A1(_08023_),
    .A2(_08027_));
 sg13g2_or2_1 _18115_ (.X(_08029_),
    .B(_08028_),
    .A(_08017_));
 sg13g2_and2_1 _18116_ (.A(_08017_),
    .B(_08028_),
    .X(_08030_));
 sg13g2_or2_1 _18117_ (.X(_08031_),
    .B(net2738),
    .A(net2324));
 sg13g2_nand2_1 _18118_ (.Y(_08032_),
    .A(net2324),
    .B(net2738));
 sg13g2_nand3_1 _18119_ (.B(_08031_),
    .C(_08032_),
    .A(_02647_),
    .Y(_08033_));
 sg13g2_nor2_1 _18120_ (.A(net2388),
    .B(net2194),
    .Y(_08034_));
 sg13g2_nor2b_1 _18121_ (.A(net2656),
    .B_N(net2282),
    .Y(_08035_));
 sg13g2_xnor2_1 _18122_ (.Y(_08037_),
    .A(_08034_),
    .B(_08035_));
 sg13g2_nor2_1 _18123_ (.A(_08033_),
    .B(_08037_),
    .Y(_08038_));
 sg13g2_nor2_1 _18124_ (.A(net2530),
    .B(net2756),
    .Y(_08039_));
 sg13g2_a21oi_1 _18125_ (.A1(_08033_),
    .A2(_08037_),
    .Y(_08040_),
    .B1(_08039_));
 sg13g2_nor2_2 _18126_ (.A(_08038_),
    .B(_08040_),
    .Y(_08041_));
 sg13g2_a21oi_1 _18127_ (.A1(_08029_),
    .A2(_08041_),
    .Y(_08042_),
    .B1(_08030_));
 sg13g2_and2_1 _18128_ (.A(_08006_),
    .B(_08042_),
    .X(_08043_));
 sg13g2_nor2_1 _18129_ (.A(_08006_),
    .B(_08042_),
    .Y(_08044_));
 sg13g2_xnor2_1 _18130_ (.Y(_08045_),
    .A(net2190),
    .B(net2638));
 sg13g2_xnor2_1 _18131_ (.Y(_08046_),
    .A(net2728),
    .B(net2725));
 sg13g2_nand2_1 _18132_ (.Y(_08048_),
    .A(_08045_),
    .B(_08046_));
 sg13g2_o21ai_1 _18133_ (.B1(_08048_),
    .Y(_08049_),
    .A1(net2482),
    .A2(net2447));
 sg13g2_nand4_1 _18134_ (.B(_05407_),
    .C(_08045_),
    .A(net2184),
    .Y(_08050_),
    .D(_08046_));
 sg13g2_a22oi_1 _18135_ (.Y(_08051_),
    .B1(net2287),
    .B2(net2244),
    .A2(net2319),
    .A1(net2324));
 sg13g2_o21ai_1 _18136_ (.B1(_08051_),
    .Y(_08052_),
    .A1(net2324),
    .A2(net2319));
 sg13g2_nand2_1 _18137_ (.Y(_08053_),
    .A(_08049_),
    .B(_08052_));
 sg13g2_xnor2_1 _18138_ (.Y(_08054_),
    .A(net2437),
    .B(net2292));
 sg13g2_xnor2_1 _18139_ (.Y(_08055_),
    .A(net2677),
    .B(net2372));
 sg13g2_nor2_2 _18140_ (.A(_08054_),
    .B(_08055_),
    .Y(_08056_));
 sg13g2_or2_2 _18141_ (.X(_08057_),
    .B(\net.in[175] ),
    .A(net2239));
 sg13g2_nand2_1 _18142_ (.Y(_08059_),
    .A(_08056_),
    .B(_08057_));
 sg13g2_a21oi_2 _18143_ (.B1(net2805),
    .Y(_08060_),
    .A2(net2776),
    .A1(net2668));
 sg13g2_nor2b_2 _18144_ (.A(net2276),
    .B_N(_08060_),
    .Y(_08061_));
 sg13g2_nand2_1 _18145_ (.Y(_08062_),
    .A(_08059_),
    .B(_08061_));
 sg13g2_o21ai_1 _18146_ (.B1(_08062_),
    .Y(_08063_),
    .A1(_08056_),
    .A2(_08057_));
 sg13g2_nand3_1 _18147_ (.B(_08053_),
    .C(_08063_),
    .A(_08050_),
    .Y(_08064_));
 sg13g2_inv_1 _18148_ (.Y(_08065_),
    .A(_08064_));
 sg13g2_a21o_1 _18149_ (.A2(_08053_),
    .A1(_08050_),
    .B1(_08063_),
    .X(_08066_));
 sg13g2_xnor2_1 _18150_ (.Y(_08067_),
    .A(net2787),
    .B(net2668));
 sg13g2_nor3_2 _18151_ (.A(_05187_),
    .B(net2413),
    .C(_08067_),
    .Y(_08068_));
 sg13g2_xnor2_1 _18152_ (.Y(_08070_),
    .A(net2796),
    .B(net2690));
 sg13g2_xnor2_1 _18153_ (.Y(_08071_),
    .A(net2807),
    .B(_08070_));
 sg13g2_nand2b_1 _18154_ (.Y(_08072_),
    .B(_08071_),
    .A_N(_08068_));
 sg13g2_nor2b_1 _18155_ (.A(_08071_),
    .B_N(_08068_),
    .Y(_08073_));
 sg13g2_nor2_1 _18156_ (.A(net2740),
    .B(net2562),
    .Y(_08074_));
 sg13g2_xnor2_1 _18157_ (.Y(_08075_),
    .A(net2716),
    .B(_08074_));
 sg13g2_inv_1 _18158_ (.Y(_08076_),
    .A(_08075_));
 sg13g2_a21oi_1 _18159_ (.A1(_08072_),
    .A2(_08076_),
    .Y(_08077_),
    .B1(_08073_));
 sg13g2_o21ai_1 _18160_ (.B1(_08066_),
    .Y(_08078_),
    .A1(_08065_),
    .A2(_08077_));
 sg13g2_nor2_1 _18161_ (.A(_08044_),
    .B(_08078_),
    .Y(_08079_));
 sg13g2_nor2_2 _18162_ (.A(_08043_),
    .B(_08079_),
    .Y(_08081_));
 sg13g2_a21oi_2 _18163_ (.B1(_07969_),
    .Y(_08082_),
    .A2(_08081_),
    .A1(_07968_));
 sg13g2_inv_1 _18164_ (.Y(_08083_),
    .A(_08082_));
 sg13g2_nor2b_1 _18165_ (.A(_07930_),
    .B_N(_07931_),
    .Y(_08084_));
 sg13g2_xnor2_1 _18166_ (.Y(_08085_),
    .A(_07934_),
    .B(_08084_));
 sg13g2_xnor2_1 _18167_ (.Y(_08086_),
    .A(_07898_),
    .B(_07902_));
 sg13g2_xnor2_1 _18168_ (.Y(_08087_),
    .A(_07907_),
    .B(_08086_));
 sg13g2_xnor2_1 _18169_ (.Y(_08088_),
    .A(_07911_),
    .B(_07912_));
 sg13g2_xnor2_1 _18170_ (.Y(_08089_),
    .A(_07917_),
    .B(_08088_));
 sg13g2_nor2_1 _18171_ (.A(_08087_),
    .B(_08089_),
    .Y(_08090_));
 sg13g2_nand2_1 _18172_ (.Y(_08092_),
    .A(_08087_),
    .B(_08089_));
 sg13g2_xnor2_1 _18173_ (.Y(_08093_),
    .A(_08087_),
    .B(_08089_));
 sg13g2_xnor2_1 _18174_ (.Y(_08094_),
    .A(_08085_),
    .B(_08093_));
 sg13g2_xor2_1 _18175_ (.B(_07881_),
    .A(_07877_),
    .X(_08095_));
 sg13g2_xnor2_1 _18176_ (.Y(_08096_),
    .A(_07885_),
    .B(_08095_));
 sg13g2_xnor2_1 _18177_ (.Y(_08097_),
    .A(_07862_),
    .B(_07866_));
 sg13g2_xnor2_1 _18178_ (.Y(_08098_),
    .A(_07870_),
    .B(_08097_));
 sg13g2_xnor2_1 _18179_ (.Y(_08099_),
    .A(_08096_),
    .B(_08098_));
 sg13g2_and2_1 _18180_ (.A(_07891_),
    .B(_07892_),
    .X(_08100_));
 sg13g2_xnor2_1 _18181_ (.Y(_08101_),
    .A(_07895_),
    .B(_08100_));
 sg13g2_xnor2_1 _18182_ (.Y(_08103_),
    .A(_08099_),
    .B(_08101_));
 sg13g2_inv_1 _18183_ (.Y(_08104_),
    .A(_08103_));
 sg13g2_nor2_1 _18184_ (.A(_08094_),
    .B(_08104_),
    .Y(_08105_));
 sg13g2_xor2_1 _18185_ (.B(_07727_),
    .A(_07724_),
    .X(_08106_));
 sg13g2_xnor2_1 _18186_ (.Y(_08107_),
    .A(_07731_),
    .B(_08106_));
 sg13g2_xnor2_1 _18187_ (.Y(_08108_),
    .A(_07939_),
    .B(_07942_));
 sg13g2_xnor2_1 _18188_ (.Y(_08109_),
    .A(_07947_),
    .B(_08108_));
 sg13g2_or2_1 _18189_ (.X(_08110_),
    .B(_07962_),
    .A(_07958_));
 sg13g2_a22oi_1 _18190_ (.Y(_08111_),
    .B1(_07963_),
    .B2(_08110_),
    .A2(_07962_),
    .A1(_07957_));
 sg13g2_nor2b_1 _18191_ (.A(_08109_),
    .B_N(_08111_),
    .Y(_08112_));
 sg13g2_nand2b_1 _18192_ (.Y(_08114_),
    .B(_08109_),
    .A_N(_08111_));
 sg13g2_xnor2_1 _18193_ (.Y(_08115_),
    .A(_08109_),
    .B(_08111_));
 sg13g2_xor2_1 _18194_ (.B(_08115_),
    .A(_08107_),
    .X(_08116_));
 sg13g2_a21oi_1 _18195_ (.A1(_08094_),
    .A2(_08104_),
    .Y(_08117_),
    .B1(_08116_));
 sg13g2_nor2_1 _18196_ (.A(_08105_),
    .B(_08117_),
    .Y(_08118_));
 sg13g2_a21o_1 _18197_ (.A2(_07767_),
    .A1(_07765_),
    .B1(_07768_),
    .X(_08119_));
 sg13g2_o21ai_1 _18198_ (.B1(_08119_),
    .Y(_08120_),
    .A1(_07762_),
    .A2(_07765_));
 sg13g2_xor2_1 _18199_ (.B(_07752_),
    .A(_07748_),
    .X(_08121_));
 sg13g2_xnor2_1 _18200_ (.Y(_08122_),
    .A(_07757_),
    .B(_08121_));
 sg13g2_nand2_1 _18201_ (.Y(_08123_),
    .A(_07737_),
    .B(_07738_));
 sg13g2_xnor2_1 _18202_ (.Y(_08125_),
    .A(_07741_),
    .B(_08123_));
 sg13g2_nor2b_1 _18203_ (.A(_08125_),
    .B_N(_08122_),
    .Y(_08126_));
 sg13g2_nand2b_1 _18204_ (.Y(_08127_),
    .B(_08125_),
    .A_N(_08122_));
 sg13g2_xor2_1 _18205_ (.B(_08125_),
    .A(_08122_),
    .X(_08128_));
 sg13g2_xnor2_1 _18206_ (.Y(_08129_),
    .A(_08120_),
    .B(_08128_));
 sg13g2_nor2b_1 _18207_ (.A(_07784_),
    .B_N(_07785_),
    .Y(_08130_));
 sg13g2_xnor2_1 _18208_ (.Y(_08131_),
    .A(_07787_),
    .B(_08130_));
 sg13g2_nand2b_1 _18209_ (.Y(_08132_),
    .B(_07773_),
    .A_N(_07771_));
 sg13g2_xnor2_1 _18210_ (.Y(_08133_),
    .A(_07775_),
    .B(_08132_));
 sg13g2_nor2_1 _18211_ (.A(_08131_),
    .B(_08133_),
    .Y(_08134_));
 sg13g2_xnor2_1 _18212_ (.Y(_08136_),
    .A(_08131_),
    .B(_08133_));
 sg13g2_nand2_1 _18213_ (.Y(_08137_),
    .A(_07795_),
    .B(_07796_));
 sg13g2_xnor2_1 _18214_ (.Y(_08138_),
    .A(_07799_),
    .B(_08137_));
 sg13g2_xnor2_1 _18215_ (.Y(_08139_),
    .A(_08136_),
    .B(_08138_));
 sg13g2_nand2_1 _18216_ (.Y(_08140_),
    .A(_08129_),
    .B(_08139_));
 sg13g2_nor2_1 _18217_ (.A(_08129_),
    .B(_08139_),
    .Y(_08141_));
 sg13g2_xor2_1 _18218_ (.B(_07818_),
    .A(_07815_),
    .X(_08142_));
 sg13g2_xnor2_1 _18219_ (.Y(_08143_),
    .A(_07823_),
    .B(_08142_));
 sg13g2_xor2_1 _18220_ (.B(_07804_),
    .A(_07802_),
    .X(_08144_));
 sg13g2_xnor2_1 _18221_ (.Y(_08145_),
    .A(_07810_),
    .B(_08144_));
 sg13g2_nand2_1 _18222_ (.Y(_08147_),
    .A(_08143_),
    .B(_08145_));
 sg13g2_or2_1 _18223_ (.X(_08148_),
    .B(_08145_),
    .A(_08143_));
 sg13g2_nand2_1 _18224_ (.Y(_08149_),
    .A(_08147_),
    .B(_08148_));
 sg13g2_nand2b_1 _18225_ (.Y(_08150_),
    .B(_08024_),
    .A_N(_08023_));
 sg13g2_xnor2_1 _18226_ (.Y(_08151_),
    .A(_08027_),
    .B(_08150_));
 sg13g2_xor2_1 _18227_ (.B(_08151_),
    .A(_08149_),
    .X(_08152_));
 sg13g2_a21oi_1 _18228_ (.A1(_08140_),
    .A2(_08152_),
    .Y(_08153_),
    .B1(_08141_));
 sg13g2_nor2b_1 _18229_ (.A(_08118_),
    .B_N(_08153_),
    .Y(_08154_));
 sg13g2_nor3_1 _18230_ (.A(_08105_),
    .B(_08117_),
    .C(_08153_),
    .Y(_08155_));
 sg13g2_nand2b_1 _18231_ (.Y(_08156_),
    .B(_07976_),
    .A_N(_07975_));
 sg13g2_xnor2_1 _18232_ (.Y(_08158_),
    .A(_07979_),
    .B(_08156_));
 sg13g2_xnor2_1 _18233_ (.Y(_08159_),
    .A(_08007_),
    .B(_08010_));
 sg13g2_xnor2_1 _18234_ (.Y(_08160_),
    .A(_08016_),
    .B(_08159_));
 sg13g2_xnor2_1 _18235_ (.Y(_08161_),
    .A(_08033_),
    .B(_08037_));
 sg13g2_xnor2_1 _18236_ (.Y(_08162_),
    .A(_08039_),
    .B(_08161_));
 sg13g2_xnor2_1 _18237_ (.Y(_08163_),
    .A(_08160_),
    .B(_08162_));
 sg13g2_a21o_1 _18238_ (.A2(_08162_),
    .A1(_08160_),
    .B1(_08158_),
    .X(_08164_));
 sg13g2_o21ai_1 _18239_ (.B1(_08164_),
    .Y(_08165_),
    .A1(_08160_),
    .A2(_08162_));
 sg13g2_xnor2_1 _18240_ (.Y(_08166_),
    .A(_08158_),
    .B(_08163_));
 sg13g2_nand2_1 _18241_ (.Y(_08167_),
    .A(_08049_),
    .B(_08050_));
 sg13g2_xor2_1 _18242_ (.B(_08167_),
    .A(_08052_),
    .X(_08169_));
 sg13g2_xor2_1 _18243_ (.B(_07985_),
    .A(_07983_),
    .X(_08170_));
 sg13g2_xnor2_1 _18244_ (.Y(_08171_),
    .A(_07988_),
    .B(_08170_));
 sg13g2_xnor2_1 _18245_ (.Y(_08172_),
    .A(_07996_),
    .B(_07998_));
 sg13g2_xnor2_1 _18246_ (.Y(_08173_),
    .A(_08004_),
    .B(_08172_));
 sg13g2_xor2_1 _18247_ (.B(_08173_),
    .A(_08171_),
    .X(_08174_));
 sg13g2_xnor2_1 _18248_ (.Y(_08175_),
    .A(_08169_),
    .B(_08174_));
 sg13g2_nor2_1 _18249_ (.A(_08166_),
    .B(_08175_),
    .Y(_08176_));
 sg13g2_nand2_1 _18250_ (.Y(_08177_),
    .A(_08166_),
    .B(_08175_));
 sg13g2_and3_2 _18251_ (.X(_08178_),
    .A(_05495_),
    .B(_05858_),
    .C(_00022_));
 sg13g2_xor2_1 _18252_ (.B(net2748),
    .A(net2668),
    .X(_08180_));
 sg13g2_xnor2_1 _18253_ (.Y(_08181_),
    .A(net2194),
    .B(net2282));
 sg13g2_nor3_1 _18254_ (.A(_02558_),
    .B(_08180_),
    .C(_08181_),
    .Y(_08182_));
 sg13g2_o21ai_1 _18255_ (.B1(_08181_),
    .Y(_08183_),
    .A1(_02558_),
    .A2(_08180_));
 sg13g2_nor2b_1 _18256_ (.A(_08182_),
    .B_N(_08183_),
    .Y(_08184_));
 sg13g2_xnor2_1 _18257_ (.Y(_08185_),
    .A(_08178_),
    .B(_08184_));
 sg13g2_xnor2_1 _18258_ (.Y(_08186_),
    .A(_08068_),
    .B(_08071_));
 sg13g2_xnor2_1 _18259_ (.Y(_08187_),
    .A(_08075_),
    .B(_08186_));
 sg13g2_xor2_1 _18260_ (.B(_08057_),
    .A(_08056_),
    .X(_08188_));
 sg13g2_xnor2_1 _18261_ (.Y(_08189_),
    .A(_08061_),
    .B(_08188_));
 sg13g2_nand2_1 _18262_ (.Y(_08191_),
    .A(_08187_),
    .B(_08189_));
 sg13g2_or2_1 _18263_ (.X(_08192_),
    .B(_08191_),
    .A(_08185_));
 sg13g2_nor2_1 _18264_ (.A(_08187_),
    .B(_08189_),
    .Y(_08193_));
 sg13g2_a21oi_1 _18265_ (.A1(_08185_),
    .A2(_08191_),
    .Y(_08194_),
    .B1(_08193_));
 sg13g2_and2_1 _18266_ (.A(_08185_),
    .B(_08193_),
    .X(_08195_));
 sg13g2_o21ai_1 _18267_ (.B1(_08192_),
    .Y(_08196_),
    .A1(_08194_),
    .A2(_08195_));
 sg13g2_inv_1 _18268_ (.Y(_08197_),
    .A(_08196_));
 sg13g2_o21ai_1 _18269_ (.B1(_08177_),
    .Y(_08198_),
    .A1(_08176_),
    .A2(_08197_));
 sg13g2_nor2_1 _18270_ (.A(_08155_),
    .B(_08198_),
    .Y(_08199_));
 sg13g2_nor2_1 _18271_ (.A(_08154_),
    .B(_08199_),
    .Y(_08200_));
 sg13g2_xor2_1 _18272_ (.B(net2766),
    .A(net2370),
    .X(_08202_));
 sg13g2_nor3_2 _18273_ (.A(net2505),
    .B(net2596),
    .C(_08202_),
    .Y(_08203_));
 sg13g2_nor2_1 _18274_ (.A(net2725),
    .B(net2552),
    .Y(_08204_));
 sg13g2_xnor2_1 _18275_ (.Y(_08205_),
    .A(_00024_),
    .B(_08204_));
 sg13g2_nor2_1 _18276_ (.A(net2800),
    .B(net2220),
    .Y(_08206_));
 sg13g2_xnor2_1 _18277_ (.Y(_08207_),
    .A(net2322),
    .B(net2728));
 sg13g2_xnor2_1 _18278_ (.Y(_08208_),
    .A(_08206_),
    .B(_08207_));
 sg13g2_nor2_1 _18279_ (.A(_08205_),
    .B(_08208_),
    .Y(_08209_));
 sg13g2_xnor2_1 _18280_ (.Y(_08210_),
    .A(_08205_),
    .B(_08208_));
 sg13g2_xnor2_1 _18281_ (.Y(_08211_),
    .A(_08203_),
    .B(_08210_));
 sg13g2_nor2_1 _18282_ (.A(net2460),
    .B(net2743),
    .Y(_08213_));
 sg13g2_o21ai_1 _18283_ (.B1(_08213_),
    .Y(_08214_),
    .A1(net2571),
    .A2(net2269));
 sg13g2_xnor2_1 _18284_ (.Y(_08215_),
    .A(net2558),
    .B(net2746));
 sg13g2_nand3_1 _18285_ (.B(_05968_),
    .C(_08215_),
    .A(net2570),
    .Y(_08216_));
 sg13g2_xnor2_1 _18286_ (.Y(_08217_),
    .A(net2505),
    .B(net2668));
 sg13g2_nand2b_1 _18287_ (.Y(_08218_),
    .B(_08217_),
    .A_N(_08216_));
 sg13g2_nor2b_1 _18288_ (.A(_08217_),
    .B_N(_08216_),
    .Y(_08219_));
 sg13g2_xnor2_1 _18289_ (.Y(_08220_),
    .A(_08216_),
    .B(_08217_));
 sg13g2_o21ai_1 _18290_ (.B1(_08218_),
    .Y(_08221_),
    .A1(_08214_),
    .A2(_08219_));
 sg13g2_xnor2_1 _18291_ (.Y(_08222_),
    .A(_08214_),
    .B(_08220_));
 sg13g2_xor2_1 _18292_ (.B(_08222_),
    .A(_08211_),
    .X(_08224_));
 sg13g2_xor2_1 _18293_ (.B(net2418),
    .A(net2525),
    .X(_08225_));
 sg13g2_nand2b_1 _18294_ (.Y(_08226_),
    .B(net2252),
    .A_N(net2270));
 sg13g2_nor2_1 _18295_ (.A(net2437),
    .B(net2397),
    .Y(_08227_));
 sg13g2_a22oi_1 _18296_ (.Y(_08228_),
    .B1(_08226_),
    .B2(_08227_),
    .A2(_08225_),
    .A1(_06584_));
 sg13g2_nand4_1 _18297_ (.B(_08225_),
    .C(_08226_),
    .A(_06584_),
    .Y(_08229_),
    .D(_08227_));
 sg13g2_nand2b_1 _18298_ (.Y(_08230_),
    .B(_08229_),
    .A_N(_08228_));
 sg13g2_nand2_1 _18299_ (.Y(_08231_),
    .A(net2194),
    .B(net2702));
 sg13g2_o21ai_1 _18300_ (.B1(_08231_),
    .Y(_08232_),
    .A1(net2702),
    .A2(_08181_));
 sg13g2_xnor2_1 _18301_ (.Y(_08233_),
    .A(_08230_),
    .B(_08232_));
 sg13g2_xnor2_1 _18302_ (.Y(_08235_),
    .A(_08224_),
    .B(_08233_));
 sg13g2_xor2_1 _18303_ (.B(net2199),
    .A(net2269),
    .X(_08236_));
 sg13g2_nor2b_1 _18304_ (.A(net2397),
    .B_N(net2505),
    .Y(_08237_));
 sg13g2_nor2b_1 _18305_ (.A(net2505),
    .B_N(net2397),
    .Y(_08238_));
 sg13g2_nor3_1 _18306_ (.A(_07828_),
    .B(_08237_),
    .C(_08238_),
    .Y(_08239_));
 sg13g2_nand3_1 _18307_ (.B(net2289),
    .C(net2463),
    .A(_05066_),
    .Y(_08240_));
 sg13g2_nor4_1 _18308_ (.A(_07828_),
    .B(_08237_),
    .C(_08238_),
    .D(_08240_),
    .Y(_08241_));
 sg13g2_nand2b_1 _18309_ (.Y(_08242_),
    .B(_08240_),
    .A_N(_08239_));
 sg13g2_xnor2_1 _18310_ (.Y(_08243_),
    .A(_08239_),
    .B(_08240_));
 sg13g2_o21ai_1 _18311_ (.B1(_08242_),
    .Y(_08244_),
    .A1(_08236_),
    .A2(_08241_));
 sg13g2_xnor2_1 _18312_ (.Y(_08246_),
    .A(_08236_),
    .B(_08243_));
 sg13g2_xnor2_1 _18313_ (.Y(_08247_),
    .A(net2434),
    .B(net2376));
 sg13g2_nor2b_1 _18314_ (.A(net2558),
    .B_N(net2673),
    .Y(_08248_));
 sg13g2_nor2b_1 _18315_ (.A(net2673),
    .B_N(net2558),
    .Y(_08249_));
 sg13g2_nor2_1 _18316_ (.A(net2332),
    .B(net2235),
    .Y(_08250_));
 sg13g2_nor3_2 _18317_ (.A(_08248_),
    .B(_08249_),
    .C(_08250_),
    .Y(_08251_));
 sg13g2_nor2b_1 _18318_ (.A(_08251_),
    .B_N(_08060_),
    .Y(_08252_));
 sg13g2_nand2b_1 _18319_ (.Y(_08253_),
    .B(_08251_),
    .A_N(_08060_));
 sg13g2_xor2_1 _18320_ (.B(_08251_),
    .A(_08060_),
    .X(_08254_));
 sg13g2_xnor2_1 _18321_ (.Y(_08255_),
    .A(_08247_),
    .B(_08254_));
 sg13g2_nor2_1 _18322_ (.A(_08246_),
    .B(_08255_),
    .Y(_08257_));
 sg13g2_xor2_1 _18323_ (.B(_08255_),
    .A(_08246_),
    .X(_08258_));
 sg13g2_nor2_1 _18324_ (.A(net2769),
    .B(net2177),
    .Y(_08259_));
 sg13g2_xnor2_1 _18325_ (.Y(_08260_),
    .A(net2269),
    .B(_08259_));
 sg13g2_xnor2_1 _18326_ (.Y(_08261_),
    .A(net2800),
    .B(net2534));
 sg13g2_xnor2_1 _18327_ (.Y(_08262_),
    .A(net2686),
    .B(net2792));
 sg13g2_xor2_1 _18328_ (.B(net2328),
    .A(net2389),
    .X(_08263_));
 sg13g2_nand3_1 _18329_ (.B(_08262_),
    .C(_08263_),
    .A(_08261_),
    .Y(_08264_));
 sg13g2_a21o_1 _18330_ (.A2(_08262_),
    .A1(_08261_),
    .B1(_08263_),
    .X(_08265_));
 sg13g2_nand2_1 _18331_ (.Y(_08266_),
    .A(_08264_),
    .B(_08265_));
 sg13g2_xor2_1 _18332_ (.B(_08266_),
    .A(_08260_),
    .X(_08268_));
 sg13g2_xnor2_1 _18333_ (.Y(_08269_),
    .A(_08258_),
    .B(_08268_));
 sg13g2_nand2_1 _18334_ (.Y(_08270_),
    .A(_08235_),
    .B(_08269_));
 sg13g2_or2_1 _18335_ (.X(_08271_),
    .B(_08269_),
    .A(_08235_));
 sg13g2_nand2_1 _18336_ (.Y(_08272_),
    .A(net2422),
    .B(_08215_));
 sg13g2_nor2_2 _18337_ (.A(net2530),
    .B(_08272_),
    .Y(_08273_));
 sg13g2_xnor2_1 _18338_ (.Y(_08274_),
    .A(net2652),
    .B(net2287));
 sg13g2_xnor2_1 _18339_ (.Y(_08275_),
    .A(net2299),
    .B(_08274_));
 sg13g2_nor2_1 _18340_ (.A(net2412),
    .B(_07763_),
    .Y(_08276_));
 sg13g2_and2_1 _18341_ (.A(net2412),
    .B(net2816),
    .X(_08277_));
 sg13g2_nor3_1 _18342_ (.A(_08275_),
    .B(_08276_),
    .C(_08277_),
    .Y(_08279_));
 sg13g2_o21ai_1 _18343_ (.B1(_08275_),
    .Y(_08280_),
    .A1(_08276_),
    .A2(_08277_));
 sg13g2_nand2b_1 _18344_ (.Y(_08281_),
    .B(_08280_),
    .A_N(_08279_));
 sg13g2_xor2_1 _18345_ (.B(_08281_),
    .A(_08273_),
    .X(_08282_));
 sg13g2_nor2_1 _18346_ (.A(net2367),
    .B(net2746),
    .Y(_08283_));
 sg13g2_xnor2_1 _18347_ (.Y(_08284_),
    .A(net2769),
    .B(net2309));
 sg13g2_xnor2_1 _18348_ (.Y(_08285_),
    .A(_08283_),
    .B(_08284_));
 sg13g2_nor2_1 _18349_ (.A(net2769),
    .B(net2618),
    .Y(_08286_));
 sg13g2_nor2_1 _18350_ (.A(net2725),
    .B(net2457),
    .Y(_08287_));
 sg13g2_xor2_1 _18351_ (.B(_08287_),
    .A(_08286_),
    .X(_08288_));
 sg13g2_nor2_1 _18352_ (.A(_08285_),
    .B(_08288_),
    .Y(_08290_));
 sg13g2_xor2_1 _18353_ (.B(_08288_),
    .A(_08285_),
    .X(_08291_));
 sg13g2_xor2_1 _18354_ (.B(net2766),
    .A(net2677),
    .X(_08292_));
 sg13g2_xnor2_1 _18355_ (.Y(_08293_),
    .A(_07875_),
    .B(_08292_));
 sg13g2_xnor2_1 _18356_ (.Y(_08294_),
    .A(_08291_),
    .B(_08293_));
 sg13g2_nand2_1 _18357_ (.Y(_08295_),
    .A(_08282_),
    .B(_08294_));
 sg13g2_or2_1 _18358_ (.X(_08296_),
    .B(_08294_),
    .A(_08282_));
 sg13g2_nand2_1 _18359_ (.Y(_08297_),
    .A(_08295_),
    .B(_08296_));
 sg13g2_nand2_1 _18360_ (.Y(_08298_),
    .A(net2380),
    .B(_07984_));
 sg13g2_nor2_1 _18361_ (.A(net2413),
    .B(net2738),
    .Y(_08299_));
 sg13g2_nand2_1 _18362_ (.Y(_08301_),
    .A(_05352_),
    .B(_05946_));
 sg13g2_xnor2_1 _18363_ (.Y(_08302_),
    .A(net2477),
    .B(net2252));
 sg13g2_o21ai_1 _18364_ (.B1(_08302_),
    .Y(_08303_),
    .A1(_00874_),
    .A2(_08301_));
 sg13g2_or3_1 _18365_ (.A(_00874_),
    .B(_08301_),
    .C(_08302_),
    .X(_08304_));
 sg13g2_nand2_1 _18366_ (.Y(_08305_),
    .A(_08303_),
    .B(_08304_));
 sg13g2_xor2_1 _18367_ (.B(_08305_),
    .A(_08298_),
    .X(_08306_));
 sg13g2_xnor2_1 _18368_ (.Y(_08307_),
    .A(_08297_),
    .B(_08306_));
 sg13g2_nand2_1 _18369_ (.Y(_08308_),
    .A(_08270_),
    .B(_08307_));
 sg13g2_xnor2_1 _18370_ (.Y(_08309_),
    .A(net2462),
    .B(net2667));
 sg13g2_xnor2_1 _18371_ (.Y(_08310_),
    .A(net2615),
    .B(net2746));
 sg13g2_nand3_1 _18372_ (.B(_08309_),
    .C(_08310_),
    .A(_06573_),
    .Y(_08312_));
 sg13g2_a21o_1 _18373_ (.A2(_08309_),
    .A1(_06573_),
    .B1(_08310_),
    .X(_08313_));
 sg13g2_nand2_1 _18374_ (.Y(_08314_),
    .A(_08312_),
    .B(_08313_));
 sg13g2_xnor2_1 _18375_ (.Y(_08315_),
    .A(net2509),
    .B(net2714));
 sg13g2_xnor2_1 _18376_ (.Y(_08316_),
    .A(_08314_),
    .B(_08315_));
 sg13g2_xnor2_1 _18377_ (.Y(_08317_),
    .A(net2231),
    .B(net2638));
 sg13g2_nor2_2 _18378_ (.A(_00886_),
    .B(_08317_),
    .Y(_08318_));
 sg13g2_xor2_1 _18379_ (.B(net2269),
    .A(net2517),
    .X(_08319_));
 sg13g2_xor2_1 _18380_ (.B(net2677),
    .A(net2694),
    .X(_08320_));
 sg13g2_nand2_2 _18381_ (.Y(_08321_),
    .A(_08319_),
    .B(_08320_));
 sg13g2_nand2_2 _18382_ (.Y(_08323_),
    .A(_00011_),
    .B(_07763_));
 sg13g2_nand2b_1 _18383_ (.Y(_08324_),
    .B(_08321_),
    .A_N(_08323_));
 sg13g2_nor2b_1 _18384_ (.A(_08321_),
    .B_N(_08323_),
    .Y(_08325_));
 sg13g2_xor2_1 _18385_ (.B(_08323_),
    .A(_08321_),
    .X(_08326_));
 sg13g2_xnor2_1 _18386_ (.Y(_08327_),
    .A(_08318_),
    .B(_08326_));
 sg13g2_nor2_1 _18387_ (.A(_08316_),
    .B(_08327_),
    .Y(_08328_));
 sg13g2_nand2_1 _18388_ (.Y(_08329_),
    .A(_08316_),
    .B(_08327_));
 sg13g2_xnor2_1 _18389_ (.Y(_08330_),
    .A(_08316_),
    .B(_08327_));
 sg13g2_xnor2_1 _18390_ (.Y(_08331_),
    .A(net2392),
    .B(net2285));
 sg13g2_nor2b_1 _18391_ (.A(net2743),
    .B_N(net2516),
    .Y(_08332_));
 sg13g2_xnor2_1 _18392_ (.Y(_08334_),
    .A(net2629),
    .B(net2597));
 sg13g2_xnor2_1 _18393_ (.Y(_08335_),
    .A(_08332_),
    .B(_08334_));
 sg13g2_nand2_1 _18394_ (.Y(_08336_),
    .A(_08331_),
    .B(_08335_));
 sg13g2_nor2_1 _18395_ (.A(_08331_),
    .B(_08335_),
    .Y(_08337_));
 sg13g2_xor2_1 _18396_ (.B(_08335_),
    .A(_08331_),
    .X(_08338_));
 sg13g2_nor2_1 _18397_ (.A(net2800),
    .B(net2748),
    .Y(_08339_));
 sg13g2_nor2_1 _18398_ (.A(net2505),
    .B(net2177),
    .Y(_08340_));
 sg13g2_xnor2_1 _18399_ (.Y(_08341_),
    .A(_08339_),
    .B(_08340_));
 sg13g2_xnor2_1 _18400_ (.Y(_08342_),
    .A(_08338_),
    .B(_08341_));
 sg13g2_xnor2_1 _18401_ (.Y(_08343_),
    .A(_08330_),
    .B(_08342_));
 sg13g2_xnor2_1 _18402_ (.Y(_08345_),
    .A(_07840_),
    .B(_07846_));
 sg13g2_xnor2_1 _18403_ (.Y(_08346_),
    .A(_07859_),
    .B(_08345_));
 sg13g2_nand2_1 _18404_ (.Y(_08347_),
    .A(_08343_),
    .B(_08346_));
 sg13g2_or2_1 _18405_ (.X(_08348_),
    .B(_08346_),
    .A(_08343_));
 sg13g2_o21ai_1 _18406_ (.B1(_08299_),
    .Y(_08349_),
    .A1(net2572),
    .A2(_05693_));
 sg13g2_nand2b_1 _18407_ (.Y(_08350_),
    .B(_08347_),
    .A_N(_08349_));
 sg13g2_and4_1 _18408_ (.A(_08271_),
    .B(_08308_),
    .C(_08348_),
    .D(_08350_),
    .X(_08351_));
 sg13g2_a22oi_1 _18409_ (.Y(_08352_),
    .B1(_08348_),
    .B2(_08350_),
    .A2(_08308_),
    .A1(_08271_));
 sg13g2_a21o_1 _18410_ (.A2(_08098_),
    .A1(_08096_),
    .B1(_08101_),
    .X(_08353_));
 sg13g2_o21ai_1 _18411_ (.B1(_08353_),
    .Y(_08354_),
    .A1(_08096_),
    .A2(_08098_));
 sg13g2_nor2_1 _18412_ (.A(_08352_),
    .B(_08354_),
    .Y(_08356_));
 sg13g2_or2_2 _18413_ (.X(_08357_),
    .B(_08356_),
    .A(_08351_));
 sg13g2_o21ai_1 _18414_ (.B1(_08357_),
    .Y(_08358_),
    .A1(_08154_),
    .A2(_08199_));
 sg13g2_nor3_1 _18415_ (.A(_08154_),
    .B(_08199_),
    .C(_08357_),
    .Y(_08359_));
 sg13g2_a21oi_1 _18416_ (.A1(_08085_),
    .A2(_08092_),
    .Y(_08360_),
    .B1(_08090_));
 sg13g2_a21oi_1 _18417_ (.A1(_08107_),
    .A2(_08114_),
    .Y(_08361_),
    .B1(_08112_));
 sg13g2_nand2_1 _18418_ (.Y(_08362_),
    .A(_08360_),
    .B(_08361_));
 sg13g2_nor2_1 _18419_ (.A(_08360_),
    .B(_08361_),
    .Y(_08363_));
 sg13g2_a21oi_2 _18420_ (.B1(_08126_),
    .Y(_08364_),
    .A2(_08127_),
    .A1(_08120_));
 sg13g2_a21oi_2 _18421_ (.B1(_08363_),
    .Y(_08365_),
    .A2(_08364_),
    .A1(_08362_));
 sg13g2_inv_1 _18422_ (.Y(_08367_),
    .A(_08365_));
 sg13g2_a21oi_2 _18423_ (.B1(_08359_),
    .Y(_08368_),
    .A2(_08367_),
    .A1(_08358_));
 sg13g2_nand2b_1 _18424_ (.Y(_08369_),
    .B(_08232_),
    .A_N(_08228_));
 sg13g2_nand2b_1 _18425_ (.Y(_08370_),
    .B(_08273_),
    .A_N(_08279_));
 sg13g2_a22oi_1 _18426_ (.Y(_08371_),
    .B1(_08370_),
    .B2(_08280_),
    .A2(_08369_),
    .A1(_08229_));
 sg13g2_nand4_1 _18427_ (.B(_08280_),
    .C(_08369_),
    .A(_08229_),
    .Y(_08372_),
    .D(_08370_));
 sg13g2_nor2b_1 _18428_ (.A(_08371_),
    .B_N(_08372_),
    .Y(_08373_));
 sg13g2_a21oi_1 _18429_ (.A1(_08285_),
    .A2(_08288_),
    .Y(_08374_),
    .B1(_08293_));
 sg13g2_nor2_1 _18430_ (.A(_08290_),
    .B(_08374_),
    .Y(_08375_));
 sg13g2_xnor2_1 _18431_ (.Y(_08376_),
    .A(_08373_),
    .B(_08375_));
 sg13g2_nand2_1 _18432_ (.Y(_08378_),
    .A(_08313_),
    .B(_08315_));
 sg13g2_and2_1 _18433_ (.A(_08312_),
    .B(_08378_),
    .X(_08379_));
 sg13g2_nand2b_1 _18434_ (.Y(_08380_),
    .B(_08303_),
    .A_N(_08298_));
 sg13g2_a21o_1 _18435_ (.A2(_08380_),
    .A1(_08304_),
    .B1(_08379_),
    .X(_08381_));
 sg13g2_nand3_1 _18436_ (.B(_08379_),
    .C(_08380_),
    .A(_08304_),
    .Y(_08382_));
 sg13g2_nand2_1 _18437_ (.Y(_08383_),
    .A(_08381_),
    .B(_08382_));
 sg13g2_a21oi_1 _18438_ (.A1(_08318_),
    .A2(_08324_),
    .Y(_08384_),
    .B1(_08325_));
 sg13g2_xnor2_1 _18439_ (.Y(_08385_),
    .A(_08383_),
    .B(_08384_));
 sg13g2_nand2_1 _18440_ (.Y(_08386_),
    .A(_08376_),
    .B(_08385_));
 sg13g2_nor2_1 _18441_ (.A(_08376_),
    .B(_08385_),
    .Y(_08387_));
 sg13g2_a21oi_1 _18442_ (.A1(_08336_),
    .A2(_08341_),
    .Y(_08389_),
    .B1(_08337_));
 sg13g2_a21oi_1 _18443_ (.A1(_07829_),
    .A2(_07836_),
    .Y(_08390_),
    .B1(_07837_));
 sg13g2_and2_1 _18444_ (.A(_08389_),
    .B(_08390_),
    .X(_08391_));
 sg13g2_nor2_1 _18445_ (.A(_08389_),
    .B(_08390_),
    .Y(_08392_));
 sg13g2_nor2_1 _18446_ (.A(_08391_),
    .B(_08392_),
    .Y(_08393_));
 sg13g2_a21oi_1 _18447_ (.A1(_07841_),
    .A2(_07842_),
    .Y(_08394_),
    .B1(_07845_));
 sg13g2_nor2_2 _18448_ (.A(_07843_),
    .B(_08394_),
    .Y(_08395_));
 sg13g2_xnor2_1 _18449_ (.Y(_08396_),
    .A(_08393_),
    .B(_08395_));
 sg13g2_a21oi_2 _18450_ (.B1(_08387_),
    .Y(_08397_),
    .A2(_08396_),
    .A1(_08386_));
 sg13g2_nand2_1 _18451_ (.Y(_08398_),
    .A(_08064_),
    .B(_08066_));
 sg13g2_xor2_1 _18452_ (.B(_08398_),
    .A(_08077_),
    .X(_08400_));
 sg13g2_a21oi_2 _18453_ (.B1(_08182_),
    .Y(_08401_),
    .A2(_08183_),
    .A1(_08178_));
 sg13g2_nand2_1 _18454_ (.Y(_08402_),
    .A(_08244_),
    .B(_08401_));
 sg13g2_nor2_1 _18455_ (.A(_08244_),
    .B(_08401_),
    .Y(_08403_));
 sg13g2_xnor2_1 _18456_ (.Y(_08404_),
    .A(_08244_),
    .B(_08401_));
 sg13g2_o21ai_1 _18457_ (.B1(_08253_),
    .Y(_08405_),
    .A1(_08247_),
    .A2(_08252_));
 sg13g2_xnor2_1 _18458_ (.Y(_08406_),
    .A(_08404_),
    .B(_08405_));
 sg13g2_nand2_1 _18459_ (.Y(_08407_),
    .A(_08400_),
    .B(_08406_));
 sg13g2_a21oi_1 _18460_ (.A1(_08205_),
    .A2(_08208_),
    .Y(_08408_),
    .B1(_08203_));
 sg13g2_nor2_1 _18461_ (.A(_08209_),
    .B(_08408_),
    .Y(_08409_));
 sg13g2_nand2_1 _18462_ (.Y(_08411_),
    .A(_08260_),
    .B(_08264_));
 sg13g2_and2_1 _18463_ (.A(_08265_),
    .B(_08411_),
    .X(_08412_));
 sg13g2_xor2_1 _18464_ (.B(_08412_),
    .A(_08409_),
    .X(_08413_));
 sg13g2_xnor2_1 _18465_ (.Y(_08414_),
    .A(_08221_),
    .B(_08413_));
 sg13g2_nand2_1 _18466_ (.Y(_08415_),
    .A(_08407_),
    .B(_08414_));
 sg13g2_o21ai_1 _18467_ (.B1(_08415_),
    .Y(_08416_),
    .A1(_08400_),
    .A2(_08406_));
 sg13g2_nand2_1 _18468_ (.Y(_08417_),
    .A(_08397_),
    .B(_08416_));
 sg13g2_nor2_1 _18469_ (.A(_08397_),
    .B(_08416_),
    .Y(_08418_));
 sg13g2_nand2_1 _18470_ (.Y(_08419_),
    .A(_08347_),
    .B(_08348_));
 sg13g2_xor2_1 _18471_ (.B(_08419_),
    .A(_08349_),
    .X(_08420_));
 sg13g2_nand2_1 _18472_ (.Y(_08422_),
    .A(_08270_),
    .B(_08271_));
 sg13g2_xor2_1 _18473_ (.B(_08422_),
    .A(_08307_),
    .X(_08423_));
 sg13g2_nor2b_1 _18474_ (.A(_08423_),
    .B_N(_08420_),
    .Y(_08424_));
 sg13g2_xnor2_1 _18475_ (.Y(_08425_),
    .A(_08420_),
    .B(_08423_));
 sg13g2_xor2_1 _18476_ (.B(_08103_),
    .A(_08094_),
    .X(_08426_));
 sg13g2_xnor2_1 _18477_ (.Y(_08427_),
    .A(_08116_),
    .B(_08426_));
 sg13g2_xor2_1 _18478_ (.B(_08139_),
    .A(_08129_),
    .X(_08428_));
 sg13g2_xnor2_1 _18479_ (.Y(_08429_),
    .A(_08152_),
    .B(_08428_));
 sg13g2_nand2b_1 _18480_ (.Y(_08430_),
    .B(_08429_),
    .A_N(_08427_));
 sg13g2_nor2b_1 _18481_ (.A(_08429_),
    .B_N(_08427_),
    .Y(_08431_));
 sg13g2_xor2_1 _18482_ (.B(_08429_),
    .A(_08427_),
    .X(_08433_));
 sg13g2_nand2b_1 _18483_ (.Y(_08434_),
    .B(_08177_),
    .A_N(_08176_));
 sg13g2_xnor2_1 _18484_ (.Y(_08435_),
    .A(_08196_),
    .B(_08434_));
 sg13g2_xnor2_1 _18485_ (.Y(_08436_),
    .A(_08433_),
    .B(_08435_));
 sg13g2_a21oi_1 _18486_ (.A1(_08425_),
    .A2(_08436_),
    .Y(_08437_),
    .B1(_08424_));
 sg13g2_a21oi_1 _18487_ (.A1(_08430_),
    .A2(_08435_),
    .Y(_08438_),
    .B1(_08431_));
 sg13g2_nor2_1 _18488_ (.A(_08437_),
    .B(_08438_),
    .Y(_08439_));
 sg13g2_a21oi_1 _18489_ (.A1(_08417_),
    .A2(_08439_),
    .Y(_08440_),
    .B1(_08418_));
 sg13g2_nand2_1 _18490_ (.Y(_08441_),
    .A(_08368_),
    .B(_08440_));
 sg13g2_or2_1 _18491_ (.X(_08442_),
    .B(_08440_),
    .A(_08368_));
 sg13g2_inv_1 _18492_ (.Y(_08444_),
    .A(_08442_));
 sg13g2_nor2_1 _18493_ (.A(_08134_),
    .B(_08138_),
    .Y(_08445_));
 sg13g2_a21oi_1 _18494_ (.A1(_08131_),
    .A2(_08133_),
    .Y(_08446_),
    .B1(_08445_));
 sg13g2_nand2b_1 _18495_ (.Y(_08447_),
    .B(_08147_),
    .A_N(_08151_));
 sg13g2_nand3_1 _18496_ (.B(_08446_),
    .C(_08447_),
    .A(_08148_),
    .Y(_08448_));
 sg13g2_a21o_1 _18497_ (.A2(_08447_),
    .A1(_08148_),
    .B1(_08446_),
    .X(_08449_));
 sg13g2_nand2_1 _18498_ (.Y(_08450_),
    .A(_08165_),
    .B(_08449_));
 sg13g2_nand2_1 _18499_ (.Y(_08451_),
    .A(_08448_),
    .B(_08450_));
 sg13g2_a21o_1 _18500_ (.A2(_08173_),
    .A1(_08171_),
    .B1(_08169_),
    .X(_08452_));
 sg13g2_o21ai_1 _18501_ (.B1(_08452_),
    .Y(_08453_),
    .A1(_08171_),
    .A2(_08173_));
 sg13g2_or2_1 _18502_ (.X(_08455_),
    .B(_08453_),
    .A(_08194_));
 sg13g2_nand2_1 _18503_ (.Y(_08456_),
    .A(_08194_),
    .B(_08453_));
 sg13g2_nor2_1 _18504_ (.A(_08257_),
    .B(_08268_),
    .Y(_08457_));
 sg13g2_a21oi_2 _18505_ (.B1(_08457_),
    .Y(_08458_),
    .A2(_08255_),
    .A1(_08246_));
 sg13g2_nand2_1 _18506_ (.Y(_08459_),
    .A(_08455_),
    .B(_08458_));
 sg13g2_nand3_1 _18507_ (.B(_08456_),
    .C(_08459_),
    .A(_08451_),
    .Y(_08460_));
 sg13g2_inv_1 _18508_ (.Y(_08461_),
    .A(_08460_));
 sg13g2_a21o_1 _18509_ (.A2(_08459_),
    .A1(_08456_),
    .B1(_08451_),
    .X(_08462_));
 sg13g2_a21o_1 _18510_ (.A2(_08222_),
    .A1(_08211_),
    .B1(_08233_),
    .X(_08463_));
 sg13g2_o21ai_1 _18511_ (.B1(_08463_),
    .Y(_08464_),
    .A1(_08211_),
    .A2(_08222_));
 sg13g2_nand2_1 _18512_ (.Y(_08466_),
    .A(_08295_),
    .B(_08306_));
 sg13g2_nand3_1 _18513_ (.B(_08464_),
    .C(_08466_),
    .A(_08296_),
    .Y(_08467_));
 sg13g2_a21o_1 _18514_ (.A2(_08466_),
    .A1(_08296_),
    .B1(_08464_),
    .X(_08468_));
 sg13g2_inv_1 _18515_ (.Y(_08469_),
    .A(_08468_));
 sg13g2_o21ai_1 _18516_ (.B1(_08329_),
    .Y(_08470_),
    .A1(_08328_),
    .A2(_08342_));
 sg13g2_a21oi_2 _18517_ (.B1(_08469_),
    .Y(_08471_),
    .A2(_08470_),
    .A1(_08467_));
 sg13g2_o21ai_1 _18518_ (.B1(_08462_),
    .Y(_08472_),
    .A1(_08461_),
    .A2(_08471_));
 sg13g2_a21oi_2 _18519_ (.B1(_08444_),
    .Y(_08473_),
    .A2(_08472_),
    .A1(_08441_));
 sg13g2_nor2b_1 _18520_ (.A(_07921_),
    .B_N(_07922_),
    .Y(_08474_));
 sg13g2_xnor2_1 _18521_ (.Y(_08475_),
    .A(_07965_),
    .B(_08474_));
 sg13g2_nand2_1 _18522_ (.Y(_08477_),
    .A(_07790_),
    .B(_07791_));
 sg13g2_xor2_1 _18523_ (.B(_08477_),
    .A(_07825_),
    .X(_08478_));
 sg13g2_nand2_1 _18524_ (.Y(_08479_),
    .A(_08475_),
    .B(_08478_));
 sg13g2_or2_1 _18525_ (.X(_08480_),
    .B(_08478_),
    .A(_08475_));
 sg13g2_nor2_1 _18526_ (.A(_08043_),
    .B(_08044_),
    .Y(_08481_));
 sg13g2_xor2_1 _18527_ (.B(_08481_),
    .A(_08078_),
    .X(_08482_));
 sg13g2_nand2_1 _18528_ (.Y(_08483_),
    .A(_08479_),
    .B(_08482_));
 sg13g2_nand2_1 _18529_ (.Y(_08484_),
    .A(_08480_),
    .B(_08483_));
 sg13g2_xnor2_1 _18530_ (.Y(_08485_),
    .A(_08200_),
    .B(_08357_));
 sg13g2_xnor2_1 _18531_ (.Y(_08486_),
    .A(_08365_),
    .B(_08485_));
 sg13g2_xor2_1 _18532_ (.B(_08416_),
    .A(_08397_),
    .X(_08488_));
 sg13g2_xnor2_1 _18533_ (.Y(_08489_),
    .A(_08439_),
    .B(_08488_));
 sg13g2_nand2b_1 _18534_ (.Y(_08490_),
    .B(_08489_),
    .A_N(_08486_));
 sg13g2_nand2b_1 _18535_ (.Y(_08491_),
    .B(_08486_),
    .A_N(_08489_));
 sg13g2_nand2_1 _18536_ (.Y(_08492_),
    .A(_08460_),
    .B(_08462_));
 sg13g2_xor2_1 _18537_ (.B(_08492_),
    .A(_08471_),
    .X(_08493_));
 sg13g2_nand2_1 _18538_ (.Y(_08494_),
    .A(_08490_),
    .B(_08493_));
 sg13g2_nand2_1 _18539_ (.Y(_08495_),
    .A(_08491_),
    .B(_08494_));
 sg13g2_or2_1 _18540_ (.X(_08496_),
    .B(_08495_),
    .A(_08484_));
 sg13g2_and2_1 _18541_ (.A(_08484_),
    .B(_08495_),
    .X(_08497_));
 sg13g2_nand2_1 _18542_ (.Y(_08499_),
    .A(_08381_),
    .B(_08384_));
 sg13g2_a21oi_2 _18543_ (.B1(_08403_),
    .Y(_08500_),
    .A2(_08405_),
    .A1(_08402_));
 sg13g2_a21o_1 _18544_ (.A2(_08412_),
    .A1(_08409_),
    .B1(_08221_),
    .X(_08501_));
 sg13g2_o21ai_1 _18545_ (.B1(_08501_),
    .Y(_08502_),
    .A1(_08409_),
    .A2(_08412_));
 sg13g2_nand2_1 _18546_ (.Y(_08503_),
    .A(_08500_),
    .B(_08502_));
 sg13g2_xor2_1 _18547_ (.B(_08502_),
    .A(_08500_),
    .X(_08504_));
 sg13g2_o21ai_1 _18548_ (.B1(_08372_),
    .Y(_08505_),
    .A1(_08371_),
    .A2(_08375_));
 sg13g2_xnor2_1 _18549_ (.Y(_08506_),
    .A(_08504_),
    .B(_08505_));
 sg13g2_a21oi_1 _18550_ (.A1(_08382_),
    .A2(_08499_),
    .Y(_08507_),
    .B1(_08506_));
 sg13g2_nand3_1 _18551_ (.B(_08499_),
    .C(_08506_),
    .A(_08382_),
    .Y(_08508_));
 sg13g2_nor2_1 _18552_ (.A(_08391_),
    .B(_08395_),
    .Y(_08510_));
 sg13g2_nor2_1 _18553_ (.A(_08392_),
    .B(_08510_),
    .Y(_08511_));
 sg13g2_o21ai_1 _18554_ (.B1(_08508_),
    .Y(_08512_),
    .A1(_08507_),
    .A2(_08511_));
 sg13g2_a21oi_2 _18555_ (.B1(_08497_),
    .Y(_08513_),
    .A2(_08512_),
    .A1(_08496_));
 sg13g2_nand2_1 _18556_ (.Y(_08514_),
    .A(_08448_),
    .B(_08449_));
 sg13g2_xnor2_1 _18557_ (.Y(_08515_),
    .A(_08165_),
    .B(_08514_));
 sg13g2_or2_1 _18558_ (.X(_08516_),
    .B(_08364_),
    .A(_08362_));
 sg13g2_a22oi_1 _18559_ (.Y(_08517_),
    .B1(_08365_),
    .B2(_08516_),
    .A2(_08364_),
    .A1(_08363_));
 sg13g2_nand2_1 _18560_ (.Y(_08518_),
    .A(_08515_),
    .B(_08517_));
 sg13g2_inv_1 _18561_ (.Y(_08519_),
    .A(_08518_));
 sg13g2_or2_1 _18562_ (.X(_08521_),
    .B(_08517_),
    .A(_08515_));
 sg13g2_nand2_1 _18563_ (.Y(_08522_),
    .A(_08455_),
    .B(_08456_));
 sg13g2_xor2_1 _18564_ (.B(_08522_),
    .A(_08458_),
    .X(_08523_));
 sg13g2_o21ai_1 _18565_ (.B1(_08521_),
    .Y(_08524_),
    .A1(_08519_),
    .A2(_08523_));
 sg13g2_nand3_1 _18566_ (.B(_07950_),
    .C(_07963_),
    .A(_07935_),
    .Y(_08525_));
 sg13g2_nor3_1 _18567_ (.A(_07935_),
    .B(_07950_),
    .C(_07963_),
    .Y(_08526_));
 sg13g2_o21ai_1 _18568_ (.B1(_08525_),
    .Y(_08527_),
    .A1(_07965_),
    .A2(_08526_));
 sg13g2_nand2_1 _18569_ (.Y(_08528_),
    .A(_07744_),
    .B(_07745_));
 sg13g2_xnor2_1 _18570_ (.Y(_08529_),
    .A(_07758_),
    .B(_08528_));
 sg13g2_nand2_1 _18571_ (.Y(_08530_),
    .A(_08527_),
    .B(_08529_));
 sg13g2_xor2_1 _18572_ (.B(_08529_),
    .A(_08527_),
    .X(_08532_));
 sg13g2_and2_1 _18573_ (.A(_07777_),
    .B(_07778_),
    .X(_08533_));
 sg13g2_xnor2_1 _18574_ (.Y(_08534_),
    .A(_07788_),
    .B(_08533_));
 sg13g2_xnor2_1 _18575_ (.Y(_08535_),
    .A(_08532_),
    .B(_08534_));
 sg13g2_or2_1 _18576_ (.X(_08536_),
    .B(_08005_),
    .A(_07990_));
 sg13g2_a22oi_1 _18577_ (.Y(_08537_),
    .B1(_08006_),
    .B2(_08536_),
    .A2(_08005_),
    .A1(_07991_));
 sg13g2_or2_1 _18578_ (.X(_08538_),
    .B(_07824_),
    .A(_07812_));
 sg13g2_a22oi_1 _18579_ (.Y(_08539_),
    .B1(_07825_),
    .B2(_08538_),
    .A2(_07824_),
    .A1(_07813_));
 sg13g2_nor2_1 _18580_ (.A(_08029_),
    .B(_08041_),
    .Y(_08540_));
 sg13g2_a21oi_1 _18581_ (.A1(_08030_),
    .A2(_08041_),
    .Y(_08541_),
    .B1(_08042_));
 sg13g2_nor2_1 _18582_ (.A(_08540_),
    .B(_08541_),
    .Y(_08543_));
 sg13g2_or2_1 _18583_ (.X(_08544_),
    .B(_08543_),
    .A(_08539_));
 sg13g2_inv_1 _18584_ (.Y(_08545_),
    .A(_08544_));
 sg13g2_nand2_1 _18585_ (.Y(_08546_),
    .A(_08539_),
    .B(_08543_));
 sg13g2_a21oi_2 _18586_ (.B1(_08545_),
    .Y(_08547_),
    .A2(_08546_),
    .A1(_08537_));
 sg13g2_inv_1 _18587_ (.Y(_08548_),
    .A(_08547_));
 sg13g2_or2_1 _18588_ (.X(_08549_),
    .B(_08546_),
    .A(_08537_));
 sg13g2_a22oi_1 _18589_ (.Y(_08550_),
    .B1(_08547_),
    .B2(_08549_),
    .A2(_08545_),
    .A1(_08537_));
 sg13g2_nand2_1 _18590_ (.Y(_08551_),
    .A(_08535_),
    .B(_08550_));
 sg13g2_xor2_1 _18591_ (.B(_08406_),
    .A(_08400_),
    .X(_08552_));
 sg13g2_xnor2_1 _18592_ (.Y(_08554_),
    .A(_08414_),
    .B(_08552_));
 sg13g2_o21ai_1 _18593_ (.B1(_08554_),
    .Y(_08555_),
    .A1(_08535_),
    .A2(_08550_));
 sg13g2_xnor2_1 _18594_ (.Y(_08556_),
    .A(_08437_),
    .B(_08438_));
 sg13g2_nor2_1 _18595_ (.A(_08154_),
    .B(_08155_),
    .Y(_08557_));
 sg13g2_xnor2_1 _18596_ (.Y(_08558_),
    .A(_08198_),
    .B(_08557_));
 sg13g2_nand2_1 _18597_ (.Y(_08559_),
    .A(_08556_),
    .B(_08558_));
 sg13g2_nor2_1 _18598_ (.A(_08556_),
    .B(_08558_),
    .Y(_08560_));
 sg13g2_nor2_1 _18599_ (.A(_08351_),
    .B(_08352_),
    .Y(_08561_));
 sg13g2_xor2_1 _18600_ (.B(_08561_),
    .A(_08354_),
    .X(_08562_));
 sg13g2_a21oi_1 _18601_ (.A1(_08559_),
    .A2(_08562_),
    .Y(_08563_),
    .B1(_08560_));
 sg13g2_and3_1 _18602_ (.X(_08565_),
    .A(_08551_),
    .B(_08555_),
    .C(_08563_));
 sg13g2_a21oi_1 _18603_ (.A1(_08551_),
    .A2(_08555_),
    .Y(_08566_),
    .B1(_08563_));
 sg13g2_nor2_1 _18604_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sg13g2_nor2_1 _18605_ (.A(_08524_),
    .B(_08566_),
    .Y(_08568_));
 sg13g2_nor2_1 _18606_ (.A(_08565_),
    .B(_08568_),
    .Y(_08569_));
 sg13g2_xnor2_1 _18607_ (.Y(_08570_),
    .A(_08524_),
    .B(_08567_));
 sg13g2_xnor2_1 _18608_ (.Y(_08571_),
    .A(_08535_),
    .B(_08550_));
 sg13g2_xnor2_1 _18609_ (.Y(_08572_),
    .A(_08554_),
    .B(_08571_));
 sg13g2_xor2_1 _18610_ (.B(_08558_),
    .A(_08556_),
    .X(_08573_));
 sg13g2_xnor2_1 _18611_ (.Y(_08574_),
    .A(_08562_),
    .B(_08573_));
 sg13g2_nand2_1 _18612_ (.Y(_08576_),
    .A(_08518_),
    .B(_08521_));
 sg13g2_xnor2_1 _18613_ (.Y(_08577_),
    .A(_08523_),
    .B(_08576_));
 sg13g2_nor2_1 _18614_ (.A(_08574_),
    .B(_08577_),
    .Y(_08578_));
 sg13g2_xnor2_1 _18615_ (.Y(_08579_),
    .A(_08574_),
    .B(_08577_));
 sg13g2_nand2_1 _18616_ (.Y(_08580_),
    .A(_07873_),
    .B(_07874_));
 sg13g2_xnor2_1 _18617_ (.Y(_08581_),
    .A(_07886_),
    .B(_08580_));
 sg13g2_nand2_1 _18618_ (.Y(_08582_),
    .A(_08467_),
    .B(_08468_));
 sg13g2_xnor2_1 _18619_ (.Y(_08583_),
    .A(_08470_),
    .B(_08582_));
 sg13g2_nand2_1 _18620_ (.Y(_08584_),
    .A(_08581_),
    .B(_08583_));
 sg13g2_xnor2_1 _18621_ (.Y(_08585_),
    .A(_08581_),
    .B(_08583_));
 sg13g2_nor2_1 _18622_ (.A(_07909_),
    .B(_07910_),
    .Y(_08587_));
 sg13g2_xnor2_1 _18623_ (.Y(_08588_),
    .A(_07918_),
    .B(_08587_));
 sg13g2_xnor2_1 _18624_ (.Y(_08589_),
    .A(_08585_),
    .B(_08588_));
 sg13g2_xnor2_1 _18625_ (.Y(_08590_),
    .A(_08579_),
    .B(_08589_));
 sg13g2_nand2_1 _18626_ (.Y(_08591_),
    .A(_08572_),
    .B(_08590_));
 sg13g2_xor2_1 _18627_ (.B(_08385_),
    .A(_08376_),
    .X(_08592_));
 sg13g2_xnor2_1 _18628_ (.Y(_08593_),
    .A(_08396_),
    .B(_08592_));
 sg13g2_nor2_1 _18629_ (.A(_08591_),
    .B(_08593_),
    .Y(_08594_));
 sg13g2_a21oi_2 _18630_ (.B1(_07854_),
    .Y(_08595_),
    .A2(_07858_),
    .A1(_07853_));
 sg13g2_nand2_1 _18631_ (.Y(_08596_),
    .A(_08594_),
    .B(_08595_));
 sg13g2_nor2_1 _18632_ (.A(_08572_),
    .B(_08590_),
    .Y(_08598_));
 sg13g2_a21oi_1 _18633_ (.A1(_08591_),
    .A2(_08593_),
    .Y(_08599_),
    .B1(_08598_));
 sg13g2_nand2_1 _18634_ (.Y(_08600_),
    .A(_08593_),
    .B(_08598_));
 sg13g2_nor2b_1 _18635_ (.A(_08599_),
    .B_N(_08600_),
    .Y(_08601_));
 sg13g2_nor2_1 _18636_ (.A(_08594_),
    .B(_08601_),
    .Y(_08602_));
 sg13g2_a21o_1 _18637_ (.A2(_08600_),
    .A1(_08595_),
    .B1(_08599_),
    .X(_08603_));
 sg13g2_nor2_1 _18638_ (.A(_08578_),
    .B(_08589_),
    .Y(_08604_));
 sg13g2_a21oi_2 _18639_ (.B1(_08604_),
    .Y(_08605_),
    .A2(_08577_),
    .A1(_08574_));
 sg13g2_a21oi_1 _18640_ (.A1(_08596_),
    .A2(_08603_),
    .Y(_08606_),
    .B1(_08605_));
 sg13g2_and3_1 _18641_ (.X(_08607_),
    .A(_08596_),
    .B(_08603_),
    .C(_08605_));
 sg13g2_or3_1 _18642_ (.A(_08570_),
    .B(_08606_),
    .C(_08607_),
    .X(_08609_));
 sg13g2_o21ai_1 _18643_ (.B1(_08570_),
    .Y(_08610_),
    .A1(_08606_),
    .A2(_08607_));
 sg13g2_o21ai_1 _18644_ (.B1(_08588_),
    .Y(_08611_),
    .A1(_08581_),
    .A2(_08583_));
 sg13g2_nand2_2 _18645_ (.Y(_08612_),
    .A(_08584_),
    .B(_08611_));
 sg13g2_nand2_1 _18646_ (.Y(_08613_),
    .A(_08530_),
    .B(_08534_));
 sg13g2_o21ai_1 _18647_ (.B1(_08613_),
    .Y(_08614_),
    .A1(_08527_),
    .A2(_08529_));
 sg13g2_nor2b_1 _18648_ (.A(_08612_),
    .B_N(_08614_),
    .Y(_08615_));
 sg13g2_nand2b_1 _18649_ (.Y(_08616_),
    .B(_08612_),
    .A_N(_08614_));
 sg13g2_nor2b_1 _18650_ (.A(_08615_),
    .B_N(_08616_),
    .Y(_08617_));
 sg13g2_xnor2_1 _18651_ (.Y(_08618_),
    .A(_08547_),
    .B(_08617_));
 sg13g2_a21o_1 _18652_ (.A2(_08610_),
    .A1(_08609_),
    .B1(_08618_),
    .X(_08620_));
 sg13g2_nand3_1 _18653_ (.B(_08610_),
    .C(_08618_),
    .A(_08609_),
    .Y(_08621_));
 sg13g2_nand2_1 _18654_ (.Y(_08622_),
    .A(_08490_),
    .B(_08491_));
 sg13g2_xor2_1 _18655_ (.B(_08622_),
    .A(_08493_),
    .X(_08623_));
 sg13g2_nand3_1 _18656_ (.B(_08621_),
    .C(_08623_),
    .A(_08620_),
    .Y(_08624_));
 sg13g2_a21o_1 _18657_ (.A2(_08621_),
    .A1(_08620_),
    .B1(_08623_),
    .X(_08625_));
 sg13g2_nand2_1 _18658_ (.Y(_08626_),
    .A(_08479_),
    .B(_08480_));
 sg13g2_xnor2_1 _18659_ (.Y(_08627_),
    .A(_08482_),
    .B(_08626_));
 sg13g2_inv_1 _18660_ (.Y(_08628_),
    .A(_08627_));
 sg13g2_nand3_1 _18661_ (.B(_08625_),
    .C(_08628_),
    .A(_08624_),
    .Y(_08629_));
 sg13g2_a21o_1 _18662_ (.A2(_08625_),
    .A1(_08624_),
    .B1(_08628_),
    .X(_08631_));
 sg13g2_nand2b_1 _18663_ (.Y(_08632_),
    .B(_08508_),
    .A_N(_08507_));
 sg13g2_xnor2_1 _18664_ (.Y(_08633_),
    .A(_08511_),
    .B(_08632_));
 sg13g2_a21oi_2 _18665_ (.B1(_08633_),
    .Y(_08634_),
    .A2(_08631_),
    .A1(_08629_));
 sg13g2_nand2_1 _18666_ (.Y(_08635_),
    .A(_08624_),
    .B(_08627_));
 sg13g2_and2_1 _18667_ (.A(_08625_),
    .B(_08635_),
    .X(_08636_));
 sg13g2_nor2b_1 _18668_ (.A(_08634_),
    .B_N(_08636_),
    .Y(_08637_));
 sg13g2_nor3_1 _18669_ (.A(_08625_),
    .B(_08628_),
    .C(_08633_),
    .Y(_08638_));
 sg13g2_nand2_1 _18670_ (.Y(_08639_),
    .A(_08609_),
    .B(_08618_));
 sg13g2_and2_1 _18671_ (.A(_08610_),
    .B(_08639_),
    .X(_08640_));
 sg13g2_nor2_1 _18672_ (.A(_08638_),
    .B(_08640_),
    .Y(_08642_));
 sg13g2_nor2_1 _18673_ (.A(_08637_),
    .B(_08642_),
    .Y(_08643_));
 sg13g2_o21ai_1 _18674_ (.B1(_08513_),
    .Y(_08644_),
    .A1(_08637_),
    .A2(_08642_));
 sg13g2_nor3_1 _18675_ (.A(_08513_),
    .B(_08637_),
    .C(_08642_),
    .Y(_08645_));
 sg13g2_xor2_1 _18676_ (.B(_08643_),
    .A(_08513_),
    .X(_08646_));
 sg13g2_nand2_1 _18677_ (.Y(_08647_),
    .A(_08603_),
    .B(_08605_));
 sg13g2_nand2_1 _18678_ (.Y(_08648_),
    .A(_08596_),
    .B(_08647_));
 sg13g2_nor2_1 _18679_ (.A(_08569_),
    .B(_08648_),
    .Y(_08649_));
 sg13g2_nand2_1 _18680_ (.Y(_08650_),
    .A(_08569_),
    .B(_08648_));
 sg13g2_a21oi_1 _18681_ (.A1(_08548_),
    .A2(_08616_),
    .Y(_08651_),
    .B1(_08615_));
 sg13g2_inv_1 _18682_ (.Y(_08653_),
    .A(_08651_));
 sg13g2_o21ai_1 _18683_ (.B1(_08650_),
    .Y(_08654_),
    .A1(_08649_),
    .A2(_08653_));
 sg13g2_xnor2_1 _18684_ (.Y(_08655_),
    .A(_08646_),
    .B(_08654_));
 sg13g2_xor2_1 _18685_ (.B(_08636_),
    .A(_08634_),
    .X(_08656_));
 sg13g2_xor2_1 _18686_ (.B(_08656_),
    .A(_08640_),
    .X(_08657_));
 sg13g2_xor2_1 _18687_ (.B(_08495_),
    .A(_08484_),
    .X(_08658_));
 sg13g2_xnor2_1 _18688_ (.Y(_08659_),
    .A(_08512_),
    .B(_08658_));
 sg13g2_nand2_1 _18689_ (.Y(_08660_),
    .A(_08657_),
    .B(_08659_));
 sg13g2_nor2_1 _18690_ (.A(_08657_),
    .B(_08659_),
    .Y(_08661_));
 sg13g2_xnor2_1 _18691_ (.Y(_08662_),
    .A(_08657_),
    .B(_08659_));
 sg13g2_nand2b_1 _18692_ (.Y(_08664_),
    .B(_08650_),
    .A_N(_08649_));
 sg13g2_xnor2_1 _18693_ (.Y(_08665_),
    .A(_08653_),
    .B(_08664_));
 sg13g2_inv_1 _18694_ (.Y(_08666_),
    .A(_08665_));
 sg13g2_xnor2_1 _18695_ (.Y(_08667_),
    .A(_08662_),
    .B(_08666_));
 sg13g2_xnor2_1 _18696_ (.Y(_08668_),
    .A(_08662_),
    .B(_08665_));
 sg13g2_or2_1 _18697_ (.X(_08669_),
    .B(_08472_),
    .A(_08441_));
 sg13g2_a22oi_1 _18698_ (.Y(_08670_),
    .B1(_08473_),
    .B2(_08669_),
    .A2(_08472_),
    .A1(_08444_));
 sg13g2_nand2_1 _18699_ (.Y(_08671_),
    .A(_07969_),
    .B(_08081_));
 sg13g2_o21ai_1 _18700_ (.B1(_08082_),
    .Y(_08672_),
    .A1(_07968_),
    .A2(_08081_));
 sg13g2_nand2_1 _18701_ (.Y(_08673_),
    .A(_08671_),
    .B(_08672_));
 sg13g2_nand2b_1 _18702_ (.Y(_08675_),
    .B(_08673_),
    .A_N(_08670_));
 sg13g2_nor2b_1 _18703_ (.A(_08673_),
    .B_N(_08670_),
    .Y(_08676_));
 sg13g2_xnor2_1 _18704_ (.Y(_08677_),
    .A(_08670_),
    .B(_08673_));
 sg13g2_o21ai_1 _18705_ (.B1(_08505_),
    .Y(_08678_),
    .A1(_08500_),
    .A2(_08502_));
 sg13g2_nand2_2 _18706_ (.Y(_08679_),
    .A(_08503_),
    .B(_08678_));
 sg13g2_xnor2_1 _18707_ (.Y(_08680_),
    .A(_08677_),
    .B(_08679_));
 sg13g2_inv_1 _18708_ (.Y(_08681_),
    .A(_08680_));
 sg13g2_o21ai_1 _18709_ (.B1(_08665_),
    .Y(_08682_),
    .A1(_08657_),
    .A2(_08659_));
 sg13g2_nand2_1 _18710_ (.Y(_08683_),
    .A(_08660_),
    .B(_08682_));
 sg13g2_a22oi_1 _18711_ (.Y(_08684_),
    .B1(_08682_),
    .B2(_08660_),
    .A2(_08680_),
    .A1(_08667_));
 sg13g2_o21ai_1 _18712_ (.B1(_08683_),
    .Y(_08686_),
    .A1(_08668_),
    .A2(_08681_));
 sg13g2_nand3_1 _18713_ (.B(_08666_),
    .C(_08680_),
    .A(_08661_),
    .Y(_08687_));
 sg13g2_inv_1 _18714_ (.Y(_08688_),
    .A(_08687_));
 sg13g2_a21o_1 _18715_ (.A2(_08679_),
    .A1(_08675_),
    .B1(_08676_),
    .X(_08689_));
 sg13g2_inv_1 _18716_ (.Y(_08690_),
    .A(_08689_));
 sg13g2_o21ai_1 _18717_ (.B1(_08689_),
    .Y(_08691_),
    .A1(_08684_),
    .A2(_08688_));
 sg13g2_nand3_1 _18718_ (.B(_08687_),
    .C(_08690_),
    .A(_08686_),
    .Y(_08692_));
 sg13g2_nor3_1 _18719_ (.A(_08684_),
    .B(_08688_),
    .C(_08690_),
    .Y(_08693_));
 sg13g2_a21oi_1 _18720_ (.A1(_08686_),
    .A2(_08687_),
    .Y(_08694_),
    .B1(_08689_));
 sg13g2_nor3_1 _18721_ (.A(_08655_),
    .B(_08693_),
    .C(_08694_),
    .Y(_08695_));
 sg13g2_and3_1 _18722_ (.X(_08697_),
    .A(_08655_),
    .B(_08691_),
    .C(_08692_));
 sg13g2_o21ai_1 _18723_ (.B1(_08655_),
    .Y(_08698_),
    .A1(_08693_),
    .A2(_08694_));
 sg13g2_nor3_1 _18724_ (.A(_08473_),
    .B(_08695_),
    .C(_08697_),
    .Y(_08699_));
 sg13g2_o21ai_1 _18725_ (.B1(_08473_),
    .Y(_08700_),
    .A1(_08695_),
    .A2(_08697_));
 sg13g2_nor2b_1 _18726_ (.A(_08699_),
    .B_N(_08700_),
    .Y(_08701_));
 sg13g2_nand3b_1 _18727_ (.B(_08700_),
    .C(_08083_),
    .Y(_08702_),
    .A_N(_08699_));
 sg13g2_xnor2_1 _18728_ (.Y(_08703_),
    .A(_08082_),
    .B(_08701_));
 sg13g2_inv_1 _18729_ (.Y(_08704_),
    .A(_08703_));
 sg13g2_xor2_1 _18730_ (.B(net2417),
    .A(net2522),
    .X(_08705_));
 sg13g2_nand2_2 _18731_ (.Y(_08706_),
    .A(net2491),
    .B(_05847_));
 sg13g2_and2_1 _18732_ (.A(_08705_),
    .B(_08706_),
    .X(_08708_));
 sg13g2_xnor2_1 _18733_ (.Y(_08709_),
    .A(net2385),
    .B(_07453_));
 sg13g2_nand2b_1 _18734_ (.Y(_08710_),
    .B(net2478),
    .A_N(net2366));
 sg13g2_xnor2_1 _18735_ (.Y(_08711_),
    .A(net2542),
    .B(net2487));
 sg13g2_xnor2_1 _18736_ (.Y(_08712_),
    .A(_08710_),
    .B(_08711_));
 sg13g2_nand2_1 _18737_ (.Y(_08713_),
    .A(_08709_),
    .B(_08712_));
 sg13g2_xor2_1 _18738_ (.B(_08712_),
    .A(_08709_),
    .X(_08714_));
 sg13g2_xnor2_1 _18739_ (.Y(_08715_),
    .A(_08708_),
    .B(_08714_));
 sg13g2_o21ai_1 _18740_ (.B1(_06238_),
    .Y(_08716_),
    .A1(net2451),
    .A2(net2536));
 sg13g2_nor2_1 _18741_ (.A(net2337),
    .B(net2798),
    .Y(_08717_));
 sg13g2_xnor2_1 _18742_ (.Y(_08719_),
    .A(net2337),
    .B(net2798));
 sg13g2_nand3_1 _18743_ (.B(_05506_),
    .C(_08719_),
    .A(net2227),
    .Y(_08720_));
 sg13g2_nor2_1 _18744_ (.A(_08716_),
    .B(_08720_),
    .Y(_08721_));
 sg13g2_xnor2_1 _18745_ (.Y(_08722_),
    .A(_08716_),
    .B(_08720_));
 sg13g2_nor2_1 _18746_ (.A(net2472),
    .B(net2423),
    .Y(_08723_));
 sg13g2_nor2_1 _18747_ (.A(net2432),
    .B(net2494),
    .Y(_08724_));
 sg13g2_xor2_1 _18748_ (.B(_08724_),
    .A(_08723_),
    .X(_08725_));
 sg13g2_xnor2_1 _18749_ (.Y(_08726_),
    .A(_08722_),
    .B(_08725_));
 sg13g2_nor2_1 _18750_ (.A(_08715_),
    .B(_08726_),
    .Y(_08727_));
 sg13g2_xnor2_1 _18751_ (.Y(_08728_),
    .A(_08715_),
    .B(_08726_));
 sg13g2_xnor2_1 _18752_ (.Y(_08730_),
    .A(net2378),
    .B(net2594));
 sg13g2_xnor2_1 _18753_ (.Y(_08731_),
    .A(net2568),
    .B(_08730_));
 sg13g2_o21ai_1 _18754_ (.B1(_00018_),
    .Y(_08732_),
    .A1(net2439),
    .A2(net2491));
 sg13g2_inv_1 _18755_ (.Y(_08733_),
    .A(_08732_));
 sg13g2_xnor2_1 _18756_ (.Y(_08734_),
    .A(net2452),
    .B(_08732_));
 sg13g2_xnor2_1 _18757_ (.Y(_08735_),
    .A(_08731_),
    .B(_08734_));
 sg13g2_xnor2_1 _18758_ (.Y(_08736_),
    .A(_08728_),
    .B(_08735_));
 sg13g2_nor2_1 _18759_ (.A(net2180),
    .B(net2707),
    .Y(_08737_));
 sg13g2_xnor2_1 _18760_ (.Y(_08738_),
    .A(_00014_),
    .B(_08737_));
 sg13g2_nor2_1 _18761_ (.A(net2469),
    .B(\net.in[252] ),
    .Y(_08739_));
 sg13g2_nand2_1 _18762_ (.Y(_08741_),
    .A(_08738_),
    .B(_08739_));
 sg13g2_nor2_1 _18763_ (.A(_08738_),
    .B(_08739_),
    .Y(_08742_));
 sg13g2_xor2_1 _18764_ (.B(_08739_),
    .A(_08738_),
    .X(_08743_));
 sg13g2_xnor2_1 _18765_ (.Y(_08744_),
    .A(net2469),
    .B(net2631));
 sg13g2_xnor2_1 _18766_ (.Y(_08745_),
    .A(_00421_),
    .B(_08744_));
 sg13g2_xnor2_1 _18767_ (.Y(_08746_),
    .A(_08743_),
    .B(_08745_));
 sg13g2_or2_1 _18768_ (.X(_08747_),
    .B(net2425),
    .A(net2477));
 sg13g2_a21oi_1 _18769_ (.A1(_05616_),
    .A2(net2801),
    .Y(_08748_),
    .B1(_08747_));
 sg13g2_o21ai_1 _18770_ (.B1(_08748_),
    .Y(_08749_),
    .A1(_05616_),
    .A2(net2801));
 sg13g2_nand2b_1 _18771_ (.Y(_08750_),
    .B(net2462),
    .A_N(net2478));
 sg13g2_nor2b_1 _18772_ (.A(net2462),
    .B_N(net2478),
    .Y(_08752_));
 sg13g2_o21ai_1 _18773_ (.B1(_08750_),
    .Y(_08753_),
    .A1(net2494),
    .A2(_05462_));
 sg13g2_nor2_1 _18774_ (.A(_08752_),
    .B(_08753_),
    .Y(_08754_));
 sg13g2_o21ai_1 _18775_ (.B1(_08749_),
    .Y(_08755_),
    .A1(_08752_),
    .A2(_08753_));
 sg13g2_nor3_1 _18776_ (.A(_08749_),
    .B(_08752_),
    .C(_08753_),
    .Y(_08756_));
 sg13g2_xor2_1 _18777_ (.B(_08754_),
    .A(_08749_),
    .X(_08757_));
 sg13g2_nor2_1 _18778_ (.A(net2498),
    .B(net2554),
    .Y(_08758_));
 sg13g2_nor2_1 _18779_ (.A(net2519),
    .B(net2712),
    .Y(_08759_));
 sg13g2_xnor2_1 _18780_ (.Y(_08760_),
    .A(_08758_),
    .B(_08759_));
 sg13g2_xnor2_1 _18781_ (.Y(_08761_),
    .A(_08757_),
    .B(_08760_));
 sg13g2_nand2_1 _18782_ (.Y(_08763_),
    .A(_08746_),
    .B(_08761_));
 sg13g2_xnor2_1 _18783_ (.Y(_08764_),
    .A(_08746_),
    .B(_08761_));
 sg13g2_a22oi_1 _18784_ (.Y(_08765_),
    .B1(net2378),
    .B2(_05770_),
    .A2(net2511),
    .A1(net2518));
 sg13g2_nand2b_1 _18785_ (.Y(_08766_),
    .B(net2262),
    .A_N(net2512));
 sg13g2_nor2b_1 _18786_ (.A(net2472),
    .B_N(net2626),
    .Y(_08767_));
 sg13g2_xnor2_1 _18787_ (.Y(_08768_),
    .A(_08766_),
    .B(_08767_));
 sg13g2_nor2_1 _18788_ (.A(_08765_),
    .B(_08768_),
    .Y(_08769_));
 sg13g2_xnor2_1 _18789_ (.Y(_08770_),
    .A(_08765_),
    .B(_08768_));
 sg13g2_xnor2_1 _18790_ (.Y(_08771_),
    .A(_00821_),
    .B(_08770_));
 sg13g2_xnor2_1 _18791_ (.Y(_08772_),
    .A(_08764_),
    .B(_08771_));
 sg13g2_nor2_1 _18792_ (.A(net2313),
    .B(\net.in[144] ),
    .Y(_08774_));
 sg13g2_nor2_1 _18793_ (.A(net2788),
    .B(net2564),
    .Y(_08775_));
 sg13g2_xor2_1 _18794_ (.B(_08775_),
    .A(_08774_),
    .X(_08776_));
 sg13g2_or2_1 _18795_ (.X(_08777_),
    .B(net2330),
    .A(net2578));
 sg13g2_a22oi_1 _18796_ (.Y(_08778_),
    .B1(net2330),
    .B2(net2578),
    .A2(net2683),
    .A1(net2490));
 sg13g2_xnor2_1 _18797_ (.Y(_08779_),
    .A(net2188),
    .B(net2278));
 sg13g2_xnor2_1 _18798_ (.Y(_08780_),
    .A(net2806),
    .B(_08779_));
 sg13g2_a21oi_1 _18799_ (.A1(_08777_),
    .A2(_08778_),
    .Y(_08781_),
    .B1(_08780_));
 sg13g2_nand3_1 _18800_ (.B(_08778_),
    .C(_08780_),
    .A(_08777_),
    .Y(_08782_));
 sg13g2_nor2b_1 _18801_ (.A(_08781_),
    .B_N(_08782_),
    .Y(_08783_));
 sg13g2_a21oi_1 _18802_ (.A1(_08776_),
    .A2(_08782_),
    .Y(_08785_),
    .B1(_08781_));
 sg13g2_xor2_1 _18803_ (.B(_08783_),
    .A(_08776_),
    .X(_08786_));
 sg13g2_nand2_1 _18804_ (.Y(_08787_),
    .A(net2808),
    .B(_05176_));
 sg13g2_nand2b_1 _18805_ (.Y(_08788_),
    .B(net2469),
    .A_N(net2626));
 sg13g2_nand2_1 _18806_ (.Y(_08789_),
    .A(_02559_),
    .B(_02783_));
 sg13g2_a21oi_1 _18807_ (.A1(_08787_),
    .A2(_08788_),
    .Y(_08790_),
    .B1(_08789_));
 sg13g2_and3_1 _18808_ (.X(_08791_),
    .A(_08787_),
    .B(_08788_),
    .C(_08789_));
 sg13g2_nor2_1 _18809_ (.A(_08790_),
    .B(_08791_),
    .Y(_08792_));
 sg13g2_nor2b_1 _18810_ (.A(net2730),
    .B_N(net2475),
    .Y(_08793_));
 sg13g2_xor2_1 _18811_ (.B(net2369),
    .A(net2533),
    .X(_08794_));
 sg13g2_xnor2_1 _18812_ (.Y(_08796_),
    .A(_08793_),
    .B(_08794_));
 sg13g2_xnor2_1 _18813_ (.Y(_08797_),
    .A(_08792_),
    .B(_08796_));
 sg13g2_nor2b_1 _18814_ (.A(_08786_),
    .B_N(_08797_),
    .Y(_08798_));
 sg13g2_nand2b_1 _18815_ (.Y(_08799_),
    .B(_08786_),
    .A_N(_08797_));
 sg13g2_xnor2_1 _18816_ (.Y(_08800_),
    .A(_08786_),
    .B(_08797_));
 sg13g2_nor2_1 _18817_ (.A(net2217),
    .B(net2239),
    .Y(_08801_));
 sg13g2_xnor2_1 _18818_ (.Y(_08802_),
    .A(net2337),
    .B(net2227));
 sg13g2_xor2_1 _18819_ (.B(net2511),
    .A(net2464),
    .X(_08803_));
 sg13g2_nor2_1 _18820_ (.A(_08802_),
    .B(_08803_),
    .Y(_08804_));
 sg13g2_nor2_1 _18821_ (.A(_05088_),
    .B(\net.in[112] ),
    .Y(_08805_));
 sg13g2_nor2_1 _18822_ (.A(_05330_),
    .B(net2660),
    .Y(_08807_));
 sg13g2_xnor2_1 _18823_ (.Y(_08808_),
    .A(_08805_),
    .B(_08807_));
 sg13g2_nand2b_1 _18824_ (.Y(_08809_),
    .B(_08808_),
    .A_N(_08804_));
 sg13g2_nor3_1 _18825_ (.A(_08802_),
    .B(_08803_),
    .C(_08808_),
    .Y(_08810_));
 sg13g2_xnor2_1 _18826_ (.Y(_08811_),
    .A(_08804_),
    .B(_08808_));
 sg13g2_xnor2_1 _18827_ (.Y(_08812_),
    .A(_08801_),
    .B(_08811_));
 sg13g2_xnor2_1 _18828_ (.Y(_08813_),
    .A(_08800_),
    .B(_08812_));
 sg13g2_nand2_1 _18829_ (.Y(_08814_),
    .A(_08772_),
    .B(_08813_));
 sg13g2_xnor2_1 _18830_ (.Y(_08815_),
    .A(_08772_),
    .B(_08813_));
 sg13g2_xnor2_1 _18831_ (.Y(_08816_),
    .A(_08736_),
    .B(_08815_));
 sg13g2_xnor2_1 _18832_ (.Y(_08818_),
    .A(net2469),
    .B(net2772));
 sg13g2_nand2b_1 _18833_ (.Y(_08819_),
    .B(net2404),
    .A_N(net2479));
 sg13g2_xor2_1 _18834_ (.B(net2247),
    .A(net2191),
    .X(_08820_));
 sg13g2_and3_1 _18835_ (.X(_08821_),
    .A(_00898_),
    .B(_08819_),
    .C(_08820_));
 sg13g2_nand3_1 _18836_ (.B(_08819_),
    .C(_08820_),
    .A(_00898_),
    .Y(_08822_));
 sg13g2_a21oi_1 _18837_ (.A1(_00898_),
    .A2(_08819_),
    .Y(_08823_),
    .B1(_08820_));
 sg13g2_nor2_1 _18838_ (.A(_08821_),
    .B(_08823_),
    .Y(_08824_));
 sg13g2_a22oi_1 _18839_ (.Y(_08825_),
    .B1(net2501),
    .B2(net2611),
    .A2(net2568),
    .A1(net2419));
 sg13g2_o21ai_1 _18840_ (.B1(_08825_),
    .Y(_08826_),
    .A1(net2420),
    .A2(net2568));
 sg13g2_a21oi_2 _18841_ (.B1(_08823_),
    .Y(_08827_),
    .A2(_08826_),
    .A1(_08822_));
 sg13g2_inv_1 _18842_ (.Y(_08829_),
    .A(_08827_));
 sg13g2_xnor2_1 _18843_ (.Y(_08830_),
    .A(_08824_),
    .B(_08826_));
 sg13g2_nor2_1 _18844_ (.A(net2423),
    .B(\net.in[252] ),
    .Y(_08831_));
 sg13g2_xor2_1 _18845_ (.B(\net.in[4] ),
    .A(net2518),
    .X(_08832_));
 sg13g2_xnor2_1 _18846_ (.Y(_08833_),
    .A(_08831_),
    .B(_08832_));
 sg13g2_nor2b_1 _18847_ (.A(net2471),
    .B_N(net2676),
    .Y(_08834_));
 sg13g2_a21oi_1 _18848_ (.A1(net2262),
    .A2(net2712),
    .Y(_08835_),
    .B1(_08834_));
 sg13g2_nor3_2 _18849_ (.A(net2470),
    .B(_05473_),
    .C(_08758_),
    .Y(_08836_));
 sg13g2_nand2b_1 _18850_ (.Y(_08837_),
    .B(_08836_),
    .A_N(_08835_));
 sg13g2_nor2b_1 _18851_ (.A(_08836_),
    .B_N(_08835_),
    .Y(_08838_));
 sg13g2_o21ai_1 _18852_ (.B1(_08837_),
    .Y(_08840_),
    .A1(_08833_),
    .A2(_08838_));
 sg13g2_xnor2_1 _18853_ (.Y(_08841_),
    .A(_08835_),
    .B(_08836_));
 sg13g2_xnor2_1 _18854_ (.Y(_08842_),
    .A(_08833_),
    .B(_08841_));
 sg13g2_a22oi_1 _18855_ (.Y(_08843_),
    .B1(_05847_),
    .B2(net2308),
    .A2(_05638_),
    .A1(_05385_));
 sg13g2_xnor2_1 _18856_ (.Y(_08844_),
    .A(net2334),
    .B(net2785));
 sg13g2_xor2_1 _18857_ (.B(net2599),
    .A(net2533),
    .X(_08845_));
 sg13g2_nor3_1 _18858_ (.A(net2451),
    .B(_08844_),
    .C(_08845_),
    .Y(_08846_));
 sg13g2_o21ai_1 _18859_ (.B1(_08845_),
    .Y(_08847_),
    .A1(net2451),
    .A2(_08844_));
 sg13g2_nand2b_1 _18860_ (.Y(_08848_),
    .B(_08847_),
    .A_N(_08846_));
 sg13g2_xnor2_1 _18861_ (.Y(_08849_),
    .A(_08843_),
    .B(_08848_));
 sg13g2_nor2b_1 _18862_ (.A(_08842_),
    .B_N(_08849_),
    .Y(_08851_));
 sg13g2_nand2b_1 _18863_ (.Y(_08852_),
    .B(_08842_),
    .A_N(_08849_));
 sg13g2_a21oi_1 _18864_ (.A1(_08830_),
    .A2(_08852_),
    .Y(_08853_),
    .B1(_08851_));
 sg13g2_xnor2_1 _18865_ (.Y(_08854_),
    .A(_08842_),
    .B(_08849_));
 sg13g2_xnor2_1 _18866_ (.Y(_08855_),
    .A(_08830_),
    .B(_08854_));
 sg13g2_xnor2_1 _18867_ (.Y(_08856_),
    .A(net2579),
    .B(net2377));
 sg13g2_xor2_1 _18868_ (.B(net2610),
    .A(net2551),
    .X(_08857_));
 sg13g2_nor2_1 _18869_ (.A(_08856_),
    .B(_08857_),
    .Y(_08858_));
 sg13g2_xor2_1 _18870_ (.B(net2436),
    .A(net2560),
    .X(_08859_));
 sg13g2_nand2b_1 _18871_ (.Y(_08860_),
    .B(net2653),
    .A_N(net2603));
 sg13g2_nor2b_1 _18872_ (.A(net2217),
    .B_N(net2672),
    .Y(_08862_));
 sg13g2_xnor2_1 _18873_ (.Y(_08863_),
    .A(_08860_),
    .B(_08862_));
 sg13g2_nor2b_1 _18874_ (.A(_08863_),
    .B_N(_08859_),
    .Y(_08864_));
 sg13g2_nand2b_1 _18875_ (.Y(_08865_),
    .B(_08863_),
    .A_N(_08859_));
 sg13g2_xnor2_1 _18876_ (.Y(_08866_),
    .A(_08859_),
    .B(_08863_));
 sg13g2_xnor2_1 _18877_ (.Y(_08867_),
    .A(_08858_),
    .B(_08866_));
 sg13g2_nand2b_1 _18878_ (.Y(_08868_),
    .B(net2594),
    .A_N(net2528));
 sg13g2_nand2b_1 _18879_ (.Y(_08869_),
    .B(net2378),
    .A_N(\net.in[126] ));
 sg13g2_a221oi_1 _18880_ (.B2(net2183),
    .C1(_02318_),
    .B1(_08869_),
    .A1(_05242_),
    .Y(_08870_),
    .A2(net2594));
 sg13g2_a221oi_1 _18881_ (.B2(_08868_),
    .C1(net2522),
    .B1(_02319_),
    .A1(_05088_),
    .Y(_08871_),
    .A2(net2378));
 sg13g2_nor2_1 _18882_ (.A(_08870_),
    .B(_08871_),
    .Y(_08873_));
 sg13g2_xnor2_1 _18883_ (.Y(_08874_),
    .A(net2385),
    .B(net2272));
 sg13g2_xnor2_1 _18884_ (.Y(_08875_),
    .A(_08873_),
    .B(_08874_));
 sg13g2_nor2_1 _18885_ (.A(_08867_),
    .B(_08875_),
    .Y(_08876_));
 sg13g2_nand2_1 _18886_ (.Y(_08877_),
    .A(_08867_),
    .B(_08875_));
 sg13g2_xor2_1 _18887_ (.B(_08875_),
    .A(_08867_),
    .X(_08878_));
 sg13g2_nor2_1 _18888_ (.A(net2755),
    .B(net2763),
    .Y(_08879_));
 sg13g2_xnor2_1 _18889_ (.Y(_08880_),
    .A(net2522),
    .B(net2334));
 sg13g2_xnor2_1 _18890_ (.Y(_08881_),
    .A(_08879_),
    .B(_08880_));
 sg13g2_xor2_1 _18891_ (.B(net2583),
    .A(net2478),
    .X(_08882_));
 sg13g2_nor3_2 _18892_ (.A(net2334),
    .B(net2420),
    .C(_08882_),
    .Y(_08884_));
 sg13g2_xor2_1 _18893_ (.B(net2607),
    .A(net2560),
    .X(_08885_));
 sg13g2_nand2_1 _18894_ (.Y(_08886_),
    .A(_08884_),
    .B(_08885_));
 sg13g2_nor2_1 _18895_ (.A(_08884_),
    .B(_08885_),
    .Y(_08887_));
 sg13g2_xnor2_1 _18896_ (.Y(_08888_),
    .A(_08884_),
    .B(_08885_));
 sg13g2_o21ai_1 _18897_ (.B1(_08886_),
    .Y(_08889_),
    .A1(_08881_),
    .A2(_08887_));
 sg13g2_xnor2_1 _18898_ (.Y(_08890_),
    .A(_08881_),
    .B(_08888_));
 sg13g2_xnor2_1 _18899_ (.Y(_08891_),
    .A(_08878_),
    .B(_08890_));
 sg13g2_nand2_1 _18900_ (.Y(_08892_),
    .A(_08855_),
    .B(_08891_));
 sg13g2_or2_1 _18901_ (.X(_08893_),
    .B(_08891_),
    .A(_08855_));
 sg13g2_nand2_1 _18902_ (.Y(_08895_),
    .A(_08892_),
    .B(_08893_));
 sg13g2_xnor2_1 _18903_ (.Y(_08896_),
    .A(_08818_),
    .B(_08895_));
 sg13g2_nand2_1 _18904_ (.Y(_08897_),
    .A(_08816_),
    .B(_08896_));
 sg13g2_xnor2_1 _18905_ (.Y(_08898_),
    .A(_08816_),
    .B(_08896_));
 sg13g2_xnor2_1 _18906_ (.Y(_08899_),
    .A(net2653),
    .B(net2718));
 sg13g2_nor2b_1 _18907_ (.A(net2385),
    .B_N(net2266),
    .Y(_08900_));
 sg13g2_nor2_1 _18908_ (.A(net2201),
    .B(net2710),
    .Y(_08901_));
 sg13g2_xnor2_1 _18909_ (.Y(_08902_),
    .A(_08900_),
    .B(_08901_));
 sg13g2_nor2_1 _18910_ (.A(_08899_),
    .B(_08902_),
    .Y(_08903_));
 sg13g2_nand2_1 _18911_ (.Y(_08904_),
    .A(_08899_),
    .B(_08902_));
 sg13g2_xor2_1 _18912_ (.B(_08902_),
    .A(_08899_),
    .X(_08906_));
 sg13g2_xnor2_1 _18913_ (.Y(_08907_),
    .A(net2515),
    .B(net2378));
 sg13g2_xnor2_1 _18914_ (.Y(_08908_),
    .A(_08906_),
    .B(_08907_));
 sg13g2_nor2b_1 _18915_ (.A(net2384),
    .B_N(net2723),
    .Y(_08909_));
 sg13g2_nor2_1 _18916_ (.A(net2423),
    .B(\net.in[225] ),
    .Y(_08910_));
 sg13g2_o21ai_1 _18917_ (.B1(_08910_),
    .Y(_08911_),
    .A1(net2297),
    .A2(net2266));
 sg13g2_nor2_1 _18918_ (.A(net2741),
    .B(net2188),
    .Y(_08912_));
 sg13g2_nor2b_1 _18919_ (.A(net2532),
    .B_N(net2242),
    .Y(_08913_));
 sg13g2_xnor2_1 _18920_ (.Y(_08914_),
    .A(_08912_),
    .B(_08913_));
 sg13g2_nand2_1 _18921_ (.Y(_08915_),
    .A(_08911_),
    .B(_08914_));
 sg13g2_nor2_1 _18922_ (.A(_08911_),
    .B(_08914_),
    .Y(_08917_));
 sg13g2_xor2_1 _18923_ (.B(_08914_),
    .A(_08911_),
    .X(_08918_));
 sg13g2_xnor2_1 _18924_ (.Y(_08919_),
    .A(_08909_),
    .B(_08918_));
 sg13g2_nand2_1 _18925_ (.Y(_08920_),
    .A(_08908_),
    .B(_08919_));
 sg13g2_or2_1 _18926_ (.X(_08921_),
    .B(_08919_),
    .A(_08908_));
 sg13g2_nand2_1 _18927_ (.Y(_08922_),
    .A(_08920_),
    .B(_08921_));
 sg13g2_nor3_2 _18928_ (.A(net2338),
    .B(net2423),
    .C(net2514),
    .Y(_08923_));
 sg13g2_o21ai_1 _18929_ (.B1(_07984_),
    .Y(_08924_),
    .A1(net2233),
    .A2(net2257));
 sg13g2_xor2_1 _18930_ (.B(net2632),
    .A(net2464),
    .X(_08925_));
 sg13g2_nand2_1 _18931_ (.Y(_08926_),
    .A(_08924_),
    .B(_08925_));
 sg13g2_nor2_1 _18932_ (.A(_08924_),
    .B(_08925_),
    .Y(_08928_));
 sg13g2_xor2_1 _18933_ (.B(_08925_),
    .A(_08924_),
    .X(_08929_));
 sg13g2_xnor2_1 _18934_ (.Y(_08930_),
    .A(_08923_),
    .B(_08929_));
 sg13g2_xor2_1 _18935_ (.B(_08930_),
    .A(_08922_),
    .X(_08931_));
 sg13g2_nor3_2 _18936_ (.A(_05308_),
    .B(net2383),
    .C(\net.in[10] ),
    .Y(_08932_));
 sg13g2_nor2_1 _18937_ (.A(_02517_),
    .B(_08932_),
    .Y(_08933_));
 sg13g2_nor2b_1 _18938_ (.A(net2400),
    .B_N(_08932_),
    .Y(_08934_));
 sg13g2_nor2_1 _18939_ (.A(_08933_),
    .B(_08934_),
    .Y(_08935_));
 sg13g2_a22oi_1 _18940_ (.Y(_08936_),
    .B1(net2224),
    .B2(net2178),
    .A2(net2293),
    .A1(net2680));
 sg13g2_nand4_1 _18941_ (.B(net2678),
    .C(net2293),
    .A(net2178),
    .Y(_08937_),
    .D(net2224));
 sg13g2_nor2b_2 _18942_ (.A(_08936_),
    .B_N(_08937_),
    .Y(_08939_));
 sg13g2_nor2_1 _18943_ (.A(_08934_),
    .B(_08939_),
    .Y(_08940_));
 sg13g2_nor2_2 _18944_ (.A(_08933_),
    .B(_08940_),
    .Y(_08941_));
 sg13g2_xor2_1 _18945_ (.B(_08939_),
    .A(_08935_),
    .X(_08942_));
 sg13g2_nand2b_1 _18946_ (.Y(_08943_),
    .B(net2227),
    .A_N(net2797));
 sg13g2_nor2_1 _18947_ (.A(_05484_),
    .B(net2754),
    .Y(_08944_));
 sg13g2_xnor2_1 _18948_ (.Y(_08945_),
    .A(_08943_),
    .B(_08944_));
 sg13g2_a22oi_1 _18949_ (.Y(_08946_),
    .B1(net2355),
    .B2(net2611),
    .A2(_05462_),
    .A1(net2730));
 sg13g2_nor2b_1 _18950_ (.A(net2375),
    .B_N(net2495),
    .Y(_08947_));
 sg13g2_xnor2_1 _18951_ (.Y(_08948_),
    .A(_01062_),
    .B(_08947_));
 sg13g2_nand2b_1 _18952_ (.Y(_08950_),
    .B(_08946_),
    .A_N(_08948_));
 sg13g2_nor2b_1 _18953_ (.A(_08946_),
    .B_N(_08948_),
    .Y(_08951_));
 sg13g2_xnor2_1 _18954_ (.Y(_08952_),
    .A(_08946_),
    .B(_08948_));
 sg13g2_xnor2_1 _18955_ (.Y(_08953_),
    .A(_08945_),
    .B(_08952_));
 sg13g2_o21ai_1 _18956_ (.B1(net2723),
    .Y(_08954_),
    .A1(_05209_),
    .A2(net2462));
 sg13g2_a21oi_1 _18957_ (.A1(_05209_),
    .A2(net2462),
    .Y(_08955_),
    .B1(net2811));
 sg13g2_nand2b_1 _18958_ (.Y(_08956_),
    .B(_08955_),
    .A_N(_08954_));
 sg13g2_nand2_1 _18959_ (.Y(_08957_),
    .A(\net.in[126] ),
    .B(net2179));
 sg13g2_nand2b_1 _18960_ (.Y(_08958_),
    .B(net2191),
    .A_N(net2404));
 sg13g2_xnor2_1 _18961_ (.Y(_08959_),
    .A(net2212),
    .B(net2429));
 sg13g2_xnor2_1 _18962_ (.Y(_08961_),
    .A(_08958_),
    .B(_08959_));
 sg13g2_nand2b_1 _18963_ (.Y(_08962_),
    .B(_08961_),
    .A_N(_08957_));
 sg13g2_a21oi_1 _18964_ (.A1(net2498),
    .A2(net2179),
    .Y(_08963_),
    .B1(_08961_));
 sg13g2_xnor2_1 _18965_ (.Y(_08964_),
    .A(_08957_),
    .B(_08961_));
 sg13g2_o21ai_1 _18966_ (.B1(_08962_),
    .Y(_08965_),
    .A1(_08956_),
    .A2(_08963_));
 sg13g2_xnor2_1 _18967_ (.Y(_08966_),
    .A(_08956_),
    .B(_08964_));
 sg13g2_inv_1 _18968_ (.Y(_08967_),
    .A(_08966_));
 sg13g2_nand2_1 _18969_ (.Y(_08968_),
    .A(_08953_),
    .B(_08967_));
 sg13g2_nand2b_1 _18970_ (.Y(_08969_),
    .B(_08966_),
    .A_N(_08953_));
 sg13g2_xnor2_1 _18971_ (.Y(_08970_),
    .A(_08953_),
    .B(_08966_));
 sg13g2_xnor2_1 _18972_ (.Y(_08972_),
    .A(_08942_),
    .B(_08970_));
 sg13g2_nand2b_1 _18973_ (.Y(_08973_),
    .B(net2420),
    .A_N(net2352));
 sg13g2_a21oi_1 _18974_ (.A1(_00011_),
    .A2(_08973_),
    .Y(_08974_),
    .B1(_06153_));
 sg13g2_nand3_1 _18975_ (.B(_06153_),
    .C(_08973_),
    .A(_00011_),
    .Y(_08975_));
 sg13g2_nand2b_1 _18976_ (.Y(_08976_),
    .B(_08975_),
    .A_N(_08974_));
 sg13g2_xor2_1 _18977_ (.B(net2794),
    .A(net2514),
    .X(_08977_));
 sg13g2_xnor2_1 _18978_ (.Y(_08978_),
    .A(_08976_),
    .B(_08977_));
 sg13g2_nand2b_1 _18979_ (.Y(_08979_),
    .B(_03914_),
    .A_N(_02783_));
 sg13g2_nor2_1 _18980_ (.A(net2465),
    .B(net2569),
    .Y(_08980_));
 sg13g2_nor3_2 _18981_ (.A(net2680),
    .B(_07888_),
    .C(_08980_),
    .Y(_08981_));
 sg13g2_o21ai_1 _18982_ (.B1(_07888_),
    .Y(_08983_),
    .A1(net2679),
    .A2(_08980_));
 sg13g2_nand2b_1 _18983_ (.Y(_08984_),
    .B(_08983_),
    .A_N(_08981_));
 sg13g2_xnor2_1 _18984_ (.Y(_08985_),
    .A(_08979_),
    .B(_08984_));
 sg13g2_nand2_1 _18985_ (.Y(_08986_),
    .A(_08978_),
    .B(_08985_));
 sg13g2_nor2_1 _18986_ (.A(_08978_),
    .B(_08985_),
    .Y(_08987_));
 sg13g2_xnor2_1 _18987_ (.Y(_08988_),
    .A(_08978_),
    .B(_08985_));
 sg13g2_nor2_1 _18988_ (.A(net2191),
    .B(net2511),
    .Y(_08989_));
 sg13g2_nand2_1 _18989_ (.Y(_08990_),
    .A(net2402),
    .B(_08989_));
 sg13g2_nor2_1 _18990_ (.A(net2399),
    .B(net2360),
    .Y(_08991_));
 sg13g2_nor2_1 _18991_ (.A(net2498),
    .B(net2233),
    .Y(_08992_));
 sg13g2_xnor2_1 _18992_ (.Y(_08994_),
    .A(_08991_),
    .B(_08992_));
 sg13g2_nand2b_1 _18993_ (.Y(_08995_),
    .B(_08994_),
    .A_N(_08990_));
 sg13g2_a21oi_1 _18994_ (.A1(net2402),
    .A2(_08989_),
    .Y(_08996_),
    .B1(_08994_));
 sg13g2_xnor2_1 _18995_ (.Y(_08997_),
    .A(_08990_),
    .B(_08994_));
 sg13g2_xnor2_1 _18996_ (.Y(_08998_),
    .A(_02009_),
    .B(_08997_));
 sg13g2_xnor2_1 _18997_ (.Y(_08999_),
    .A(_08988_),
    .B(_08998_));
 sg13g2_inv_1 _18998_ (.Y(_09000_),
    .A(_08999_));
 sg13g2_nand2b_1 _18999_ (.Y(_09001_),
    .B(_08999_),
    .A_N(_08972_));
 sg13g2_nand2_1 _19000_ (.Y(_09002_),
    .A(_08972_),
    .B(_09000_));
 sg13g2_xnor2_1 _19001_ (.Y(_09003_),
    .A(_08972_),
    .B(_08999_));
 sg13g2_xnor2_1 _19002_ (.Y(_09005_),
    .A(_08931_),
    .B(_09003_));
 sg13g2_nor2_2 _19003_ (.A(net2480),
    .B(_05275_),
    .Y(_09006_));
 sg13g2_xnor2_1 _19004_ (.Y(_09007_),
    .A(_00004_),
    .B(_09006_));
 sg13g2_xor2_1 _19005_ (.B(net2514),
    .A(net2424),
    .X(_09008_));
 sg13g2_nand2_1 _19006_ (.Y(_09009_),
    .A(_09007_),
    .B(_09008_));
 sg13g2_xnor2_1 _19007_ (.Y(_09010_),
    .A(_09007_),
    .B(_09008_));
 sg13g2_xnor2_1 _19008_ (.Y(_09011_),
    .A(_02559_),
    .B(_09010_));
 sg13g2_xor2_1 _19009_ (.B(net2419),
    .A(net2523),
    .X(_09012_));
 sg13g2_nor2_2 _19010_ (.A(_01145_),
    .B(_09012_),
    .Y(_09013_));
 sg13g2_nor2_1 _19011_ (.A(net2185),
    .B(net2423),
    .Y(_09014_));
 sg13g2_xor2_1 _19012_ (.B(net2327),
    .A(net2337),
    .X(_09016_));
 sg13g2_xnor2_1 _19013_ (.Y(_09017_),
    .A(_09014_),
    .B(_09016_));
 sg13g2_nand2b_1 _19014_ (.Y(_09018_),
    .B(net2487),
    .A_N(net2494));
 sg13g2_nor2_1 _19015_ (.A(net2451),
    .B(net2406),
    .Y(_09019_));
 sg13g2_xnor2_1 _19016_ (.Y(_09020_),
    .A(_09018_),
    .B(_09019_));
 sg13g2_nand2_1 _19017_ (.Y(_09021_),
    .A(_09017_),
    .B(_09020_));
 sg13g2_or2_1 _19018_ (.X(_09022_),
    .B(_09020_),
    .A(_09017_));
 sg13g2_nand2_1 _19019_ (.Y(_09023_),
    .A(_09021_),
    .B(_09022_));
 sg13g2_xor2_1 _19020_ (.B(_09023_),
    .A(_09013_),
    .X(_09024_));
 sg13g2_nor2_1 _19021_ (.A(_09011_),
    .B(_09024_),
    .Y(_09025_));
 sg13g2_nand2_1 _19022_ (.Y(_09027_),
    .A(_09011_),
    .B(_09024_));
 sg13g2_xnor2_1 _19023_ (.Y(_09028_),
    .A(_09011_),
    .B(_09024_));
 sg13g2_nor2_1 _19024_ (.A(net2514),
    .B(net2414),
    .Y(_09029_));
 sg13g2_xnor2_1 _19025_ (.Y(_09030_),
    .A(net2384),
    .B(_09029_));
 sg13g2_nand2_1 _19026_ (.Y(_09031_),
    .A(net2391),
    .B(net2313));
 sg13g2_a22oi_1 _19027_ (.Y(_09032_),
    .B1(_05330_),
    .B2(_05099_),
    .A2(_05319_),
    .A1(_05308_));
 sg13g2_a22oi_1 _19028_ (.Y(_09033_),
    .B1(_05341_),
    .B2(net2455),
    .A2(net2478),
    .A1(_05044_));
 sg13g2_o21ai_1 _19029_ (.B1(_09033_),
    .Y(_09034_),
    .A1(net2455),
    .A2(_05341_));
 sg13g2_a21oi_1 _19030_ (.A1(_09031_),
    .A2(_09032_),
    .Y(_09035_),
    .B1(_09034_));
 sg13g2_nand3_1 _19031_ (.B(_09032_),
    .C(_09034_),
    .A(_09031_),
    .Y(_09036_));
 sg13g2_nand2b_1 _19032_ (.Y(_09038_),
    .B(_09036_),
    .A_N(_09035_));
 sg13g2_xor2_1 _19033_ (.B(_09038_),
    .A(_09030_),
    .X(_09039_));
 sg13g2_xnor2_1 _19034_ (.Y(_09040_),
    .A(_09028_),
    .B(_09039_));
 sg13g2_nor2_1 _19035_ (.A(_05121_),
    .B(net2358),
    .Y(_09041_));
 sg13g2_xnor2_1 _19036_ (.Y(_09042_),
    .A(net2664),
    .B(_09041_));
 sg13g2_inv_1 _19037_ (.Y(_09043_),
    .A(_09042_));
 sg13g2_xor2_1 _19038_ (.B(net2478),
    .A(net2290),
    .X(_09044_));
 sg13g2_nor2_1 _19039_ (.A(net2498),
    .B(net2551),
    .Y(_09045_));
 sg13g2_nor2b_1 _19040_ (.A(net2334),
    .B_N(net2298),
    .Y(_09046_));
 sg13g2_xnor2_1 _19041_ (.Y(_09047_),
    .A(_09045_),
    .B(_09046_));
 sg13g2_nand2b_1 _19042_ (.Y(_09049_),
    .B(_09044_),
    .A_N(_09047_));
 sg13g2_nor2b_1 _19043_ (.A(_09044_),
    .B_N(_09047_),
    .Y(_09050_));
 sg13g2_xnor2_1 _19044_ (.Y(_09051_),
    .A(_09044_),
    .B(_09047_));
 sg13g2_xnor2_1 _19045_ (.Y(_09052_),
    .A(_09042_),
    .B(_09051_));
 sg13g2_inv_1 _19046_ (.Y(_09053_),
    .A(_09052_));
 sg13g2_nand2b_1 _19047_ (.Y(_09054_),
    .B(net2219),
    .A_N(net2765));
 sg13g2_nand2b_1 _19048_ (.Y(_09055_),
    .B(net2765),
    .A_N(net2219));
 sg13g2_nand3_1 _19049_ (.B(_09054_),
    .C(_09055_),
    .A(_00004_),
    .Y(_09056_));
 sg13g2_nand2_2 _19050_ (.Y(_09057_),
    .A(net2688),
    .B(_05154_));
 sg13g2_nor2_1 _19051_ (.A(_09056_),
    .B(_09057_),
    .Y(_09058_));
 sg13g2_xor2_1 _19052_ (.B(_09057_),
    .A(_09056_),
    .X(_09060_));
 sg13g2_xor2_1 _19053_ (.B(net2554),
    .A(net2507),
    .X(_09061_));
 sg13g2_xnor2_1 _19054_ (.Y(_09062_),
    .A(_09060_),
    .B(_09061_));
 sg13g2_nor2_1 _19055_ (.A(_09053_),
    .B(_09062_),
    .Y(_09063_));
 sg13g2_xor2_1 _19056_ (.B(_09062_),
    .A(_09052_),
    .X(_09064_));
 sg13g2_nor2_1 _19057_ (.A(net2529),
    .B(net2788),
    .Y(_09065_));
 sg13g2_nor2_1 _19058_ (.A(net2417),
    .B(net2611),
    .Y(_09066_));
 sg13g2_xnor2_1 _19059_ (.Y(_09067_),
    .A(_09065_),
    .B(_09066_));
 sg13g2_or2_1 _19060_ (.X(_09068_),
    .B(net2469),
    .A(net2333));
 sg13g2_nand2b_1 _19061_ (.Y(_09069_),
    .B(net2498),
    .A_N(net2475));
 sg13g2_nand2_1 _19062_ (.Y(_09071_),
    .A(net2338),
    .B(net2560));
 sg13g2_a22oi_1 _19063_ (.Y(_09072_),
    .B1(_05209_),
    .B2(_05220_),
    .A2(net2494),
    .A1(net2182));
 sg13g2_nand4_1 _19064_ (.B(_09069_),
    .C(_09071_),
    .A(_09068_),
    .Y(_09073_),
    .D(_09072_));
 sg13g2_a22oi_1 _19065_ (.Y(_09074_),
    .B1(_09071_),
    .B2(_09072_),
    .A2(_09069_),
    .A1(_09068_));
 sg13g2_or2_1 _19066_ (.X(_09075_),
    .B(_09073_),
    .A(_09067_));
 sg13g2_o21ai_1 _19067_ (.B1(_09073_),
    .Y(_09076_),
    .A1(_09067_),
    .A2(_09074_));
 sg13g2_and2_1 _19068_ (.A(_09067_),
    .B(_09074_),
    .X(_09077_));
 sg13g2_o21ai_1 _19069_ (.B1(_09075_),
    .Y(_09078_),
    .A1(_09076_),
    .A2(_09077_));
 sg13g2_xnor2_1 _19070_ (.Y(_09079_),
    .A(_09064_),
    .B(_09078_));
 sg13g2_nor2b_1 _19071_ (.A(net2808),
    .B_N(net2262),
    .Y(_09080_));
 sg13g2_nor2b_1 _19072_ (.A(net2455),
    .B_N(net2451),
    .Y(_09082_));
 sg13g2_nor2b_1 _19073_ (.A(net2451),
    .B_N(net2455),
    .Y(_09083_));
 sg13g2_nor2_1 _19074_ (.A(net2471),
    .B(net2751),
    .Y(_09084_));
 sg13g2_nor3_2 _19075_ (.A(_09082_),
    .B(_09083_),
    .C(_09084_),
    .Y(_09085_));
 sg13g2_nand2_1 _19076_ (.Y(_09086_),
    .A(_08705_),
    .B(_09085_));
 sg13g2_nor2_1 _19077_ (.A(_08705_),
    .B(_09085_),
    .Y(_09087_));
 sg13g2_xor2_1 _19078_ (.B(_09085_),
    .A(_08705_),
    .X(_09088_));
 sg13g2_xnor2_1 _19079_ (.Y(_09089_),
    .A(_09080_),
    .B(_09088_));
 sg13g2_xnor2_1 _19080_ (.Y(_09090_),
    .A(_04094_),
    .B(_06473_));
 sg13g2_nand2_1 _19081_ (.Y(_09091_),
    .A(_01200_),
    .B(_09090_));
 sg13g2_xnor2_1 _19082_ (.Y(_09093_),
    .A(_01200_),
    .B(_09090_));
 sg13g2_xnor2_1 _19083_ (.Y(_09094_),
    .A(_02229_),
    .B(_09093_));
 sg13g2_nor2_1 _19084_ (.A(_09089_),
    .B(_09094_),
    .Y(_09095_));
 sg13g2_xor2_1 _19085_ (.B(_09094_),
    .A(_09089_),
    .X(_09096_));
 sg13g2_a22oi_1 _19086_ (.Y(_09097_),
    .B1(net2752),
    .B2(net2499),
    .A2(_05077_),
    .A1(net2305));
 sg13g2_o21ai_1 _19087_ (.B1(_09097_),
    .Y(_09098_),
    .A1(net2305),
    .A2(_05077_));
 sg13g2_o21ai_1 _19088_ (.B1(_00002_),
    .Y(_09099_),
    .A1(net2452),
    .A2(net2486));
 sg13g2_nand2b_1 _19089_ (.Y(_09100_),
    .B(_09099_),
    .A_N(_09098_));
 sg13g2_nor2b_1 _19090_ (.A(_09099_),
    .B_N(_09098_),
    .Y(_09101_));
 sg13g2_xor2_1 _19091_ (.B(_09099_),
    .A(_09098_),
    .X(_09102_));
 sg13g2_xnor2_1 _19092_ (.Y(_09104_),
    .A(_09719_),
    .B(_09102_));
 sg13g2_xnor2_1 _19093_ (.Y(_09105_),
    .A(_09096_),
    .B(_09104_));
 sg13g2_or2_1 _19094_ (.X(_09106_),
    .B(_09105_),
    .A(_09079_));
 sg13g2_nand2_1 _19095_ (.Y(_09107_),
    .A(_09079_),
    .B(_09105_));
 sg13g2_xnor2_1 _19096_ (.Y(_09108_),
    .A(_09079_),
    .B(_09105_));
 sg13g2_xnor2_1 _19097_ (.Y(_09109_),
    .A(_09040_),
    .B(_09108_));
 sg13g2_nor2b_1 _19098_ (.A(_09005_),
    .B_N(_09109_),
    .Y(_09110_));
 sg13g2_nand2b_1 _19099_ (.Y(_09111_),
    .B(_09005_),
    .A_N(_09109_));
 sg13g2_xnor2_1 _19100_ (.Y(_09112_),
    .A(_09005_),
    .B(_09109_));
 sg13g2_nor2b_1 _19101_ (.A(net2385),
    .B_N(net2670),
    .Y(_09113_));
 sg13g2_nor2_1 _19102_ (.A(_02445_),
    .B(_09113_),
    .Y(_09115_));
 sg13g2_nand2_1 _19103_ (.Y(_09116_),
    .A(_02445_),
    .B(_09113_));
 sg13g2_nor2b_1 _19104_ (.A(_09115_),
    .B_N(_09116_),
    .Y(_09117_));
 sg13g2_xor2_1 _19105_ (.B(net2657),
    .A(net2475),
    .X(_09118_));
 sg13g2_xnor2_1 _19106_ (.Y(_09119_),
    .A(_08717_),
    .B(_09118_));
 sg13g2_xnor2_1 _19107_ (.Y(_09120_),
    .A(_09117_),
    .B(_09119_));
 sg13g2_xor2_1 _19108_ (.B(net2223),
    .A(\net.in[44] ),
    .X(_09121_));
 sg13g2_nor2_1 _19109_ (.A(_01234_),
    .B(_09121_),
    .Y(_09122_));
 sg13g2_nand2_1 _19110_ (.Y(_09123_),
    .A(_01234_),
    .B(_09121_));
 sg13g2_nor2b_1 _19111_ (.A(_09122_),
    .B_N(_09123_),
    .Y(_09124_));
 sg13g2_nor2_1 _19112_ (.A(net2524),
    .B(net2469),
    .Y(_09126_));
 sg13g2_xnor2_1 _19113_ (.Y(_09127_),
    .A(_08834_),
    .B(_09126_));
 sg13g2_xnor2_1 _19114_ (.Y(_09128_),
    .A(_09124_),
    .B(_09127_));
 sg13g2_nor2_1 _19115_ (.A(_09120_),
    .B(_09128_),
    .Y(_09129_));
 sg13g2_nand2_1 _19116_ (.Y(_09130_),
    .A(_09120_),
    .B(_09128_));
 sg13g2_nand2b_1 _19117_ (.Y(_09131_),
    .B(_09130_),
    .A_N(_09129_));
 sg13g2_nand2_1 _19118_ (.Y(_09132_),
    .A(net2181),
    .B(net2257));
 sg13g2_nand2_1 _19119_ (.Y(_09133_),
    .A(_05143_),
    .B(net2636));
 sg13g2_o21ai_1 _19120_ (.B1(_00012_),
    .Y(_09134_),
    .A1(net2511),
    .A2(_05539_));
 sg13g2_a21o_2 _19121_ (.A2(_05539_),
    .A1(net2511),
    .B1(_09134_),
    .X(_09135_));
 sg13g2_a21oi_1 _19122_ (.A1(_09132_),
    .A2(_09133_),
    .Y(_09137_),
    .B1(_09135_));
 sg13g2_nand3_1 _19123_ (.B(_09133_),
    .C(_09135_),
    .A(_09132_),
    .Y(_09138_));
 sg13g2_nor2b_2 _19124_ (.A(_09137_),
    .B_N(_09138_),
    .Y(_09139_));
 sg13g2_xnor2_1 _19125_ (.Y(_09140_),
    .A(_02347_),
    .B(_09139_));
 sg13g2_xnor2_1 _19126_ (.Y(_09141_),
    .A(_09131_),
    .B(_09140_));
 sg13g2_nor4_2 _19127_ (.A(net2475),
    .B(net2186),
    .C(net2427),
    .Y(_09142_),
    .D(net2817));
 sg13g2_nor2_1 _19128_ (.A(net2518),
    .B(net2201),
    .Y(_09143_));
 sg13g2_o21ai_1 _19129_ (.B1(_09143_),
    .Y(_09144_),
    .A1(net2257),
    .A2(net2490));
 sg13g2_xnor2_1 _19130_ (.Y(_09145_),
    .A(net2420),
    .B(net2772));
 sg13g2_xnor2_1 _19131_ (.Y(_09146_),
    .A(net2213),
    .B(net2798));
 sg13g2_nand2_1 _19132_ (.Y(_09148_),
    .A(_09145_),
    .B(_09146_));
 sg13g2_nand2_1 _19133_ (.Y(_09149_),
    .A(_09144_),
    .B(_09148_));
 sg13g2_xor2_1 _19134_ (.B(_09148_),
    .A(_09144_),
    .X(_09150_));
 sg13g2_xnor2_1 _19135_ (.Y(_09151_),
    .A(_09142_),
    .B(_09150_));
 sg13g2_xor2_1 _19136_ (.B(\net.in[22] ),
    .A(net2514),
    .X(_09152_));
 sg13g2_xor2_1 _19137_ (.B(net2188),
    .A(net2213),
    .X(_09153_));
 sg13g2_nor2_2 _19138_ (.A(_09152_),
    .B(_09153_),
    .Y(_09154_));
 sg13g2_xnor2_1 _19139_ (.Y(_09155_),
    .A(net2333),
    .B(net2464));
 sg13g2_nor2_1 _19140_ (.A(net2337),
    .B(net2573),
    .Y(_09156_));
 sg13g2_nor2b_1 _19141_ (.A(net2427),
    .B_N(net2758),
    .Y(_09157_));
 sg13g2_xnor2_1 _19142_ (.Y(_09159_),
    .A(_09156_),
    .B(_09157_));
 sg13g2_nand2_1 _19143_ (.Y(_09160_),
    .A(_09155_),
    .B(_09159_));
 sg13g2_xnor2_1 _19144_ (.Y(_09161_),
    .A(_09155_),
    .B(_09159_));
 sg13g2_xor2_1 _19145_ (.B(_09161_),
    .A(_09154_),
    .X(_09162_));
 sg13g2_inv_1 _19146_ (.Y(_09163_),
    .A(_09162_));
 sg13g2_nor2b_1 _19147_ (.A(net2196),
    .B_N(net2217),
    .Y(_09164_));
 sg13g2_nor3_2 _19148_ (.A(net2423),
    .B(net2770),
    .C(_09164_),
    .Y(_09165_));
 sg13g2_a21oi_2 _19149_ (.B1(\net.in[161] ),
    .Y(_09166_),
    .A2(net2487),
    .A1(net2183));
 sg13g2_nor2b_1 _19150_ (.A(_09165_),
    .B_N(_09166_),
    .Y(_09167_));
 sg13g2_nor2b_1 _19151_ (.A(_09166_),
    .B_N(_09165_),
    .Y(_09168_));
 sg13g2_nor2_1 _19152_ (.A(_09167_),
    .B(_09168_),
    .Y(_09170_));
 sg13g2_xnor2_1 _19153_ (.Y(_09171_),
    .A(net2687),
    .B(_08856_));
 sg13g2_xnor2_1 _19154_ (.Y(_09172_),
    .A(_09170_),
    .B(_09171_));
 sg13g2_nand2_1 _19155_ (.Y(_09173_),
    .A(_09163_),
    .B(_09172_));
 sg13g2_nor2_1 _19156_ (.A(_09163_),
    .B(_09172_),
    .Y(_09174_));
 sg13g2_o21ai_1 _19157_ (.B1(_09173_),
    .Y(_09175_),
    .A1(_09151_),
    .A2(_09174_));
 sg13g2_xnor2_1 _19158_ (.Y(_09176_),
    .A(_09162_),
    .B(_09172_));
 sg13g2_xnor2_1 _19159_ (.Y(_09177_),
    .A(_09151_),
    .B(_09176_));
 sg13g2_o21ai_1 _19160_ (.B1(_00004_),
    .Y(_09178_),
    .A1(net2723),
    .A2(net2355));
 sg13g2_xor2_1 _19161_ (.B(net2579),
    .A(net2679),
    .X(_09179_));
 sg13g2_xor2_1 _19162_ (.B(\net.in[96] ),
    .A(net2578),
    .X(_09181_));
 sg13g2_xor2_1 _19163_ (.B(net2375),
    .A(net2475),
    .X(_09182_));
 sg13g2_xnor2_1 _19164_ (.Y(_09183_),
    .A(_09181_),
    .B(_09182_));
 sg13g2_inv_1 _19165_ (.Y(_09184_),
    .A(_09183_));
 sg13g2_nor2_1 _19166_ (.A(_09179_),
    .B(_09184_),
    .Y(_09185_));
 sg13g2_xnor2_1 _19167_ (.Y(_09186_),
    .A(_09179_),
    .B(_09183_));
 sg13g2_xnor2_1 _19168_ (.Y(_09187_),
    .A(_09178_),
    .B(_09186_));
 sg13g2_nor2_1 _19169_ (.A(net2424),
    .B(\net.in[161] ),
    .Y(_09188_));
 sg13g2_xor2_1 _19170_ (.B(net2568),
    .A(net2337),
    .X(_09189_));
 sg13g2_xnor2_1 _19171_ (.Y(_09190_),
    .A(_09188_),
    .B(_09189_));
 sg13g2_xnor2_1 _19172_ (.Y(_09192_),
    .A(net2399),
    .B(net2401));
 sg13g2_inv_1 _19173_ (.Y(_09193_),
    .A(_09192_));
 sg13g2_nor2_1 _19174_ (.A(net2494),
    .B(net2490),
    .Y(_09194_));
 sg13g2_nor2b_1 _19175_ (.A(net2423),
    .B_N(net2464),
    .Y(_09195_));
 sg13g2_xnor2_1 _19176_ (.Y(_09196_),
    .A(_09194_),
    .B(_09195_));
 sg13g2_nor2_1 _19177_ (.A(_09193_),
    .B(_09196_),
    .Y(_09197_));
 sg13g2_nand2_1 _19178_ (.Y(_09198_),
    .A(_09193_),
    .B(_09196_));
 sg13g2_o21ai_1 _19179_ (.B1(_09198_),
    .Y(_09199_),
    .A1(_09190_),
    .A2(_09197_));
 sg13g2_nor2b_1 _19180_ (.A(_09197_),
    .B_N(_09198_),
    .Y(_09200_));
 sg13g2_xnor2_1 _19181_ (.Y(_09201_),
    .A(_09190_),
    .B(_09200_));
 sg13g2_nand2_1 _19182_ (.Y(_09203_),
    .A(_09187_),
    .B(_09201_));
 sg13g2_xnor2_1 _19183_ (.Y(_09204_),
    .A(_09187_),
    .B(_09201_));
 sg13g2_nand2b_1 _19184_ (.Y(_09205_),
    .B(net2794),
    .A_N(net2735));
 sg13g2_xor2_1 _19185_ (.B(net2511),
    .A(net2469),
    .X(_09206_));
 sg13g2_xnor2_1 _19186_ (.Y(_09207_),
    .A(_09205_),
    .B(_09206_));
 sg13g2_nand2_1 _19187_ (.Y(_09208_),
    .A(net2427),
    .B(net2590));
 sg13g2_or2_1 _19188_ (.X(_09209_),
    .B(net2718),
    .A(net2355));
 sg13g2_xnor2_1 _19189_ (.Y(_09210_),
    .A(net2375),
    .B(net2583));
 sg13g2_and3_1 _19190_ (.X(_09211_),
    .A(_09208_),
    .B(_09209_),
    .C(_09210_));
 sg13g2_inv_1 _19191_ (.Y(_09212_),
    .A(_09211_));
 sg13g2_a21oi_1 _19192_ (.A1(_09208_),
    .A2(_09209_),
    .Y(_09214_),
    .B1(_09210_));
 sg13g2_o21ai_1 _19193_ (.B1(_09212_),
    .Y(_09215_),
    .A1(_09207_),
    .A2(_09214_));
 sg13g2_a21o_1 _19194_ (.A2(_09214_),
    .A1(_09207_),
    .B1(_09215_),
    .X(_09216_));
 sg13g2_o21ai_1 _19195_ (.B1(_09216_),
    .Y(_09217_),
    .A1(_09207_),
    .A2(_09212_));
 sg13g2_xnor2_1 _19196_ (.Y(_09218_),
    .A(_09204_),
    .B(_09217_));
 sg13g2_nand2_1 _19197_ (.Y(_09219_),
    .A(_09177_),
    .B(_09218_));
 sg13g2_nor2_1 _19198_ (.A(_09177_),
    .B(_09218_),
    .Y(_09220_));
 sg13g2_xor2_1 _19199_ (.B(_09218_),
    .A(_09177_),
    .X(_09221_));
 sg13g2_xnor2_1 _19200_ (.Y(_09222_),
    .A(_09141_),
    .B(_09221_));
 sg13g2_xnor2_1 _19201_ (.Y(_09223_),
    .A(_09112_),
    .B(_09222_));
 sg13g2_o21ai_1 _19202_ (.B1(_08897_),
    .Y(_09225_),
    .A1(_08898_),
    .A2(_09223_));
 sg13g2_a21o_1 _19203_ (.A2(_09222_),
    .A1(_09111_),
    .B1(_09110_),
    .X(_09226_));
 sg13g2_and2_1 _19204_ (.A(_09225_),
    .B(_09226_),
    .X(_09227_));
 sg13g2_xor2_1 _19205_ (.B(_09226_),
    .A(_09225_),
    .X(_09228_));
 sg13g2_xnor2_1 _19206_ (.Y(_09229_),
    .A(_09225_),
    .B(_09226_));
 sg13g2_o21ai_1 _19207_ (.B1(_09219_),
    .Y(_09230_),
    .A1(_09141_),
    .A2(_09220_));
 sg13g2_nand2_1 _19208_ (.Y(_09231_),
    .A(_09040_),
    .B(_09107_));
 sg13g2_nand2_1 _19209_ (.Y(_09232_),
    .A(_08931_),
    .B(_09002_));
 sg13g2_a22oi_1 _19210_ (.Y(_09233_),
    .B1(_09232_),
    .B2(_09001_),
    .A2(_09231_),
    .A1(_09106_));
 sg13g2_nand4_1 _19211_ (.B(_09106_),
    .C(_09231_),
    .A(_09001_),
    .Y(_09234_),
    .D(_09232_));
 sg13g2_nand2b_1 _19212_ (.Y(_09236_),
    .B(_09234_),
    .A_N(_09233_));
 sg13g2_xnor2_1 _19213_ (.Y(_09237_),
    .A(_09230_),
    .B(_09236_));
 sg13g2_nand2_1 _19214_ (.Y(_09238_),
    .A(_09228_),
    .B(_09237_));
 sg13g2_nor2_1 _19215_ (.A(_09095_),
    .B(_09104_),
    .Y(_09239_));
 sg13g2_a21oi_2 _19216_ (.B1(_09239_),
    .Y(_09240_),
    .A2(_09094_),
    .A1(_09089_));
 sg13g2_nand2_1 _19217_ (.Y(_09241_),
    .A(_08818_),
    .B(_08893_));
 sg13g2_o21ai_1 _19218_ (.B1(_08736_),
    .Y(_09242_),
    .A1(_08772_),
    .A2(_08813_));
 sg13g2_a22oi_1 _19219_ (.Y(_09243_),
    .B1(_09242_),
    .B2(_08814_),
    .A2(_09241_),
    .A1(_08892_));
 sg13g2_nand4_1 _19220_ (.B(_08892_),
    .C(_09241_),
    .A(_08814_),
    .Y(_09244_),
    .D(_09242_));
 sg13g2_nand2b_1 _19221_ (.Y(_09245_),
    .B(_09244_),
    .A_N(_09243_));
 sg13g2_xnor2_1 _19222_ (.Y(_09247_),
    .A(_09240_),
    .B(_09245_));
 sg13g2_o21ai_1 _19223_ (.B1(_09247_),
    .Y(_09248_),
    .A1(_09228_),
    .A2(_09237_));
 sg13g2_or2_1 _19224_ (.X(_09249_),
    .B(_08907_),
    .A(_08903_));
 sg13g2_a21oi_1 _19225_ (.A1(_08904_),
    .A2(_09249_),
    .Y(_09250_),
    .B1(_08941_));
 sg13g2_and3_1 _19226_ (.X(_09251_),
    .A(_08904_),
    .B(_08941_),
    .C(_09249_));
 sg13g2_nor2_1 _19227_ (.A(_09250_),
    .B(_09251_),
    .Y(_09252_));
 sg13g2_a21oi_2 _19228_ (.B1(_08917_),
    .Y(_09253_),
    .A2(_08915_),
    .A1(_08909_));
 sg13g2_xnor2_1 _19229_ (.Y(_09254_),
    .A(_09252_),
    .B(_09253_));
 sg13g2_nor2b_1 _19230_ (.A(_09168_),
    .B_N(_09171_),
    .Y(_09255_));
 sg13g2_a21oi_2 _19231_ (.B1(_08928_),
    .Y(_09256_),
    .A2(_08926_),
    .A1(_08923_));
 sg13g2_nor3_1 _19232_ (.A(_09167_),
    .B(_09255_),
    .C(_09256_),
    .Y(_09258_));
 sg13g2_o21ai_1 _19233_ (.B1(_09256_),
    .Y(_09259_),
    .A1(_09167_),
    .A2(_09255_));
 sg13g2_nand2b_1 _19234_ (.Y(_09260_),
    .B(_09259_),
    .A_N(_09258_));
 sg13g2_o21ai_1 _19235_ (.B1(_09154_),
    .Y(_09261_),
    .A1(_09155_),
    .A2(_09159_));
 sg13g2_nand2_1 _19236_ (.Y(_09262_),
    .A(_09160_),
    .B(_09261_));
 sg13g2_xnor2_1 _19237_ (.Y(_09263_),
    .A(_09260_),
    .B(_09262_));
 sg13g2_nor2_1 _19238_ (.A(_09254_),
    .B(_09263_),
    .Y(_09264_));
 sg13g2_nand2_1 _19239_ (.Y(_09265_),
    .A(_09254_),
    .B(_09263_));
 sg13g2_nand2b_1 _19240_ (.Y(_09266_),
    .B(_09265_),
    .A_N(_09264_));
 sg13g2_nand2_1 _19241_ (.Y(_09267_),
    .A(_09142_),
    .B(_09149_));
 sg13g2_o21ai_1 _19242_ (.B1(_09267_),
    .Y(_09269_),
    .A1(_09144_),
    .A2(_09148_));
 sg13g2_a21oi_1 _19243_ (.A1(_09179_),
    .A2(_09184_),
    .Y(_09270_),
    .B1(_09178_));
 sg13g2_or2_1 _19244_ (.X(_09271_),
    .B(_09270_),
    .A(_09185_));
 sg13g2_nor2_1 _19245_ (.A(_09269_),
    .B(_09271_),
    .Y(_09272_));
 sg13g2_inv_1 _19246_ (.Y(_09273_),
    .A(_09272_));
 sg13g2_and2_1 _19247_ (.A(_09269_),
    .B(_09271_),
    .X(_09274_));
 sg13g2_nor2_1 _19248_ (.A(_09272_),
    .B(_09274_),
    .Y(_09275_));
 sg13g2_xnor2_1 _19249_ (.Y(_09276_),
    .A(_09199_),
    .B(_09275_));
 sg13g2_xnor2_1 _19250_ (.Y(_09277_),
    .A(_09266_),
    .B(_09276_));
 sg13g2_nand2_1 _19251_ (.Y(_09278_),
    .A(_09013_),
    .B(_09021_));
 sg13g2_and3_1 _19252_ (.X(_09280_),
    .A(_09022_),
    .B(_09076_),
    .C(_09278_));
 sg13g2_a21o_1 _19253_ (.A2(_09278_),
    .A1(_09022_),
    .B1(_09076_),
    .X(_09281_));
 sg13g2_nor2b_1 _19254_ (.A(_09280_),
    .B_N(_09281_),
    .Y(_09282_));
 sg13g2_o21ai_1 _19255_ (.B1(_02559_),
    .Y(_09283_),
    .A1(_09007_),
    .A2(_09008_));
 sg13g2_nand2_1 _19256_ (.Y(_09284_),
    .A(_09009_),
    .B(_09283_));
 sg13g2_xnor2_1 _19257_ (.Y(_09285_),
    .A(_09282_),
    .B(_09284_));
 sg13g2_inv_1 _19258_ (.Y(_09286_),
    .A(_09285_));
 sg13g2_o21ai_1 _19259_ (.B1(_08983_),
    .Y(_09287_),
    .A1(_08979_),
    .A2(_08981_));
 sg13g2_a21oi_1 _19260_ (.A1(_08975_),
    .A2(_08977_),
    .Y(_09288_),
    .B1(_08974_));
 sg13g2_o21ai_1 _19261_ (.B1(_09036_),
    .Y(_09289_),
    .A1(_09030_),
    .A2(_09035_));
 sg13g2_and2_1 _19262_ (.A(_09288_),
    .B(_09289_),
    .X(_09291_));
 sg13g2_or2_1 _19263_ (.X(_09292_),
    .B(_09289_),
    .A(_09288_));
 sg13g2_a21oi_2 _19264_ (.B1(_09291_),
    .Y(_09293_),
    .A2(_09292_),
    .A1(_09287_));
 sg13g2_or2_1 _19265_ (.X(_09294_),
    .B(_09292_),
    .A(_09287_));
 sg13g2_a22oi_1 _19266_ (.Y(_09295_),
    .B1(_09293_),
    .B2(_09294_),
    .A2(_09291_),
    .A1(_09287_));
 sg13g2_nand2_1 _19267_ (.Y(_09296_),
    .A(_09286_),
    .B(_09295_));
 sg13g2_nor2_1 _19268_ (.A(_09286_),
    .B(_09295_),
    .Y(_09297_));
 sg13g2_xnor2_1 _19269_ (.Y(_09298_),
    .A(_09285_),
    .B(_09295_));
 sg13g2_a21oi_2 _19270_ (.B1(_08996_),
    .Y(_09299_),
    .A2(_08995_),
    .A1(_02009_));
 sg13g2_nor2_1 _19271_ (.A(_08965_),
    .B(_09299_),
    .Y(_09300_));
 sg13g2_xor2_1 _19272_ (.B(_09299_),
    .A(_08965_),
    .X(_09302_));
 sg13g2_o21ai_1 _19273_ (.B1(_08950_),
    .Y(_09303_),
    .A1(_08945_),
    .A2(_08951_));
 sg13g2_xnor2_1 _19274_ (.Y(_09304_),
    .A(_09302_),
    .B(_09303_));
 sg13g2_xnor2_1 _19275_ (.Y(_09305_),
    .A(_09298_),
    .B(_09304_));
 sg13g2_nand2_1 _19276_ (.Y(_09306_),
    .A(_09277_),
    .B(_09305_));
 sg13g2_or2_1 _19277_ (.X(_09307_),
    .B(_09305_),
    .A(_09277_));
 sg13g2_nor2_1 _19278_ (.A(_08791_),
    .B(_08796_),
    .Y(_09308_));
 sg13g2_or2_1 _19279_ (.X(_09309_),
    .B(_09308_),
    .A(_08790_));
 sg13g2_a21oi_1 _19280_ (.A1(_08765_),
    .A2(_08768_),
    .Y(_09310_),
    .B1(_00821_));
 sg13g2_o21ai_1 _19281_ (.B1(_09309_),
    .Y(_09311_),
    .A1(_08769_),
    .A2(_09310_));
 sg13g2_inv_1 _19282_ (.Y(_09313_),
    .A(_09311_));
 sg13g2_or3_1 _19283_ (.A(_08769_),
    .B(_09309_),
    .C(_09310_),
    .X(_09314_));
 sg13g2_nand2_1 _19284_ (.Y(_09315_),
    .A(_09311_),
    .B(_09314_));
 sg13g2_o21ai_1 _19285_ (.B1(_09314_),
    .Y(_09316_),
    .A1(_08785_),
    .A2(_09313_));
 sg13g2_xor2_1 _19286_ (.B(_09315_),
    .A(_08785_),
    .X(_09317_));
 sg13g2_a21oi_2 _19287_ (.B1(_09115_),
    .Y(_09318_),
    .A2(_09119_),
    .A1(_09116_));
 sg13g2_nor2_1 _19288_ (.A(_09215_),
    .B(_09318_),
    .Y(_09319_));
 sg13g2_xor2_1 _19289_ (.B(_09318_),
    .A(_09215_),
    .X(_09320_));
 sg13g2_o21ai_1 _19290_ (.B1(_09123_),
    .Y(_09321_),
    .A1(_09122_),
    .A2(_09127_));
 sg13g2_xnor2_1 _19291_ (.Y(_09322_),
    .A(_09320_),
    .B(_09321_));
 sg13g2_o21ai_1 _19292_ (.B1(_09138_),
    .Y(_09324_),
    .A1(_02347_),
    .A2(_09137_));
 sg13g2_a21oi_2 _19293_ (.B1(_08756_),
    .Y(_09325_),
    .A2(_08760_),
    .A1(_08755_));
 sg13g2_nor2_1 _19294_ (.A(_09324_),
    .B(_09325_),
    .Y(_09326_));
 sg13g2_xor2_1 _19295_ (.B(_09325_),
    .A(_09324_),
    .X(_09327_));
 sg13g2_o21ai_1 _19296_ (.B1(_08741_),
    .Y(_09328_),
    .A1(_08742_),
    .A2(_08745_));
 sg13g2_xnor2_1 _19297_ (.Y(_09329_),
    .A(_09327_),
    .B(_09328_));
 sg13g2_or2_1 _19298_ (.X(_09330_),
    .B(_09329_),
    .A(_09322_));
 sg13g2_nand2_1 _19299_ (.Y(_09331_),
    .A(_09322_),
    .B(_09329_));
 sg13g2_nand2_1 _19300_ (.Y(_09332_),
    .A(_09330_),
    .B(_09331_));
 sg13g2_xor2_1 _19301_ (.B(_09332_),
    .A(_09317_),
    .X(_09333_));
 sg13g2_nand2_1 _19302_ (.Y(_09335_),
    .A(_09307_),
    .B(_09333_));
 sg13g2_nand2_1 _19303_ (.Y(_09336_),
    .A(_09306_),
    .B(_09335_));
 sg13g2_nand3_1 _19304_ (.B(_09248_),
    .C(_09336_),
    .A(_09238_),
    .Y(_09337_));
 sg13g2_a21o_1 _19305_ (.A2(_09248_),
    .A1(_09238_),
    .B1(_09336_),
    .X(_09338_));
 sg13g2_a21oi_2 _19306_ (.B1(_08987_),
    .Y(_09339_),
    .A2(_08998_),
    .A1(_08986_));
 sg13g2_a21oi_1 _19307_ (.A1(_09027_),
    .A2(_09039_),
    .Y(_09340_),
    .B1(_09025_));
 sg13g2_a21oi_1 _19308_ (.A1(_09053_),
    .A2(_09062_),
    .Y(_09341_),
    .B1(_09078_));
 sg13g2_nor2_2 _19309_ (.A(_09063_),
    .B(_09341_),
    .Y(_09342_));
 sg13g2_nor2_1 _19310_ (.A(_09340_),
    .B(_09342_),
    .Y(_09343_));
 sg13g2_and2_1 _19311_ (.A(_09340_),
    .B(_09342_),
    .X(_09344_));
 sg13g2_nor2_1 _19312_ (.A(_09343_),
    .B(_09344_),
    .Y(_09346_));
 sg13g2_xnor2_1 _19313_ (.Y(_09347_),
    .A(_09339_),
    .B(_09346_));
 sg13g2_nand2_1 _19314_ (.Y(_09348_),
    .A(_08942_),
    .B(_08968_));
 sg13g2_nand2b_1 _19315_ (.Y(_09349_),
    .B(_08920_),
    .A_N(_08930_));
 sg13g2_a22oi_1 _19316_ (.Y(_09350_),
    .B1(_09349_),
    .B2(_08921_),
    .A2(_09348_),
    .A1(_08969_));
 sg13g2_nand4_1 _19317_ (.B(_08969_),
    .C(_09348_),
    .A(_08921_),
    .Y(_09351_),
    .D(_09349_));
 sg13g2_nand2b_1 _19318_ (.Y(_09352_),
    .B(_09351_),
    .A_N(_09350_));
 sg13g2_xnor2_1 _19319_ (.Y(_09353_),
    .A(_09175_),
    .B(_09352_));
 sg13g2_nor2_1 _19320_ (.A(_09347_),
    .B(_09353_),
    .Y(_09354_));
 sg13g2_nand2_1 _19321_ (.Y(_09355_),
    .A(_09347_),
    .B(_09353_));
 sg13g2_o21ai_1 _19322_ (.B1(_08771_),
    .Y(_09357_),
    .A1(_08746_),
    .A2(_08761_));
 sg13g2_nand2_2 _19323_ (.Y(_09358_),
    .A(_08763_),
    .B(_09357_));
 sg13g2_a21o_1 _19324_ (.A2(_09140_),
    .A1(_09130_),
    .B1(_09129_),
    .X(_09359_));
 sg13g2_o21ai_1 _19325_ (.B1(_09217_),
    .Y(_09360_),
    .A1(_09187_),
    .A2(_09201_));
 sg13g2_a21oi_1 _19326_ (.A1(_09203_),
    .A2(_09360_),
    .Y(_09361_),
    .B1(_09359_));
 sg13g2_nand3_1 _19327_ (.B(_09359_),
    .C(_09360_),
    .A(_09203_),
    .Y(_09362_));
 sg13g2_nor2b_1 _19328_ (.A(_09361_),
    .B_N(_09362_),
    .Y(_09363_));
 sg13g2_xnor2_1 _19329_ (.Y(_09364_),
    .A(_09358_),
    .B(_09363_));
 sg13g2_o21ai_1 _19330_ (.B1(_09355_),
    .Y(_09365_),
    .A1(_09354_),
    .A2(_09364_));
 sg13g2_nand2_1 _19331_ (.Y(_09366_),
    .A(_09337_),
    .B(_09365_));
 sg13g2_nand2_1 _19332_ (.Y(_09368_),
    .A(_09338_),
    .B(_09366_));
 sg13g2_nand2_1 _19333_ (.Y(_09369_),
    .A(_09306_),
    .B(_09307_));
 sg13g2_xor2_1 _19334_ (.B(_09369_),
    .A(_09333_),
    .X(_09370_));
 sg13g2_nor2b_1 _19335_ (.A(_09354_),
    .B_N(_09355_),
    .Y(_09371_));
 sg13g2_xnor2_1 _19336_ (.Y(_09372_),
    .A(_09364_),
    .B(_09371_));
 sg13g2_xnor2_1 _19337_ (.Y(_09373_),
    .A(_09229_),
    .B(_09237_));
 sg13g2_xnor2_1 _19338_ (.Y(_09374_),
    .A(_09247_),
    .B(_09373_));
 sg13g2_nor2b_1 _19339_ (.A(_09374_),
    .B_N(_09372_),
    .Y(_09375_));
 sg13g2_nand2b_1 _19340_ (.Y(_09376_),
    .B(_09374_),
    .A_N(_09372_));
 sg13g2_xnor2_1 _19341_ (.Y(_09377_),
    .A(_09372_),
    .B(_09374_));
 sg13g2_o21ai_1 _19342_ (.B1(_02229_),
    .Y(_09379_),
    .A1(_01200_),
    .A2(_09090_));
 sg13g2_a21oi_1 _19343_ (.A1(_09091_),
    .A2(_09379_),
    .Y(_09380_),
    .B1(_08853_));
 sg13g2_nand3_1 _19344_ (.B(_09091_),
    .C(_09379_),
    .A(_08853_),
    .Y(_09381_));
 sg13g2_nand2b_1 _19345_ (.Y(_09382_),
    .B(_09381_),
    .A_N(_09380_));
 sg13g2_a21oi_1 _19346_ (.A1(_09080_),
    .A2(_09086_),
    .Y(_09383_),
    .B1(_09087_));
 sg13g2_xnor2_1 _19347_ (.Y(_09384_),
    .A(_09382_),
    .B(_09383_));
 sg13g2_o21ai_1 _19348_ (.B1(_08877_),
    .Y(_09385_),
    .A1(_08876_),
    .A2(_08890_));
 sg13g2_a21oi_1 _19349_ (.A1(_08715_),
    .A2(_08726_),
    .Y(_09386_),
    .B1(_08735_));
 sg13g2_nor2_1 _19350_ (.A(_08727_),
    .B(_09386_),
    .Y(_09387_));
 sg13g2_o21ai_1 _19351_ (.B1(_08799_),
    .Y(_09388_),
    .A1(_08798_),
    .A2(_08812_));
 sg13g2_nand2_1 _19352_ (.Y(_09390_),
    .A(_09387_),
    .B(_09388_));
 sg13g2_inv_1 _19353_ (.Y(_09391_),
    .A(_09390_));
 sg13g2_or2_1 _19354_ (.X(_09392_),
    .B(_09388_),
    .A(_09387_));
 sg13g2_nand2_1 _19355_ (.Y(_09393_),
    .A(_09390_),
    .B(_09392_));
 sg13g2_xor2_1 _19356_ (.B(_09393_),
    .A(_09385_),
    .X(_09394_));
 sg13g2_nor2_1 _19357_ (.A(_09384_),
    .B(_09394_),
    .Y(_09395_));
 sg13g2_nand2_1 _19358_ (.Y(_09396_),
    .A(_09384_),
    .B(_09394_));
 sg13g2_nand2b_1 _19359_ (.Y(_09397_),
    .B(_09396_),
    .A_N(_09395_));
 sg13g2_a21oi_2 _19360_ (.B1(_09101_),
    .Y(_09398_),
    .A2(_09100_),
    .A1(_09719_));
 sg13g2_a21oi_1 _19361_ (.A1(_09043_),
    .A2(_09049_),
    .Y(_09399_),
    .B1(_09050_));
 sg13g2_and2_1 _19362_ (.A(_09398_),
    .B(_09399_),
    .X(_09401_));
 sg13g2_inv_1 _19363_ (.Y(_09402_),
    .A(_09401_));
 sg13g2_nor2_1 _19364_ (.A(_09398_),
    .B(_09399_),
    .Y(_09403_));
 sg13g2_nor2_1 _19365_ (.A(_09401_),
    .B(_09403_),
    .Y(_09404_));
 sg13g2_nor2_1 _19366_ (.A(_09058_),
    .B(_09061_),
    .Y(_09405_));
 sg13g2_a21oi_2 _19367_ (.B1(_09405_),
    .Y(_09406_),
    .A2(_09057_),
    .A1(_09056_));
 sg13g2_xor2_1 _19368_ (.B(_09406_),
    .A(_09404_),
    .X(_09407_));
 sg13g2_xnor2_1 _19369_ (.Y(_09408_),
    .A(_09397_),
    .B(_09407_));
 sg13g2_xnor2_1 _19370_ (.Y(_09409_),
    .A(_09377_),
    .B(_09408_));
 sg13g2_nand2b_1 _19371_ (.Y(_09410_),
    .B(_09409_),
    .A_N(_09370_));
 sg13g2_nor2b_1 _19372_ (.A(_09409_),
    .B_N(_09370_),
    .Y(_09412_));
 sg13g2_xor2_1 _19373_ (.B(_09409_),
    .A(_09370_),
    .X(_09413_));
 sg13g2_o21ai_1 _19374_ (.B1(_08847_),
    .Y(_09414_),
    .A1(_08843_),
    .A2(_08846_));
 sg13g2_and2_1 _19375_ (.A(_08840_),
    .B(_08889_),
    .X(_09415_));
 sg13g2_nor2_1 _19376_ (.A(_08840_),
    .B(_08889_),
    .Y(_09416_));
 sg13g2_nor2_1 _19377_ (.A(_09414_),
    .B(_09415_),
    .Y(_09417_));
 sg13g2_nor2_1 _19378_ (.A(_09416_),
    .B(_09417_),
    .Y(_09418_));
 sg13g2_nor2_1 _19379_ (.A(_09415_),
    .B(_09416_),
    .Y(_09419_));
 sg13g2_xnor2_1 _19380_ (.Y(_09420_),
    .A(_09414_),
    .B(_09419_));
 sg13g2_a21oi_1 _19381_ (.A1(_05099_),
    .A2(_08732_),
    .Y(_09421_),
    .B1(_08731_));
 sg13g2_a21oi_2 _19382_ (.B1(_09421_),
    .Y(_09423_),
    .A2(_08733_),
    .A1(net2452));
 sg13g2_nor2b_1 _19383_ (.A(_08871_),
    .B_N(_08874_),
    .Y(_09424_));
 sg13g2_o21ai_1 _19384_ (.B1(_09423_),
    .Y(_09425_),
    .A1(_08870_),
    .A2(_09424_));
 sg13g2_or3_1 _19385_ (.A(_08870_),
    .B(_09423_),
    .C(_09424_),
    .X(_09426_));
 sg13g2_nand2_1 _19386_ (.Y(_09427_),
    .A(_09425_),
    .B(_09426_));
 sg13g2_o21ai_1 _19387_ (.B1(_08865_),
    .Y(_09428_),
    .A1(_08858_),
    .A2(_08864_));
 sg13g2_xnor2_1 _19388_ (.Y(_09429_),
    .A(_09427_),
    .B(_09428_));
 sg13g2_inv_1 _19389_ (.Y(_09430_),
    .A(_09429_));
 sg13g2_nor2_1 _19390_ (.A(_08721_),
    .B(_08725_),
    .Y(_09431_));
 sg13g2_a21oi_1 _19391_ (.A1(_08716_),
    .A2(_08720_),
    .Y(_09432_),
    .B1(_09431_));
 sg13g2_inv_1 _19392_ (.Y(_09434_),
    .A(_09432_));
 sg13g2_or2_1 _19393_ (.X(_09435_),
    .B(_08810_),
    .A(_08801_));
 sg13g2_o21ai_1 _19394_ (.B1(_08708_),
    .Y(_09436_),
    .A1(_08709_),
    .A2(_08712_));
 sg13g2_nand4_1 _19395_ (.B(_08809_),
    .C(_09435_),
    .A(_08713_),
    .Y(_09437_),
    .D(_09436_));
 sg13g2_a22oi_1 _19396_ (.Y(_09438_),
    .B1(_09436_),
    .B2(_08713_),
    .A2(_09435_),
    .A1(_08809_));
 sg13g2_o21ai_1 _19397_ (.B1(_09437_),
    .Y(_09439_),
    .A1(_09434_),
    .A2(_09438_));
 sg13g2_o21ai_1 _19398_ (.B1(_09439_),
    .Y(_09440_),
    .A1(_09434_),
    .A2(_09437_));
 sg13g2_nand2_1 _19399_ (.Y(_09441_),
    .A(_09434_),
    .B(_09438_));
 sg13g2_nand2_2 _19400_ (.Y(_09442_),
    .A(_09440_),
    .B(_09441_));
 sg13g2_inv_1 _19401_ (.Y(_09443_),
    .A(_09442_));
 sg13g2_xnor2_1 _19402_ (.Y(_09445_),
    .A(_09429_),
    .B(_09442_));
 sg13g2_xnor2_1 _19403_ (.Y(_09446_),
    .A(_09420_),
    .B(_09445_));
 sg13g2_xnor2_1 _19404_ (.Y(_09447_),
    .A(_09413_),
    .B(_09446_));
 sg13g2_or2_1 _19405_ (.X(_09448_),
    .B(_09446_),
    .A(_09412_));
 sg13g2_nand3_1 _19406_ (.B(_09412_),
    .C(_09446_),
    .A(_08829_),
    .Y(_09449_));
 sg13g2_inv_1 _19407_ (.Y(_09450_),
    .A(_09449_));
 sg13g2_a22oi_1 _19408_ (.Y(_09451_),
    .B1(_09448_),
    .B2(_09410_),
    .A2(_09447_),
    .A1(_08829_));
 sg13g2_o21ai_1 _19409_ (.B1(_09376_),
    .Y(_09452_),
    .A1(_09375_),
    .A2(_09408_));
 sg13g2_a21o_1 _19410_ (.A2(_09452_),
    .A1(_09449_),
    .B1(_09451_),
    .X(_09453_));
 sg13g2_nor2b_1 _19411_ (.A(_09368_),
    .B_N(_09453_),
    .Y(_09454_));
 sg13g2_nand2b_1 _19412_ (.Y(_09456_),
    .B(_09368_),
    .A_N(_09453_));
 sg13g2_o21ai_1 _19413_ (.B1(_09396_),
    .Y(_09457_),
    .A1(_09395_),
    .A2(_09407_));
 sg13g2_a21oi_1 _19414_ (.A1(_09296_),
    .A2(_09304_),
    .Y(_09458_),
    .B1(_09297_));
 sg13g2_nor2_1 _19415_ (.A(_09457_),
    .B(_09458_),
    .Y(_09459_));
 sg13g2_a21oi_2 _19416_ (.B1(_09264_),
    .Y(_09460_),
    .A2(_09276_),
    .A1(_09265_));
 sg13g2_nand2_1 _19417_ (.Y(_09461_),
    .A(_09457_),
    .B(_09458_));
 sg13g2_o21ai_1 _19418_ (.B1(_09461_),
    .Y(_09462_),
    .A1(_09459_),
    .A2(_09460_));
 sg13g2_o21ai_1 _19419_ (.B1(_09456_),
    .Y(_09463_),
    .A1(_09454_),
    .A2(_09462_));
 sg13g2_nor2_1 _19420_ (.A(_09339_),
    .B(_09344_),
    .Y(_09464_));
 sg13g2_nor2_1 _19421_ (.A(_09343_),
    .B(_09464_),
    .Y(_09465_));
 sg13g2_a21oi_2 _19422_ (.B1(_09233_),
    .Y(_09467_),
    .A2(_09234_),
    .A1(_09230_));
 sg13g2_a21oi_2 _19423_ (.B1(_09243_),
    .Y(_09468_),
    .A2(_09244_),
    .A1(_09240_));
 sg13g2_nand2_1 _19424_ (.Y(_09469_),
    .A(_09467_),
    .B(_09468_));
 sg13g2_xor2_1 _19425_ (.B(_09468_),
    .A(_09467_),
    .X(_09470_));
 sg13g2_o21ai_1 _19426_ (.B1(_09465_),
    .Y(_09471_),
    .A1(_09467_),
    .A2(_09468_));
 sg13g2_nand2_1 _19427_ (.Y(_09472_),
    .A(_09469_),
    .B(_09471_));
 sg13g2_xnor2_1 _19428_ (.Y(_09473_),
    .A(_09465_),
    .B(_09470_));
 sg13g2_a21oi_1 _19429_ (.A1(_09430_),
    .A2(_09442_),
    .Y(_09474_),
    .B1(_09420_));
 sg13g2_a21oi_1 _19430_ (.A1(_09429_),
    .A2(_09443_),
    .Y(_09475_),
    .B1(_09474_));
 sg13g2_nand2_1 _19431_ (.Y(_09476_),
    .A(_09317_),
    .B(_09331_));
 sg13g2_a21o_1 _19432_ (.A2(_09476_),
    .A1(_09330_),
    .B1(_09475_),
    .X(_09478_));
 sg13g2_nand3_1 _19433_ (.B(_09475_),
    .C(_09476_),
    .A(_09330_),
    .Y(_09479_));
 sg13g2_nand2_1 _19434_ (.Y(_09480_),
    .A(_09478_),
    .B(_09479_));
 sg13g2_xnor2_1 _19435_ (.Y(_09481_),
    .A(_09227_),
    .B(_09480_));
 sg13g2_nor2_1 _19436_ (.A(_09473_),
    .B(_09481_),
    .Y(_09482_));
 sg13g2_and2_1 _19437_ (.A(_09473_),
    .B(_09481_),
    .X(_09483_));
 sg13g2_nor2_1 _19438_ (.A(_09482_),
    .B(_09483_),
    .Y(_09484_));
 sg13g2_a21oi_1 _19439_ (.A1(_09175_),
    .A2(_09351_),
    .Y(_09485_),
    .B1(_09350_));
 sg13g2_a21oi_1 _19440_ (.A1(_09358_),
    .A2(_09362_),
    .Y(_09486_),
    .B1(_09361_));
 sg13g2_nand2_1 _19441_ (.Y(_09487_),
    .A(_09485_),
    .B(_09486_));
 sg13g2_or2_1 _19442_ (.X(_09489_),
    .B(_09486_),
    .A(_09485_));
 sg13g2_nand2_1 _19443_ (.Y(_09490_),
    .A(_09487_),
    .B(_09489_));
 sg13g2_a21oi_2 _19444_ (.B1(_09391_),
    .Y(_09491_),
    .A2(_09392_),
    .A1(_09385_));
 sg13g2_xor2_1 _19445_ (.B(_09491_),
    .A(_09490_),
    .X(_09492_));
 sg13g2_xor2_1 _19446_ (.B(_09492_),
    .A(_09484_),
    .X(_09493_));
 sg13g2_nand2_1 _19447_ (.Y(_09494_),
    .A(_09337_),
    .B(_09338_));
 sg13g2_xor2_1 _19448_ (.B(_09494_),
    .A(_09365_),
    .X(_09495_));
 sg13g2_inv_1 _19449_ (.Y(_09496_),
    .A(_09495_));
 sg13g2_or3_1 _19450_ (.A(_09450_),
    .B(_09451_),
    .C(_09452_),
    .X(_09497_));
 sg13g2_o21ai_1 _19451_ (.B1(_09452_),
    .Y(_09498_),
    .A1(_09450_),
    .A2(_09451_));
 sg13g2_a21o_1 _19452_ (.A2(_09498_),
    .A1(_09497_),
    .B1(_09496_),
    .X(_09500_));
 sg13g2_nand3_1 _19453_ (.B(_09497_),
    .C(_09498_),
    .A(_09496_),
    .Y(_09501_));
 sg13g2_nand2b_1 _19454_ (.Y(_09502_),
    .B(_09461_),
    .A_N(_09459_));
 sg13g2_xnor2_1 _19455_ (.Y(_09503_),
    .A(_09460_),
    .B(_09502_));
 sg13g2_inv_1 _19456_ (.Y(_09504_),
    .A(_09503_));
 sg13g2_and3_1 _19457_ (.X(_09505_),
    .A(_09500_),
    .B(_09501_),
    .C(_09504_));
 sg13g2_a21oi_1 _19458_ (.A1(_09500_),
    .A2(_09501_),
    .Y(_09506_),
    .B1(_09504_));
 sg13g2_or3_1 _19459_ (.A(_09493_),
    .B(_09505_),
    .C(_09506_),
    .X(_09507_));
 sg13g2_o21ai_1 _19460_ (.B1(_09493_),
    .Y(_09508_),
    .A1(_09505_),
    .A2(_09506_));
 sg13g2_nor2_1 _19461_ (.A(_09300_),
    .B(_09303_),
    .Y(_09509_));
 sg13g2_a21oi_2 _19462_ (.B1(_09509_),
    .Y(_09511_),
    .A2(_09299_),
    .A1(_08965_));
 sg13g2_nand2_1 _19463_ (.Y(_09512_),
    .A(_09293_),
    .B(_09511_));
 sg13g2_xor2_1 _19464_ (.B(_09511_),
    .A(_09293_),
    .X(_09513_));
 sg13g2_nor2_1 _19465_ (.A(_09250_),
    .B(_09253_),
    .Y(_09514_));
 sg13g2_nor2_1 _19466_ (.A(_09251_),
    .B(_09514_),
    .Y(_09515_));
 sg13g2_xnor2_1 _19467_ (.Y(_09516_),
    .A(_09513_),
    .B(_09515_));
 sg13g2_o21ai_1 _19468_ (.B1(_09281_),
    .Y(_09517_),
    .A1(_09280_),
    .A2(_09284_));
 sg13g2_and2_1 _19469_ (.A(_09381_),
    .B(_09383_),
    .X(_09518_));
 sg13g2_a21oi_2 _19470_ (.B1(_09403_),
    .Y(_09519_),
    .A2(_09406_),
    .A1(_09402_));
 sg13g2_o21ai_1 _19471_ (.B1(_09519_),
    .Y(_09520_),
    .A1(_09380_),
    .A2(_09518_));
 sg13g2_nor3_1 _19472_ (.A(_09380_),
    .B(_09518_),
    .C(_09519_),
    .Y(_09522_));
 sg13g2_nor2_1 _19473_ (.A(_09517_),
    .B(_09520_),
    .Y(_09523_));
 sg13g2_o21ai_1 _19474_ (.B1(_09520_),
    .Y(_09524_),
    .A1(_09517_),
    .A2(_09522_));
 sg13g2_a21oi_1 _19475_ (.A1(_09517_),
    .A2(_09522_),
    .Y(_09525_),
    .B1(_09524_));
 sg13g2_nor2_2 _19476_ (.A(_09523_),
    .B(_09525_),
    .Y(_09526_));
 sg13g2_or2_1 _19477_ (.X(_09527_),
    .B(_09526_),
    .A(_09516_));
 sg13g2_nand2_1 _19478_ (.Y(_09528_),
    .A(_09516_),
    .B(_09526_));
 sg13g2_nand2_1 _19479_ (.Y(_09529_),
    .A(_09527_),
    .B(_09528_));
 sg13g2_a21oi_1 _19480_ (.A1(_09215_),
    .A2(_09318_),
    .Y(_09530_),
    .B1(_09321_));
 sg13g2_nor2_1 _19481_ (.A(_09319_),
    .B(_09530_),
    .Y(_09531_));
 sg13g2_a21oi_2 _19482_ (.B1(_09258_),
    .Y(_09533_),
    .A2(_09262_),
    .A1(_09259_));
 sg13g2_a21oi_2 _19483_ (.B1(_09274_),
    .Y(_09534_),
    .A2(_09273_),
    .A1(_09199_));
 sg13g2_nor2_1 _19484_ (.A(_09533_),
    .B(_09534_),
    .Y(_09535_));
 sg13g2_xor2_1 _19485_ (.B(_09534_),
    .A(_09533_),
    .X(_09536_));
 sg13g2_xnor2_1 _19486_ (.Y(_09537_),
    .A(_09531_),
    .B(_09536_));
 sg13g2_nand2_1 _19487_ (.Y(_09538_),
    .A(_09528_),
    .B(_09537_));
 sg13g2_xnor2_1 _19488_ (.Y(_09539_),
    .A(_09529_),
    .B(_09537_));
 sg13g2_nand3_1 _19489_ (.B(_09508_),
    .C(_09539_),
    .A(_09507_),
    .Y(_09540_));
 sg13g2_a21o_1 _19490_ (.A2(_09508_),
    .A1(_09507_),
    .B1(_09539_),
    .X(_09541_));
 sg13g2_nand2_1 _19491_ (.Y(_09542_),
    .A(_09425_),
    .B(_09428_));
 sg13g2_nand2_2 _19492_ (.Y(_09544_),
    .A(_09426_),
    .B(_09542_));
 sg13g2_nor2_1 _19493_ (.A(_09326_),
    .B(_09328_),
    .Y(_09545_));
 sg13g2_a21oi_2 _19494_ (.B1(_09545_),
    .Y(_09546_),
    .A2(_09325_),
    .A1(_09324_));
 sg13g2_and2_1 _19495_ (.A(_09316_),
    .B(_09546_),
    .X(_09547_));
 sg13g2_xnor2_1 _19496_ (.Y(_09548_),
    .A(_09316_),
    .B(_09546_));
 sg13g2_xnor2_1 _19497_ (.Y(_09549_),
    .A(_09439_),
    .B(_09548_));
 sg13g2_nor2_1 _19498_ (.A(_09544_),
    .B(_09549_),
    .Y(_09550_));
 sg13g2_xor2_1 _19499_ (.B(_09549_),
    .A(_09544_),
    .X(_09551_));
 sg13g2_xnor2_1 _19500_ (.Y(_09552_),
    .A(_09418_),
    .B(_09551_));
 sg13g2_a21oi_2 _19501_ (.B1(_09552_),
    .Y(_09553_),
    .A2(_09541_),
    .A1(_09540_));
 sg13g2_nand2_1 _19502_ (.Y(_09555_),
    .A(_09508_),
    .B(_09539_));
 sg13g2_and2_1 _19503_ (.A(_09507_),
    .B(_09555_),
    .X(_09556_));
 sg13g2_nor2_1 _19504_ (.A(_09553_),
    .B(_09556_),
    .Y(_09557_));
 sg13g2_nand2_1 _19505_ (.Y(_09558_),
    .A(_09500_),
    .B(_09503_));
 sg13g2_and2_1 _19506_ (.A(_09501_),
    .B(_09558_),
    .X(_09559_));
 sg13g2_nor2_1 _19507_ (.A(_09557_),
    .B(_09559_),
    .Y(_09560_));
 sg13g2_a21o_1 _19508_ (.A2(_09556_),
    .A1(_09553_),
    .B1(_09560_),
    .X(_09561_));
 sg13g2_nor2_1 _19509_ (.A(_09483_),
    .B(_09492_),
    .Y(_09562_));
 sg13g2_nor2_1 _19510_ (.A(_09482_),
    .B(_09562_),
    .Y(_09563_));
 sg13g2_a21oi_1 _19511_ (.A1(_09527_),
    .A2(_09538_),
    .Y(_09564_),
    .B1(_09563_));
 sg13g2_and3_1 _19512_ (.X(_09566_),
    .A(_09527_),
    .B(_09538_),
    .C(_09563_));
 sg13g2_a21oi_1 _19513_ (.A1(_09544_),
    .A2(_09549_),
    .Y(_09567_),
    .B1(_09418_));
 sg13g2_nor2_1 _19514_ (.A(_09550_),
    .B(_09567_),
    .Y(_09568_));
 sg13g2_nor2_1 _19515_ (.A(_09566_),
    .B(_09568_),
    .Y(_09569_));
 sg13g2_nor2_1 _19516_ (.A(_09564_),
    .B(_09569_),
    .Y(_09570_));
 sg13g2_and2_1 _19517_ (.A(_09561_),
    .B(_09570_),
    .X(_09571_));
 sg13g2_nor2_1 _19518_ (.A(_09561_),
    .B(_09570_),
    .Y(_09572_));
 sg13g2_nor2_1 _19519_ (.A(_09571_),
    .B(_09572_),
    .Y(_09573_));
 sg13g2_xnor2_1 _19520_ (.Y(_09574_),
    .A(_09463_),
    .B(_09573_));
 sg13g2_nand2_1 _19521_ (.Y(_09575_),
    .A(_09227_),
    .B(_09479_));
 sg13g2_nand3_1 _19522_ (.B(_09478_),
    .C(_09575_),
    .A(_09472_),
    .Y(_09577_));
 sg13g2_inv_1 _19523_ (.Y(_09578_),
    .A(_09577_));
 sg13g2_a21o_1 _19524_ (.A2(_09575_),
    .A1(_09478_),
    .B1(_09472_),
    .X(_09579_));
 sg13g2_nand2_1 _19525_ (.Y(_09580_),
    .A(_09577_),
    .B(_09579_));
 sg13g2_nand2_1 _19526_ (.Y(_09581_),
    .A(_09489_),
    .B(_09491_));
 sg13g2_nand2_1 _19527_ (.Y(_09582_),
    .A(_09487_),
    .B(_09581_));
 sg13g2_xnor2_1 _19528_ (.Y(_09583_),
    .A(_09580_),
    .B(_09582_));
 sg13g2_o21ai_1 _19529_ (.B1(_09515_),
    .Y(_09584_),
    .A1(_09293_),
    .A2(_09511_));
 sg13g2_nand2_1 _19530_ (.Y(_09585_),
    .A(_09512_),
    .B(_09584_));
 sg13g2_nand2_1 _19531_ (.Y(_09586_),
    .A(_09524_),
    .B(_09585_));
 sg13g2_or2_1 _19532_ (.X(_09588_),
    .B(_09585_),
    .A(_09524_));
 sg13g2_nand2_1 _19533_ (.Y(_09589_),
    .A(_09586_),
    .B(_09588_));
 sg13g2_nor2_1 _19534_ (.A(_09531_),
    .B(_09535_),
    .Y(_09590_));
 sg13g2_a21o_1 _19535_ (.A2(_09534_),
    .A1(_09533_),
    .B1(_09590_),
    .X(_09591_));
 sg13g2_xnor2_1 _19536_ (.Y(_09592_),
    .A(_09589_),
    .B(_09591_));
 sg13g2_nor2_1 _19537_ (.A(_09583_),
    .B(_09592_),
    .Y(_09593_));
 sg13g2_nand2_1 _19538_ (.Y(_09594_),
    .A(_09583_),
    .B(_09592_));
 sg13g2_o21ai_1 _19539_ (.B1(_09439_),
    .Y(_09595_),
    .A1(_09316_),
    .A2(_09546_));
 sg13g2_nand2b_1 _19540_ (.Y(_09596_),
    .B(_09595_),
    .A_N(_09547_));
 sg13g2_o21ai_1 _19541_ (.B1(_09594_),
    .Y(_09597_),
    .A1(_09593_),
    .A2(_09596_));
 sg13g2_inv_1 _19542_ (.Y(_09599_),
    .A(_09597_));
 sg13g2_xnor2_1 _19543_ (.Y(_09600_),
    .A(_09553_),
    .B(_09556_));
 sg13g2_xnor2_1 _19544_ (.Y(_09601_),
    .A(_09559_),
    .B(_09600_));
 sg13g2_nor2_1 _19545_ (.A(_09564_),
    .B(_09566_),
    .Y(_09602_));
 sg13g2_xnor2_1 _19546_ (.Y(_09603_),
    .A(_09568_),
    .B(_09602_));
 sg13g2_nand2_1 _19547_ (.Y(_09604_),
    .A(_09601_),
    .B(_09603_));
 sg13g2_nor2_1 _19548_ (.A(_09601_),
    .B(_09603_),
    .Y(_09605_));
 sg13g2_xor2_1 _19549_ (.B(_09603_),
    .A(_09601_),
    .X(_09606_));
 sg13g2_nor2b_1 _19550_ (.A(_09454_),
    .B_N(_09456_),
    .Y(_09607_));
 sg13g2_xnor2_1 _19551_ (.Y(_09608_),
    .A(_09462_),
    .B(_09607_));
 sg13g2_xnor2_1 _19552_ (.Y(_09610_),
    .A(_09606_),
    .B(_09608_));
 sg13g2_nand2b_1 _19553_ (.Y(_09611_),
    .B(_09594_),
    .A_N(_09593_));
 sg13g2_xnor2_1 _19554_ (.Y(_09612_),
    .A(_09596_),
    .B(_09611_));
 sg13g2_inv_1 _19555_ (.Y(_09613_),
    .A(_09612_));
 sg13g2_a21oi_1 _19556_ (.A1(_09604_),
    .A2(_09608_),
    .Y(_09614_),
    .B1(_09605_));
 sg13g2_o21ai_1 _19557_ (.B1(_09614_),
    .Y(_09615_),
    .A1(_09610_),
    .A2(_09613_));
 sg13g2_and3_1 _19558_ (.X(_09616_),
    .A(_09605_),
    .B(_09608_),
    .C(_09612_));
 sg13g2_inv_1 _19559_ (.Y(_09617_),
    .A(_09616_));
 sg13g2_a21oi_1 _19560_ (.A1(_09615_),
    .A2(_09617_),
    .Y(_09618_),
    .B1(_09599_));
 sg13g2_and3_1 _19561_ (.X(_09619_),
    .A(_09599_),
    .B(_09615_),
    .C(_09617_));
 sg13g2_o21ai_1 _19562_ (.B1(_09574_),
    .Y(_09621_),
    .A1(_09618_),
    .A2(_09619_));
 sg13g2_nor3_1 _19563_ (.A(_09574_),
    .B(_09618_),
    .C(_09619_),
    .Y(_09622_));
 sg13g2_or3_1 _19564_ (.A(_09574_),
    .B(_09618_),
    .C(_09619_),
    .X(_09623_));
 sg13g2_o21ai_1 _19565_ (.B1(_09579_),
    .Y(_09624_),
    .A1(_09578_),
    .A2(_09582_));
 sg13g2_nand3_1 _19566_ (.B(_09623_),
    .C(_09624_),
    .A(_09621_),
    .Y(_09625_));
 sg13g2_a21o_1 _19567_ (.A2(_09623_),
    .A1(_09621_),
    .B1(_09624_),
    .X(_09626_));
 sg13g2_nand2_1 _19568_ (.Y(_09627_),
    .A(_09588_),
    .B(_09591_));
 sg13g2_nand2_1 _19569_ (.Y(_09628_),
    .A(_09586_),
    .B(_09627_));
 sg13g2_inv_1 _19570_ (.Y(_09629_),
    .A(_09628_));
 sg13g2_nand3_1 _19571_ (.B(_09626_),
    .C(_09629_),
    .A(_09625_),
    .Y(_09630_));
 sg13g2_a21o_1 _19572_ (.A2(_09626_),
    .A1(_09625_),
    .B1(_09629_),
    .X(_09632_));
 sg13g2_nand2_2 _19573_ (.Y(_09633_),
    .A(_09630_),
    .B(_09632_));
 sg13g2_inv_1 _19574_ (.Y(_09634_),
    .A(_09633_));
 sg13g2_xnor2_1 _19575_ (.Y(_09635_),
    .A(_08668_),
    .B(_08681_));
 sg13g2_nand3_1 _19576_ (.B(_08631_),
    .C(_08633_),
    .A(_08629_),
    .Y(_09636_));
 sg13g2_nand2b_2 _19577_ (.Y(_09637_),
    .B(_09636_),
    .A_N(_08634_));
 sg13g2_inv_1 _19578_ (.Y(_09638_),
    .A(_09637_));
 sg13g2_xnor2_1 _19579_ (.Y(_09639_),
    .A(_08595_),
    .B(_08602_));
 sg13g2_inv_1 _19580_ (.Y(_09640_),
    .A(_09639_));
 sg13g2_xnor2_1 _19581_ (.Y(_09641_),
    .A(_08827_),
    .B(_09447_));
 sg13g2_inv_1 _19582_ (.Y(_09643_),
    .A(_09641_));
 sg13g2_xor2_1 _19583_ (.B(_08436_),
    .A(_08425_),
    .X(_09644_));
 sg13g2_inv_1 _19584_ (.Y(_09645_),
    .A(_09644_));
 sg13g2_xnor2_1 _19585_ (.Y(_09646_),
    .A(_08898_),
    .B(_09223_));
 sg13g2_nor2_1 _19586_ (.A(_09644_),
    .B(_09646_),
    .Y(_09647_));
 sg13g2_a21oi_1 _19587_ (.A1(_09640_),
    .A2(_09641_),
    .Y(_09648_),
    .B1(_09647_));
 sg13g2_a21oi_1 _19588_ (.A1(_09639_),
    .A2(_09643_),
    .Y(_09649_),
    .B1(_09648_));
 sg13g2_nand2_1 _19589_ (.Y(_09650_),
    .A(_09637_),
    .B(_09649_));
 sg13g2_nor2_1 _19590_ (.A(_09637_),
    .B(_09649_),
    .Y(_09651_));
 sg13g2_nand3_1 _19591_ (.B(_09541_),
    .C(_09552_),
    .A(_09540_),
    .Y(_09652_));
 sg13g2_nand2b_2 _19592_ (.Y(_09654_),
    .B(_09652_),
    .A_N(_09553_));
 sg13g2_inv_1 _19593_ (.Y(_09655_),
    .A(_09654_));
 sg13g2_a21oi_1 _19594_ (.A1(_09650_),
    .A2(_09654_),
    .Y(_09656_),
    .B1(_09651_));
 sg13g2_xnor2_1 _19595_ (.Y(_09657_),
    .A(_09610_),
    .B(_09612_));
 sg13g2_inv_1 _19596_ (.Y(_09658_),
    .A(_09657_));
 sg13g2_a21o_1 _19597_ (.A2(_09657_),
    .A1(_09635_),
    .B1(_09656_),
    .X(_09659_));
 sg13g2_nor2_1 _19598_ (.A(_09635_),
    .B(_09657_),
    .Y(_09660_));
 sg13g2_a21oi_1 _19599_ (.A1(_08703_),
    .A2(_09633_),
    .Y(_09661_),
    .B1(_09660_));
 sg13g2_a22oi_1 _19600_ (.Y(_09662_),
    .B1(_09659_),
    .B2(_09661_),
    .A2(_09634_),
    .A1(_08704_));
 sg13g2_a21oi_2 _19601_ (.B1(_09622_),
    .Y(_09663_),
    .A2(_09624_),
    .A1(_09621_));
 sg13g2_xor2_1 _19602_ (.B(_09663_),
    .A(_09630_),
    .X(_09665_));
 sg13g2_a21oi_1 _19603_ (.A1(_09599_),
    .A2(_09615_),
    .Y(_09666_),
    .B1(_09616_));
 sg13g2_a21o_1 _19604_ (.A2(_09663_),
    .A1(_09630_),
    .B1(_09666_),
    .X(_09667_));
 sg13g2_xnor2_1 _19605_ (.Y(_09668_),
    .A(_09665_),
    .B(_09666_));
 sg13g2_nor2_1 _19606_ (.A(_09463_),
    .B(_09571_),
    .Y(_09669_));
 sg13g2_or2_2 _19607_ (.X(_09670_),
    .B(_09669_),
    .A(_09572_));
 sg13g2_inv_1 _19608_ (.Y(_09671_),
    .A(_09670_));
 sg13g2_xnor2_1 _19609_ (.Y(_09672_),
    .A(_09668_),
    .B(_09671_));
 sg13g2_inv_1 _19610_ (.Y(_09673_),
    .A(_09672_));
 sg13g2_o21ai_1 _19611_ (.B1(_08698_),
    .Y(_09674_),
    .A1(_08473_),
    .A2(_08695_));
 sg13g2_nor3_1 _19612_ (.A(_08082_),
    .B(_08473_),
    .C(_08698_),
    .Y(_09676_));
 sg13g2_a21o_1 _19613_ (.A2(_08701_),
    .A1(_08083_),
    .B1(_09674_),
    .X(_09677_));
 sg13g2_xnor2_1 _19614_ (.Y(_09678_),
    .A(_08702_),
    .B(_09674_));
 sg13g2_a21oi_1 _19615_ (.A1(_08687_),
    .A2(_08689_),
    .Y(_09679_),
    .B1(_08684_));
 sg13g2_xnor2_1 _19616_ (.Y(_09680_),
    .A(_09678_),
    .B(_09679_));
 sg13g2_a21oi_2 _19617_ (.B1(_08645_),
    .Y(_09681_),
    .A2(_08654_),
    .A1(_08644_));
 sg13g2_xor2_1 _19618_ (.B(_09681_),
    .A(_09680_),
    .X(_09682_));
 sg13g2_a21oi_1 _19619_ (.A1(_09677_),
    .A2(_09679_),
    .Y(_09683_),
    .B1(_09676_));
 sg13g2_o21ai_1 _19620_ (.B1(_09683_),
    .Y(_09684_),
    .A1(_09680_),
    .A2(_09681_));
 sg13g2_inv_1 _19621_ (.Y(_09685_),
    .A(_09684_));
 sg13g2_o21ai_1 _19622_ (.B1(_09667_),
    .Y(_09687_),
    .A1(_09630_),
    .A2(_09663_));
 sg13g2_a21oi_1 _19623_ (.A1(_09668_),
    .A2(_09671_),
    .Y(_09688_),
    .B1(_09687_));
 sg13g2_a21o_1 _19624_ (.A2(_09671_),
    .A1(_09668_),
    .B1(_09687_),
    .X(_09689_));
 sg13g2_o21ai_1 _19625_ (.B1(_09682_),
    .Y(_09690_),
    .A1(_09662_),
    .A2(_09672_));
 sg13g2_a22oi_1 _19626_ (.Y(_09691_),
    .B1(_09684_),
    .B2(_09688_),
    .A2(_09672_),
    .A1(_09662_));
 sg13g2_a22oi_1 _19627_ (.Y(_09692_),
    .B1(_09690_),
    .B2(_09691_),
    .A2(_09689_),
    .A1(_09685_));
 sg13g2_mux2_2 _19628_ (.A0(_09633_),
    .A1(_08704_),
    .S(net2168),
    .X(_09693_));
 sg13g2_a21o_1 _19629_ (.A2(net2169),
    .A1(net2172),
    .B1(_07687_),
    .X(_09694_));
 sg13g2_nand3_1 _19630_ (.B(_07688_),
    .C(net2170),
    .A(net2172),
    .Y(_09695_));
 sg13g2_nand2_1 _19631_ (.Y(_09696_),
    .A(_09694_),
    .B(_09695_));
 sg13g2_a21oi_1 _19632_ (.A1(_09694_),
    .A2(_09695_),
    .Y(_09698_),
    .B1(_09693_));
 sg13g2_mux2_2 _19633_ (.A0(_09673_),
    .A1(_09682_),
    .S(net2168),
    .X(_09699_));
 sg13g2_nand3b_1 _19634_ (.B(net2170),
    .C(net2172),
    .Y(_09700_),
    .A_N(_07711_));
 sg13g2_a21o_1 _19635_ (.A2(net2170),
    .A1(net2172),
    .B1(_07686_),
    .X(_09701_));
 sg13g2_and2_1 _19636_ (.A(_09700_),
    .B(_09701_),
    .X(_09702_));
 sg13g2_inv_1 _19637_ (.Y(_09703_),
    .A(_09702_));
 sg13g2_and3_1 _19638_ (.X(_09704_),
    .A(_09699_),
    .B(_09700_),
    .C(_09701_));
 sg13g2_or2_1 _19639_ (.X(_09705_),
    .B(_09704_),
    .A(_09698_));
 sg13g2_and3_1 _19640_ (.X(_09706_),
    .A(_09693_),
    .B(_09694_),
    .C(_09695_));
 sg13g2_a21oi_1 _19641_ (.A1(_09700_),
    .A2(_09701_),
    .Y(_09707_),
    .B1(_09699_));
 sg13g2_or2_1 _19642_ (.X(_09709_),
    .B(_09702_),
    .A(_09699_));
 sg13g2_nor4_2 _19643_ (.A(_09698_),
    .B(_09704_),
    .C(_09706_),
    .Y(_09710_),
    .D(_09707_));
 sg13g2_a21o_1 _19644_ (.A2(net2169),
    .A1(net2171),
    .B1(_07703_),
    .X(_09711_));
 sg13g2_nand3_1 _19645_ (.B(_07693_),
    .C(net2169),
    .A(net2171),
    .Y(_09712_));
 sg13g2_mux2_1 _19646_ (.A0(_09655_),
    .A1(_09638_),
    .S(net2168),
    .X(_09713_));
 sg13g2_nand3_1 _19647_ (.B(_09712_),
    .C(_09713_),
    .A(_09711_),
    .Y(_09714_));
 sg13g2_mux2_1 _19648_ (.A0(_09658_),
    .A1(_09635_),
    .S(net2168),
    .X(_09715_));
 sg13g2_a21o_1 _19649_ (.A2(net2169),
    .A1(net2171),
    .B1(_07691_),
    .X(_09716_));
 sg13g2_nand3_1 _19650_ (.B(_07689_),
    .C(net2169),
    .A(net2171),
    .Y(_09717_));
 sg13g2_nand2_1 _19651_ (.Y(_09718_),
    .A(_09716_),
    .B(_09717_));
 sg13g2_a21o_1 _19652_ (.A2(_09717_),
    .A1(_09716_),
    .B1(_09715_),
    .X(_09720_));
 sg13g2_a21o_1 _19653_ (.A2(_09712_),
    .A1(_09711_),
    .B1(_09713_),
    .X(_09721_));
 sg13g2_and3_1 _19654_ (.X(_09722_),
    .A(_09715_),
    .B(_09716_),
    .C(_09717_));
 sg13g2_nand3_1 _19655_ (.B(_09716_),
    .C(_09717_),
    .A(_09715_),
    .Y(_09723_));
 sg13g2_and4_1 _19656_ (.A(_09714_),
    .B(_09720_),
    .C(_09721_),
    .D(_09723_),
    .X(_09724_));
 sg13g2_a21oi_1 _19657_ (.A1(net2171),
    .A2(net2169),
    .Y(_09725_),
    .B1(_07696_));
 sg13g2_o21ai_1 _19658_ (.B1(_07694_),
    .Y(_09726_),
    .A1(_07682_),
    .A2(_07718_));
 sg13g2_nor3_1 _19659_ (.A(_07682_),
    .B(_07698_),
    .C(_07718_),
    .Y(_09727_));
 sg13g2_nand3_1 _19660_ (.B(_07697_),
    .C(net2169),
    .A(net2171),
    .Y(_09728_));
 sg13g2_nand2_1 _19661_ (.Y(_09729_),
    .A(_09726_),
    .B(_09728_));
 sg13g2_mux2_1 _19662_ (.A0(_09643_),
    .A1(_09640_),
    .S(net2168),
    .X(_09731_));
 sg13g2_mux2_1 _19663_ (.A0(_09641_),
    .A1(_09639_),
    .S(_09692_),
    .X(_09732_));
 sg13g2_a21oi_1 _19664_ (.A1(_09726_),
    .A2(_09728_),
    .Y(_09733_),
    .B1(_09731_));
 sg13g2_o21ai_1 _19665_ (.B1(_09732_),
    .Y(_09734_),
    .A1(_09725_),
    .A2(_09727_));
 sg13g2_nor3_1 _19666_ (.A(_09725_),
    .B(_09727_),
    .C(_09732_),
    .Y(_09735_));
 sg13g2_nand2_1 _19667_ (.Y(_09736_),
    .A(_09644_),
    .B(net2168));
 sg13g2_mux2_1 _19668_ (.A0(_09646_),
    .A1(_09645_),
    .S(net2168),
    .X(_09737_));
 sg13g2_o21ai_1 _19669_ (.B1(_09736_),
    .Y(_09738_),
    .A1(_09646_),
    .A2(net2168));
 sg13g2_and3_1 _19670_ (.X(_09739_),
    .A(_07721_),
    .B(_07722_),
    .C(_09737_));
 sg13g2_nor3_1 _19671_ (.A(_09733_),
    .B(_09735_),
    .C(_09739_),
    .Y(_09740_));
 sg13g2_o21ai_1 _19672_ (.B1(_09734_),
    .Y(_09742_),
    .A1(_09735_),
    .A2(_09739_));
 sg13g2_a21oi_1 _19673_ (.A1(_09714_),
    .A2(_09720_),
    .Y(_09743_),
    .B1(_09722_));
 sg13g2_a21o_1 _19674_ (.A2(_09742_),
    .A1(_09724_),
    .B1(_09743_),
    .X(_09744_));
 sg13g2_nor2_1 _19675_ (.A(_07272_),
    .B(net9),
    .Y(_09745_));
 sg13g2_nor2_2 _19676_ (.A(_09684_),
    .B(_09689_),
    .Y(_09746_));
 sg13g2_nor3_1 _19677_ (.A(_07272_),
    .B(net9),
    .C(_09746_),
    .Y(_09747_));
 sg13g2_a21o_1 _19678_ (.A2(_09709_),
    .A1(_09705_),
    .B1(_09747_),
    .X(_09748_));
 sg13g2_a21oi_2 _19679_ (.B1(_09748_),
    .Y(_09749_),
    .A2(_09744_),
    .A1(_09710_));
 sg13g2_a21o_1 _19680_ (.A2(_09744_),
    .A1(_09710_),
    .B1(_09748_),
    .X(_09750_));
 sg13g2_o21ai_1 _19681_ (.B1(_09746_),
    .Y(_09751_),
    .A1(_07272_),
    .A2(net9));
 sg13g2_a21oi_1 _19682_ (.A1(_07723_),
    .A2(_09738_),
    .Y(_09753_),
    .B1(_09747_));
 sg13g2_nand4_1 _19683_ (.B(_09724_),
    .C(_09740_),
    .A(_09710_),
    .Y(_09754_),
    .D(_09753_));
 sg13g2_and2_1 _19684_ (.A(_09751_),
    .B(_09754_),
    .X(_09755_));
 sg13g2_nand2_1 _19685_ (.Y(_09756_),
    .A(_09751_),
    .B(_09754_));
 sg13g2_nor2_2 _19686_ (.A(_09749_),
    .B(_09756_),
    .Y(_09757_));
 sg13g2_inv_1 _19687_ (.Y(_09758_),
    .A(_09757_));
 sg13g2_o21ai_1 _19688_ (.B1(_07723_),
    .Y(_09759_),
    .A1(_09749_),
    .A2(_09756_));
 sg13g2_nand3_1 _19689_ (.B(_09750_),
    .C(_09755_),
    .A(_09737_),
    .Y(_09760_));
 sg13g2_and2_1 _19690_ (.A(_09759_),
    .B(_09760_),
    .X(_09761_));
 sg13g2_nand3_1 _19691_ (.B(_09759_),
    .C(_09760_),
    .A(_05719_),
    .Y(_09762_));
 sg13g2_o21ai_1 _19692_ (.B1(_09729_),
    .Y(_09764_),
    .A1(_09749_),
    .A2(_09756_));
 sg13g2_nand3_1 _19693_ (.B(_09750_),
    .C(_09755_),
    .A(_09731_),
    .Y(_09765_));
 sg13g2_nand2_1 _19694_ (.Y(_09766_),
    .A(_09764_),
    .B(_09765_));
 sg13g2_mux2_2 _19695_ (.A0(_05688_),
    .A1(_05692_),
    .S(_05714_),
    .X(_09767_));
 sg13g2_nand3_1 _19696_ (.B(_09765_),
    .C(_09767_),
    .A(_09764_),
    .Y(_09768_));
 sg13g2_and3_1 _19697_ (.X(_09769_),
    .A(_09713_),
    .B(_09750_),
    .C(_09755_));
 sg13g2_a22oi_1 _19698_ (.Y(_09770_),
    .B1(_09750_),
    .B2(_09755_),
    .A2(_09712_),
    .A1(_09711_));
 sg13g2_nor2_1 _19699_ (.A(_09769_),
    .B(_09770_),
    .Y(_09771_));
 sg13g2_mux2_2 _19700_ (.A0(_05677_),
    .A1(_05674_),
    .S(_05714_),
    .X(_09772_));
 sg13g2_inv_1 _19701_ (.Y(_09773_),
    .A(_09772_));
 sg13g2_a21oi_1 _19702_ (.A1(_09764_),
    .A2(_09765_),
    .Y(_09775_),
    .B1(_09767_));
 sg13g2_a221oi_1 _19703_ (.B2(_09773_),
    .C1(_09775_),
    .B1(_09771_),
    .A1(_09762_),
    .Y(_09776_),
    .A2(_09768_));
 sg13g2_o21ai_1 _19704_ (.B1(_09772_),
    .Y(_09777_),
    .A1(_09769_),
    .A2(_09770_));
 sg13g2_mux2_2 _19705_ (.A0(_09718_),
    .A1(_09715_),
    .S(_09757_),
    .X(_09778_));
 sg13g2_mux2_2 _19706_ (.A0(_05672_),
    .A1(_05669_),
    .S(_05714_),
    .X(_09779_));
 sg13g2_inv_1 _19707_ (.Y(_09780_),
    .A(_09779_));
 sg13g2_o21ai_1 _19708_ (.B1(_09777_),
    .Y(_09781_),
    .A1(_09778_),
    .A2(_09780_));
 sg13g2_mux2_2 _19709_ (.A0(_09696_),
    .A1(_09693_),
    .S(_09757_),
    .X(_09782_));
 sg13g2_inv_1 _19710_ (.Y(_09783_),
    .A(_09782_));
 sg13g2_mux2_2 _19711_ (.A0(_05657_),
    .A1(_05662_),
    .S(_05714_),
    .X(_09784_));
 sg13g2_inv_1 _19712_ (.Y(_09786_),
    .A(_09784_));
 sg13g2_a22oi_1 _19713_ (.Y(_09787_),
    .B1(_09782_),
    .B2(_09786_),
    .A2(_09780_),
    .A1(_09778_));
 sg13g2_o21ai_1 _19714_ (.B1(_09787_),
    .Y(_09788_),
    .A1(_09776_),
    .A2(_09781_));
 sg13g2_mux2_2 _19715_ (.A0(_09703_),
    .A1(_09699_),
    .S(_09757_),
    .X(_09789_));
 sg13g2_inv_1 _19716_ (.Y(_09790_),
    .A(_09789_));
 sg13g2_mux2_2 _19717_ (.A0(_05651_),
    .A1(_05645_),
    .S(_05714_),
    .X(_09791_));
 sg13g2_inv_1 _19718_ (.Y(_09792_),
    .A(_09791_));
 sg13g2_a22oi_1 _19719_ (.Y(_09793_),
    .B1(_09789_),
    .B2(_09791_),
    .A2(_09784_),
    .A1(_09783_));
 sg13g2_nand2_1 _19720_ (.Y(_09794_),
    .A(_09745_),
    .B(_09746_));
 sg13g2_nand2b_2 _19721_ (.Y(_09795_),
    .B(_05706_),
    .A_N(_05705_));
 sg13g2_nand3_1 _19722_ (.B(_09746_),
    .C(_09795_),
    .A(_09745_),
    .Y(_09797_));
 sg13g2_o21ai_1 _19723_ (.B1(_09797_),
    .Y(_09798_),
    .A1(_09789_),
    .A2(_09791_));
 sg13g2_a21o_1 _19724_ (.A2(_09793_),
    .A1(_09788_),
    .B1(_09798_),
    .X(_09799_));
 sg13g2_nand2b_1 _19725_ (.Y(_09800_),
    .B(_09794_),
    .A_N(_09795_));
 sg13g2_and2_1 _19726_ (.A(_09799_),
    .B(_09800_),
    .X(_09801_));
 sg13g2_nand3_1 _19727_ (.B(_09759_),
    .C(_09760_),
    .A(_01962_),
    .Y(_09802_));
 sg13g2_mux2_2 _19728_ (.A0(_01938_),
    .A1(_01937_),
    .S(_01960_),
    .X(_09803_));
 sg13g2_inv_1 _19729_ (.Y(_09804_),
    .A(_09803_));
 sg13g2_nand3_1 _19730_ (.B(_09765_),
    .C(_09803_),
    .A(_09764_),
    .Y(_09805_));
 sg13g2_a21oi_1 _19731_ (.A1(_09764_),
    .A2(_09765_),
    .Y(_09806_),
    .B1(_09803_));
 sg13g2_mux2_2 _19732_ (.A0(_01943_),
    .A1(_01942_),
    .S(_01960_),
    .X(_09808_));
 sg13g2_inv_1 _19733_ (.Y(_09809_),
    .A(_09808_));
 sg13g2_a221oi_1 _19734_ (.B2(_09771_),
    .C1(_09806_),
    .B1(_09809_),
    .A1(_09802_),
    .Y(_09810_),
    .A2(_09805_));
 sg13g2_o21ai_1 _19735_ (.B1(_09808_),
    .Y(_09811_),
    .A1(_09769_),
    .A2(_09770_));
 sg13g2_mux2_2 _19736_ (.A0(_01934_),
    .A1(_01933_),
    .S(_01960_),
    .X(_09812_));
 sg13g2_o21ai_1 _19737_ (.B1(_09811_),
    .Y(_09813_),
    .A1(_09778_),
    .A2(_09812_));
 sg13g2_mux2_2 _19738_ (.A0(_01951_),
    .A1(_01950_),
    .S(_01960_),
    .X(_09814_));
 sg13g2_inv_1 _19739_ (.Y(_09815_),
    .A(_09814_));
 sg13g2_a22oi_1 _19740_ (.Y(_09816_),
    .B1(_09815_),
    .B2(_09782_),
    .A2(_09812_),
    .A1(_09778_));
 sg13g2_o21ai_1 _19741_ (.B1(_09816_),
    .Y(_09817_),
    .A1(_09810_),
    .A2(_09813_));
 sg13g2_mux2_2 _19742_ (.A0(_01931_),
    .A1(_01932_),
    .S(_01960_),
    .X(_09819_));
 sg13g2_inv_1 _19743_ (.Y(_09820_),
    .A(_09819_));
 sg13g2_a22oi_1 _19744_ (.Y(_09821_),
    .B1(_09819_),
    .B2(_09789_),
    .A2(_09814_),
    .A1(_09783_));
 sg13g2_nor2_2 _19745_ (.A(_01548_),
    .B(_01930_),
    .Y(_09822_));
 sg13g2_or2_1 _19746_ (.X(_09823_),
    .B(_09822_),
    .A(_09794_));
 sg13g2_o21ai_1 _19747_ (.B1(_09823_),
    .Y(_09824_),
    .A1(_09789_),
    .A2(_09819_));
 sg13g2_a21o_1 _19748_ (.A2(_09821_),
    .A1(_09817_),
    .B1(_09824_),
    .X(_09825_));
 sg13g2_nand2_1 _19749_ (.Y(_09826_),
    .A(_09794_),
    .B(_09822_));
 sg13g2_a22oi_1 _19750_ (.Y(_09827_),
    .B1(_09825_),
    .B2(_09826_),
    .A2(_09800_),
    .A1(_09799_));
 sg13g2_nand3b_1 _19751_ (.B(_05718_),
    .C(_01962_),
    .Y(_09828_),
    .A_N(_05717_));
 sg13g2_o21ai_1 _19752_ (.B1(_09828_),
    .Y(_09830_),
    .A1(_09767_),
    .A2(_09804_));
 sg13g2_a22oi_1 _19753_ (.Y(_09831_),
    .B1(_09809_),
    .B2(_09772_),
    .A2(_09804_),
    .A1(_09767_));
 sg13g2_nor2_1 _19754_ (.A(_09779_),
    .B(_09812_),
    .Y(_09832_));
 sg13g2_a221oi_1 _19755_ (.B2(_09831_),
    .C1(_09832_),
    .B1(_09830_),
    .A1(_09773_),
    .Y(_09833_),
    .A2(_09808_));
 sg13g2_a22oi_1 _19756_ (.Y(_09834_),
    .B1(_09815_),
    .B2(_09784_),
    .A2(_09812_),
    .A1(_09779_));
 sg13g2_inv_1 _19757_ (.Y(_09835_),
    .A(_09834_));
 sg13g2_a22oi_1 _19758_ (.Y(_09836_),
    .B1(_09819_),
    .B2(_09792_),
    .A2(_09814_),
    .A1(_09786_));
 sg13g2_o21ai_1 _19759_ (.B1(_09836_),
    .Y(_09837_),
    .A1(_09833_),
    .A2(_09835_));
 sg13g2_nor2_1 _19760_ (.A(_09795_),
    .B(_09822_),
    .Y(_09838_));
 sg13g2_a21oi_1 _19761_ (.A1(_09791_),
    .A2(_09820_),
    .Y(_09839_),
    .B1(_09838_));
 sg13g2_and2_1 _19762_ (.A(_09795_),
    .B(_09822_),
    .X(_09841_));
 sg13g2_a21oi_1 _19763_ (.A1(_09837_),
    .A2(_09839_),
    .Y(_09842_),
    .B1(_09841_));
 sg13g2_a21o_1 _19764_ (.A2(_09839_),
    .A1(_09837_),
    .B1(_09841_),
    .X(_09843_));
 sg13g2_and2_2 _19765_ (.A(_09801_),
    .B(_09843_),
    .X(_09844_));
 sg13g2_nand3_1 _19766_ (.B(_09800_),
    .C(_09843_),
    .A(_09799_),
    .Y(_09845_));
 sg13g2_nor2_2 _19767_ (.A(net2167),
    .B(_09844_),
    .Y(_09846_));
 sg13g2_inv_1 _19768_ (.Y(_09847_),
    .A(_09846_));
 sg13g2_a22oi_1 _19769_ (.Y(_09848_),
    .B1(_09844_),
    .B2(_05720_),
    .A2(net2166),
    .A1(_09761_));
 sg13g2_o21ai_1 _19770_ (.B1(_09848_),
    .Y(uio_out[0]),
    .A1(_01962_),
    .A2(_09847_));
 sg13g2_nor2b_1 _19771_ (.A(_09845_),
    .B_N(_09767_),
    .Y(_09849_));
 sg13g2_a221oi_1 _19772_ (.B2(_09803_),
    .C1(_09849_),
    .B1(_09846_),
    .A1(_09766_),
    .Y(uio_out[1]),
    .A2(net2166));
 sg13g2_nor2_1 _19773_ (.A(_09773_),
    .B(_09845_),
    .Y(_09851_));
 sg13g2_a221oi_1 _19774_ (.B2(_09808_),
    .C1(_09851_),
    .B1(_09846_),
    .A1(_09771_),
    .Y(uio_out[2]),
    .A2(net2166));
 sg13g2_nor3_1 _19775_ (.A(_09812_),
    .B(net2166),
    .C(_09844_),
    .Y(_09852_));
 sg13g2_a221oi_1 _19776_ (.B2(_09779_),
    .C1(_09852_),
    .B1(_09844_),
    .A1(_09778_),
    .Y(uio_out[3]),
    .A2(net2166));
 sg13g2_nor2_1 _19777_ (.A(_09786_),
    .B(_09845_),
    .Y(_09853_));
 sg13g2_a221oi_1 _19778_ (.B2(_09814_),
    .C1(_09853_),
    .B1(_09846_),
    .A1(_09782_),
    .Y(uio_out[4]),
    .A2(net2166));
 sg13g2_nor2_1 _19779_ (.A(_09792_),
    .B(_09845_),
    .Y(_09854_));
 sg13g2_a221oi_1 _19780_ (.B2(_09819_),
    .C1(_09854_),
    .B1(_09846_),
    .A1(_09790_),
    .Y(uio_out[5]),
    .A2(net2166));
 sg13g2_or4_2 _19781_ (.A(_01548_),
    .B(_01930_),
    .C(_09794_),
    .D(_09795_),
    .X(uio_out[6]));
 sg13g2_mux2_1 _19782_ (.A0(_07720_),
    .A1(_09692_),
    .S(_09757_),
    .X(_09856_));
 sg13g2_nor2b_1 _19783_ (.A(_09856_),
    .B_N(net2167),
    .Y(_09857_));
 sg13g2_nor2_1 _19784_ (.A(_03802_),
    .B(_05714_),
    .Y(_09858_));
 sg13g2_a21oi_2 _19785_ (.B1(_09858_),
    .Y(_09859_),
    .A2(_05714_),
    .A1(_05641_));
 sg13g2_nor2_1 _19786_ (.A(_09842_),
    .B(_09859_),
    .Y(_09860_));
 sg13g2_a221oi_1 _19787_ (.B2(_09801_),
    .C1(net2166),
    .B1(_09860_),
    .A1(_01961_),
    .Y(_09861_),
    .A2(_09845_));
 sg13g2_nor2_1 _19788_ (.A(_09857_),
    .B(_09861_),
    .Y(_09862_));
 sg13g2_or2_1 _19789_ (.X(_09863_),
    .B(_09861_),
    .A(_09857_));
 sg13g2_o21ai_1 _19790_ (.B1(_09845_),
    .Y(_09864_),
    .A1(_09857_),
    .A2(_09861_));
 sg13g2_nand2_1 _19791_ (.Y(_09865_),
    .A(_09758_),
    .B(net2167));
 sg13g2_and2_1 _19792_ (.A(_09864_),
    .B(_09865_),
    .X(_00280_));
 sg13g2_o21ai_1 _19793_ (.B1(_00280_),
    .Y(uo_out[0]),
    .A1(net2167),
    .A2(_09861_));
 sg13g2_a22oi_1 _19794_ (.Y(_00281_),
    .B1(_09844_),
    .B2(_05716_),
    .A2(net2167),
    .A1(_09758_));
 sg13g2_and2_1 _19795_ (.A(_09863_),
    .B(_00281_),
    .X(_00282_));
 sg13g2_o21ai_1 _19796_ (.B1(_09844_),
    .Y(_00283_),
    .A1(_09863_),
    .A2(_00281_));
 sg13g2_or2_1 _19797_ (.X(uo_out[1]),
    .B(_00283_),
    .A(_00282_));
 sg13g2_nand2b_1 _19798_ (.Y(uo_out[2]),
    .B(_09857_),
    .A_N(_00281_));
 sg13g2_o21ai_1 _19799_ (.B1(_00280_),
    .Y(uo_out[3]),
    .A1(_00282_),
    .A2(_00283_));
 sg13g2_a21oi_1 _19800_ (.A1(_09844_),
    .A2(_00281_),
    .Y(uo_out[4]),
    .B1(_09862_));
 sg13g2_nand2b_1 _19801_ (.Y(_00284_),
    .B(_09865_),
    .A_N(_09864_));
 sg13g2_nand3_1 _19802_ (.B(_00283_),
    .C(_00284_),
    .A(_09847_),
    .Y(uo_out[5]));
 sg13g2_nand3_1 _19803_ (.B(_09865_),
    .C(_00283_),
    .A(_09847_),
    .Y(uo_out[6]));
 sg13g2_mux2_1 _19804_ (.A0(net1),
    .A1(net292),
    .S(net2845),
    .X(_00025_));
 sg13g2_mux2_1 _19805_ (.A0(net2),
    .A1(net294),
    .S(net2846),
    .X(_00026_));
 sg13g2_mux2_1 _19806_ (.A0(net3),
    .A1(net279),
    .S(net2849),
    .X(_00027_));
 sg13g2_mux2_1 _19807_ (.A0(net4),
    .A1(net299),
    .S(net2845),
    .X(_00028_));
 sg13g2_mux2_1 _19808_ (.A0(net5),
    .A1(\net.in[4] ),
    .S(net2849),
    .X(_00029_));
 sg13g2_mux2_1 _19809_ (.A0(net6),
    .A1(net2817),
    .S(net2845),
    .X(_00030_));
 sg13g2_mux2_1 _19810_ (.A0(net7),
    .A1(net2814),
    .S(net2844),
    .X(_00031_));
 sg13g2_nor2_1 _19811_ (.A(net2844),
    .B(net8),
    .Y(_00286_));
 sg13g2_a21oi_1 _19812_ (.A1(_06045_),
    .A2(net2844),
    .Y(_00032_),
    .B1(_00286_));
 sg13g2_mux2_1 _19813_ (.A0(net292),
    .A1(net2809),
    .S(net2845),
    .X(_00033_));
 sg13g2_mux2_1 _19814_ (.A0(net294),
    .A1(net2807),
    .S(net2846),
    .X(_00034_));
 sg13g2_nor2_1 _19815_ (.A(net2849),
    .B(net279),
    .Y(_00288_));
 sg13g2_a21oi_1 _19816_ (.A1(_05506_),
    .A2(net2849),
    .Y(_00035_),
    .B1(_00288_));
 sg13g2_nor2_1 _19817_ (.A(net2844),
    .B(net299),
    .Y(_00289_));
 sg13g2_a21oi_1 _19818_ (.A1(_05154_),
    .A2(net2847),
    .Y(_00036_),
    .B1(_00289_));
 sg13g2_mux2_1 _19819_ (.A0(\net.in[4] ),
    .A1(net2804),
    .S(net2849),
    .X(_00037_));
 sg13g2_mux2_1 _19820_ (.A0(net2817),
    .A1(net380),
    .S(net2886),
    .X(_00038_));
 sg13g2_mux2_1 _19821_ (.A0(net2814),
    .A1(net290),
    .S(net2844),
    .X(_00039_));
 sg13g2_nand2_1 _19822_ (.Y(_00291_),
    .A(net2844),
    .B(net286));
 sg13g2_o21ai_1 _19823_ (.B1(_00291_),
    .Y(_00040_),
    .A1(_06045_),
    .A2(net2844));
 sg13g2_mux2_1 _19824_ (.A0(net2811),
    .A1(net273),
    .S(net2846),
    .X(_00041_));
 sg13g2_mux2_1 _19825_ (.A0(net2807),
    .A1(net295),
    .S(net2818),
    .X(_00042_));
 sg13g2_nand2_1 _19826_ (.Y(_00292_),
    .A(net280),
    .B(net2877));
 sg13g2_o21ai_1 _19827_ (.B1(_00292_),
    .Y(_00043_),
    .A1(_05506_),
    .A2(net2877));
 sg13g2_nand2_1 _19828_ (.Y(_00293_),
    .A(net2802),
    .B(net2878));
 sg13g2_o21ai_1 _19829_ (.B1(_00293_),
    .Y(_00044_),
    .A1(_05154_),
    .A2(net2878));
 sg13g2_mux2_1 _19830_ (.A0(net2804),
    .A1(net2801),
    .S(net2849),
    .X(_00045_));
 sg13g2_mux2_1 _19831_ (.A0(net380),
    .A1(net2798),
    .S(net2886),
    .X(_00046_));
 sg13g2_mux2_1 _19832_ (.A0(net290),
    .A1(net2796),
    .S(net2844),
    .X(_00047_));
 sg13g2_mux2_1 _19833_ (.A0(net286),
    .A1(net2793),
    .S(net2847),
    .X(_00048_));
 sg13g2_nor2_1 _19834_ (.A(net2846),
    .B(net273),
    .Y(_00295_));
 sg13g2_a21oi_1 _19835_ (.A1(_05913_),
    .A2(net2839),
    .Y(_00049_),
    .B1(_00295_));
 sg13g2_mux2_1 _19836_ (.A0(net295),
    .A1(net2787),
    .S(net2818),
    .X(_00050_));
 sg13g2_nor2_1 _19837_ (.A(net280),
    .B(net2872),
    .Y(_00296_));
 sg13g2_a21oi_1 _19838_ (.A1(_05869_),
    .A2(net2872),
    .Y(_00051_),
    .B1(_00296_));
 sg13g2_mux2_1 _19839_ (.A0(net2802),
    .A1(net2783),
    .S(net2870),
    .X(_00052_));
 sg13g2_mux2_1 _19840_ (.A0(net2801),
    .A1(net2779),
    .S(net2849),
    .X(_00053_));
 sg13g2_mux2_1 _19841_ (.A0(net2799),
    .A1(net2776),
    .S(net2823),
    .X(_00054_));
 sg13g2_mux2_1 _19842_ (.A0(net2795),
    .A1(net2775),
    .S(net2885),
    .X(_00055_));
 sg13g2_mux2_1 _19843_ (.A0(net2793),
    .A1(net330),
    .S(net2846),
    .X(_00056_));
 sg13g2_nand2_1 _19844_ (.Y(_00298_),
    .A(net2838),
    .B(net282));
 sg13g2_o21ai_1 _19845_ (.B1(_00298_),
    .Y(_00057_),
    .A1(_05913_),
    .A2(net2838));
 sg13g2_mux2_1 _19846_ (.A0(net2787),
    .A1(net293),
    .S(net2818),
    .X(_00058_));
 sg13g2_nand2_1 _19847_ (.Y(_00299_),
    .A(net2773),
    .B(net2871));
 sg13g2_o21ai_1 _19848_ (.B1(_00299_),
    .Y(_00059_),
    .A1(_05869_),
    .A2(net2871));
 sg13g2_mux2_1 _19849_ (.A0(net2782),
    .A1(net2772),
    .S(net2871),
    .X(_00060_));
 sg13g2_nor2_1 _19850_ (.A(net2778),
    .B(net2826),
    .Y(_00300_));
 sg13g2_a21oi_1 _19851_ (.A1(_05627_),
    .A2(net2827),
    .Y(_00061_),
    .B1(_00300_));
 sg13g2_mux2_1 _19852_ (.A0(net2776),
    .A1(net2766),
    .S(net2823),
    .X(_00062_));
 sg13g2_nor2_1 _19853_ (.A(net2774),
    .B(net2883),
    .Y(_00302_));
 sg13g2_a21oi_1 _19854_ (.A1(_05143_),
    .A2(net2883),
    .Y(_00063_),
    .B1(_00302_));
 sg13g2_mux2_1 _19855_ (.A0(net330),
    .A1(net2762),
    .S(net2841),
    .X(_00064_));
 sg13g2_nor2_1 _19856_ (.A(net2838),
    .B(net282),
    .Y(_00303_));
 sg13g2_a21oi_1 _19857_ (.A1(_06023_),
    .A2(net2838),
    .Y(_00065_),
    .B1(_00303_));
 sg13g2_mux2_1 _19858_ (.A0(net293),
    .A1(net2757),
    .S(net2818),
    .X(_00066_));
 sg13g2_nor2_1 _19859_ (.A(net2773),
    .B(net2858),
    .Y(_00304_));
 sg13g2_a21oi_1 _19860_ (.A1(_05495_),
    .A2(net2859),
    .Y(_00067_),
    .B1(_00304_));
 sg13g2_mux2_1 _19861_ (.A0(net2772),
    .A1(net2753),
    .S(net2855),
    .X(_00068_));
 sg13g2_nand2_1 _19862_ (.Y(_00306_),
    .A(net2750),
    .B(net2828));
 sg13g2_o21ai_1 _19863_ (.B1(_00306_),
    .Y(_00069_),
    .A1(_05627_),
    .A2(net2828));
 sg13g2_mux2_1 _19864_ (.A0(net2766),
    .A1(net2748),
    .S(net2838),
    .X(_00070_));
 sg13g2_nor2_1 _19865_ (.A(net2764),
    .B(net2840),
    .Y(_00307_));
 sg13g2_a21oi_1 _19866_ (.A1(_05891_),
    .A2(net2840),
    .Y(_00071_),
    .B1(_00307_));
 sg13g2_mux2_1 _19867_ (.A0(net2763),
    .A1(net302),
    .S(net2852),
    .X(_00072_));
 sg13g2_nand2_1 _19868_ (.Y(_00308_),
    .A(net2838),
    .B(net275));
 sg13g2_o21ai_1 _19869_ (.B1(_00308_),
    .Y(_00073_),
    .A1(_06023_),
    .A2(net2838));
 sg13g2_mux2_1 _19870_ (.A0(net2757),
    .A1(\net.in[49] ),
    .S(net2824),
    .X(_00074_));
 sg13g2_nor2_1 _19871_ (.A(net2755),
    .B(net2874),
    .Y(_00309_));
 sg13g2_a21oi_1 _19872_ (.A1(_06001_),
    .A2(net2874),
    .Y(_00075_),
    .B1(_00309_));
 sg13g2_mux2_1 _19873_ (.A0(net2753),
    .A1(net2742),
    .S(net2823),
    .X(_00076_));
 sg13g2_nor2_1 _19874_ (.A(net2750),
    .B(net2839),
    .Y(_00311_));
 sg13g2_a21oi_1 _19875_ (.A1(_05946_),
    .A2(net2839),
    .Y(_00077_),
    .B1(_00311_));
 sg13g2_mux2_1 _19876_ (.A0(net2748),
    .A1(net2734),
    .S(net2846),
    .X(_00078_));
 sg13g2_nand2_1 _19877_ (.Y(_00312_),
    .A(net2731),
    .B(net2840));
 sg13g2_o21ai_1 _19878_ (.B1(_00312_),
    .Y(_00079_),
    .A1(_05891_),
    .A2(net2840));
 sg13g2_nor2_1 _19879_ (.A(net2745),
    .B(net2857),
    .Y(_00313_));
 sg13g2_a21oi_1 _19880_ (.A1(_05451_),
    .A2(net2857),
    .Y(_00080_),
    .B1(_00313_));
 sg13g2_mux2_1 _19881_ (.A0(net275),
    .A1(net2726),
    .S(net2838),
    .X(_00081_));
 sg13g2_mux2_1 _19882_ (.A0(\net.in[49] ),
    .A1(net2722),
    .S(net2824),
    .X(_00082_));
 sg13g2_nand2_1 _19883_ (.Y(_00315_),
    .A(net2718),
    .B(net2873));
 sg13g2_o21ai_1 _19884_ (.B1(_00315_),
    .Y(_00083_),
    .A1(_06001_),
    .A2(net2873));
 sg13g2_nor2_1 _19885_ (.A(net2741),
    .B(net2854),
    .Y(_00316_));
 sg13g2_a21oi_1 _19886_ (.A1(_05957_),
    .A2(net2856),
    .Y(_00084_),
    .B1(_00316_));
 sg13g2_nand2_1 _19887_ (.Y(_00317_),
    .A(net2711),
    .B(net2840));
 sg13g2_o21ai_1 _19888_ (.B1(_00317_),
    .Y(_00085_),
    .A1(_05946_),
    .A2(net2839));
 sg13g2_nor2_1 _19889_ (.A(net2736),
    .B(net2877),
    .Y(_00318_));
 sg13g2_a21oi_1 _19890_ (.A1(_05561_),
    .A2(net2877),
    .Y(_00086_),
    .B1(_00318_));
 sg13g2_nor2_1 _19891_ (.A(net2731),
    .B(net2839),
    .Y(_00319_));
 sg13g2_a21oi_1 _19892_ (.A1(_05748_),
    .A2(net2839),
    .Y(_00087_),
    .B1(_00319_));
 sg13g2_nand2_1 _19893_ (.Y(_00321_),
    .A(net2705),
    .B(net2858));
 sg13g2_o21ai_1 _19894_ (.B1(_00321_),
    .Y(_00088_),
    .A1(_05451_),
    .A2(net2858));
 sg13g2_mux2_1 _19895_ (.A0(net2725),
    .A1(net291),
    .S(net2818),
    .X(_00089_));
 sg13g2_mux2_1 _19896_ (.A0(net2723),
    .A1(net2704),
    .S(net2870),
    .X(_00090_));
 sg13g2_mux2_1 _19897_ (.A0(net2717),
    .A1(net2702),
    .S(net2834),
    .X(_00091_));
 sg13g2_nand2_1 _19898_ (.Y(_00322_),
    .A(net2701),
    .B(net2831));
 sg13g2_o21ai_1 _19899_ (.B1(_00322_),
    .Y(_00092_),
    .A1(_05957_),
    .A2(net2831));
 sg13g2_nor2_1 _19900_ (.A(net2711),
    .B(net2843),
    .Y(_00323_));
 sg13g2_a21oi_1 _19901_ (.A1(_05011_),
    .A2(net2843),
    .Y(_00093_),
    .B1(_00323_));
 sg13g2_nand2_1 _19902_ (.Y(_00325_),
    .A(net2697),
    .B(net2878));
 sg13g2_o21ai_1 _19903_ (.B1(_00325_),
    .Y(_00094_),
    .A1(_05561_),
    .A2(net2878));
 sg13g2_nand2_1 _19904_ (.Y(_00326_),
    .A(net2690),
    .B(net2839));
 sg13g2_o21ai_1 _19905_ (.B1(_00326_),
    .Y(_00095_),
    .A1(_05748_),
    .A2(net2839));
 sg13g2_mux2_1 _19906_ (.A0(net2705),
    .A1(net2688),
    .S(net2872),
    .X(_00096_));
 sg13g2_nor2_1 _19907_ (.A(net2818),
    .B(net291),
    .Y(_00327_));
 sg13g2_a21oi_1 _19908_ (.A1(net2177),
    .A2(net2819),
    .Y(_00097_),
    .B1(_00327_));
 sg13g2_mux2_1 _19909_ (.A0(net2704),
    .A1(net2679),
    .S(net2870),
    .X(_00098_));
 sg13g2_nor2_1 _19910_ (.A(net2702),
    .B(net2842),
    .Y(_00328_));
 sg13g2_a21oi_1 _19911_ (.A1(_05715_),
    .A2(net2842),
    .Y(_00099_),
    .B1(_00328_));
 sg13g2_mux2_1 _19912_ (.A0(net2700),
    .A1(net2673),
    .S(net2835),
    .X(_00100_));
 sg13g2_nand2_1 _19913_ (.Y(_00330_),
    .A(net2668),
    .B(net2840));
 sg13g2_o21ai_1 _19914_ (.B1(_00330_),
    .Y(_00101_),
    .A1(_05011_),
    .A2(net2840));
 sg13g2_mux2_1 _19915_ (.A0(net2697),
    .A1(net2667),
    .S(net2871),
    .X(_00102_));
 sg13g2_mux2_1 _19916_ (.A0(net2692),
    .A1(net2663),
    .S(net2887),
    .X(_00103_));
 sg13g2_nor2_1 _19917_ (.A(net2687),
    .B(net2876),
    .Y(_00331_));
 sg13g2_a21oi_1 _19918_ (.A1(_05836_),
    .A2(net2876),
    .Y(_00104_),
    .B1(_00331_));
 sg13g2_nand2_1 _19919_ (.Y(_00332_),
    .A(\net.in[80] ),
    .B(net2855));
 sg13g2_o21ai_1 _19920_ (.B1(_00332_),
    .Y(_00105_),
    .A1(net2177),
    .A2(net2855));
 sg13g2_mux2_1 _19921_ (.A0(net2678),
    .A1(net304),
    .S(net2882),
    .X(_00106_));
 sg13g2_nand2_1 _19922_ (.Y(_00334_),
    .A(net2656),
    .B(net2842));
 sg13g2_o21ai_1 _19923_ (.B1(_00334_),
    .Y(_00107_),
    .A1(_05715_),
    .A2(net2842));
 sg13g2_nor2_1 _19924_ (.A(net2672),
    .B(net2859),
    .Y(_00335_));
 sg13g2_a21oi_1 _19925_ (.A1(_05572_),
    .A2(net2859),
    .Y(_00108_),
    .B1(_00335_));
 sg13g2_mux2_1 _19926_ (.A0(net2670),
    .A1(net2650),
    .S(net2871),
    .X(_00109_));
 sg13g2_nor2_1 _19927_ (.A(net2667),
    .B(net2852),
    .Y(_00336_));
 sg13g2_a21oi_1 _19928_ (.A1(_05880_),
    .A2(net2851),
    .Y(_00110_),
    .B1(_00336_));
 sg13g2_mux2_1 _19929_ (.A0(net2662),
    .A1(net2642),
    .S(net2822),
    .X(_00111_));
 sg13g2_nand2_1 _19930_ (.Y(_00337_),
    .A(net2640),
    .B(net2879));
 sg13g2_o21ai_1 _19931_ (.B1(_00337_),
    .Y(_00112_),
    .A1(_05836_),
    .A2(net2879));
 sg13g2_nor2_1 _19932_ (.A(\net.in[80] ),
    .B(net2861),
    .Y(_00339_));
 sg13g2_a21oi_1 _19933_ (.A1(_05726_),
    .A2(net2861),
    .Y(_00113_),
    .B1(_00339_));
 sg13g2_nor2_1 _19934_ (.A(net304),
    .B(net2881),
    .Y(_00340_));
 sg13g2_a21oi_1 _19935_ (.A1(_05594_),
    .A2(net2881),
    .Y(_00114_),
    .B1(_00340_));
 sg13g2_mux2_1 _19936_ (.A0(net2657),
    .A1(net2628),
    .S(net2857),
    .X(_00115_));
 sg13g2_nand2_1 _19937_ (.Y(_00341_),
    .A(net2621),
    .B(net2859));
 sg13g2_o21ai_1 _19938_ (.B1(_00341_),
    .Y(_00116_),
    .A1(_05572_),
    .A2(net2859));
 sg13g2_nor2_1 _19939_ (.A(net2651),
    .B(net2887),
    .Y(_00342_));
 sg13g2_a21oi_1 _19940_ (.A1(_05770_),
    .A2(net2887),
    .Y(_00117_),
    .B1(_00342_));
 sg13g2_nor2_1 _19941_ (.A(net2647),
    .B(net2848),
    .Y(_00343_));
 sg13g2_a21oi_1 _19942_ (.A1(_05231_),
    .A2(net2848),
    .Y(_00118_),
    .B1(_00343_));
 sg13g2_mux2_1 _19943_ (.A0(net2644),
    .A1(net2608),
    .S(net2858),
    .X(_00119_));
 sg13g2_mux2_1 _19944_ (.A0(net2640),
    .A1(net2604),
    .S(net2870),
    .X(_00120_));
 sg13g2_nand2_1 _19945_ (.Y(_00345_),
    .A(net321),
    .B(net2859));
 sg13g2_o21ai_1 _19946_ (.B1(_00345_),
    .Y(_00121_),
    .A1(_05726_),
    .A2(net2859));
 sg13g2_nand2_1 _19947_ (.Y(_00346_),
    .A(net2603),
    .B(net2883));
 sg13g2_o21ai_1 _19948_ (.B1(_00346_),
    .Y(_00122_),
    .A1(_05594_),
    .A2(net2883));
 sg13g2_mux2_1 _19949_ (.A0(net2627),
    .A1(net2601),
    .S(net2873),
    .X(_00123_));
 sg13g2_mux2_1 _19950_ (.A0(net2618),
    .A1(net2596),
    .S(net2820),
    .X(_00124_));
 sg13g2_nor2_1 _19951_ (.A(net2615),
    .B(net2834),
    .Y(_00347_));
 sg13g2_a21oi_1 _19952_ (.A1(_05858_),
    .A2(net2834),
    .Y(_00125_),
    .B1(_00347_));
 sg13g2_nor2_1 _19953_ (.A(net2612),
    .B(net2866),
    .Y(_00349_));
 sg13g2_a21oi_1 _19954_ (.A1(_05682_),
    .A2(net2866),
    .Y(_00126_),
    .B1(_00349_));
 sg13g2_nor2_1 _19955_ (.A(net2607),
    .B(net2875),
    .Y(_00350_));
 sg13g2_a21oi_1 _19956_ (.A1(_05693_),
    .A2(net2875),
    .Y(_00127_),
    .B1(_00350_));
 sg13g2_mux2_1 _19957_ (.A0(net2604),
    .A1(net2577),
    .S(net2871),
    .X(_00128_));
 sg13g2_mux2_1 _19958_ (.A0(net321),
    .A1(net2573),
    .S(net2865),
    .X(_00129_));
 sg13g2_nor2_1 _19959_ (.A(net2603),
    .B(net2853),
    .Y(_00351_));
 sg13g2_a21oi_1 _19960_ (.A1(net2178),
    .A2(net2853),
    .Y(_00130_),
    .B1(_00351_));
 sg13g2_nor2_1 _19961_ (.A(net320),
    .B(net2867),
    .Y(_00352_));
 sg13g2_a21oi_1 _19962_ (.A1(_05814_),
    .A2(net2866),
    .Y(_00131_),
    .B1(_00352_));
 sg13g2_nor2_1 _19963_ (.A(net2599),
    .B(net2885),
    .Y(_00354_));
 sg13g2_a21oi_2 _19964_ (.B1(_00354_),
    .Y(_00132_),
    .A2(net2885),
    .A1(_05220_));
 sg13g2_nor2_1 _19965_ (.A(net2595),
    .B(net2857),
    .Y(_00355_));
 sg13g2_a21oi_1 _19966_ (.A1(_05330_),
    .A2(net2857),
    .Y(_00133_),
    .B1(_00355_));
 sg13g2_nor2_1 _19967_ (.A(net2590),
    .B(net2870),
    .Y(_00356_));
 sg13g2_a21oi_1 _19968_ (.A1(_05176_),
    .A2(net2870),
    .Y(_00134_),
    .B1(_00356_));
 sg13g2_nand2_1 _19969_ (.Y(_00357_),
    .A(net2552),
    .B(net2826));
 sg13g2_o21ai_1 _19970_ (.B1(_00357_),
    .Y(_00135_),
    .A1(_05693_),
    .A2(net2826));
 sg13g2_mux2_1 _19971_ (.A0(net2577),
    .A1(net2551),
    .S(net2870),
    .X(_00136_));
 sg13g2_nor2_1 _19972_ (.A(net2572),
    .B(net2848),
    .Y(_00359_));
 sg13g2_a21oi_1 _19973_ (.A1(_05825_),
    .A2(net2848),
    .Y(_00137_),
    .B1(_00359_));
 sg13g2_nand2_1 _19974_ (.Y(_00360_),
    .A(net2548),
    .B(net2830));
 sg13g2_o21ai_1 _19975_ (.B1(_00360_),
    .Y(_00138_),
    .A1(_05385_),
    .A2(net2830));
 sg13g2_nand2_1 _19976_ (.Y(_00361_),
    .A(net2546),
    .B(net2866));
 sg13g2_o21ai_1 _19977_ (.B1(_00361_),
    .Y(_00139_),
    .A1(_05814_),
    .A2(net2866));
 sg13g2_nand2_1 _19978_ (.Y(_00362_),
    .A(net2542),
    .B(net2884));
 sg13g2_o21ai_1 _19979_ (.B1(_00362_),
    .Y(_00140_),
    .A1(_05220_),
    .A2(net2884));
 sg13g2_nand2_1 _19980_ (.Y(_00363_),
    .A(net2538),
    .B(net2860));
 sg13g2_o21ai_1 _19981_ (.B1(_00363_),
    .Y(_00141_),
    .A1(_05330_),
    .A2(net2860));
 sg13g2_nand2_1 _19982_ (.Y(_00365_),
    .A(net2532),
    .B(net2871));
 sg13g2_o21ai_1 _19983_ (.B1(_00365_),
    .Y(_00142_),
    .A1(_05176_),
    .A2(net2870));
 sg13g2_nor2_1 _19984_ (.A(net2552),
    .B(net2881),
    .Y(_00366_));
 sg13g2_a21oi_1 _19985_ (.A1(_05242_),
    .A2(net2881),
    .Y(_00143_),
    .B1(_00366_));
 sg13g2_nor2_1 _19986_ (.A(net2550),
    .B(net2883),
    .Y(_00367_));
 sg13g2_a21oi_1 _19987_ (.A1(net2183),
    .A2(net2883),
    .Y(_00144_),
    .B1(_00367_));
 sg13g2_nor2_1 _19988_ (.A(net381),
    .B(net2882),
    .Y(_00368_));
 sg13g2_a21oi_1 _19989_ (.A1(net2181),
    .A2(net2882),
    .Y(_00145_),
    .B1(_00368_));
 sg13g2_mux2_1 _19990_ (.A0(net2548),
    .A1(net2513),
    .S(net2825),
    .X(_00146_));
 sg13g2_mux2_1 _19991_ (.A0(net2547),
    .A1(net2509),
    .S(net2822),
    .X(_00147_));
 sg13g2_nor2_1 _19992_ (.A(net2539),
    .B(net2827),
    .Y(_00370_));
 sg13g2_a21oi_1 _19993_ (.A1(_05165_),
    .A2(net2826),
    .Y(_00148_),
    .B1(_00370_));
 sg13g2_mux2_1 _19994_ (.A0(net2534),
    .A1(net2502),
    .S(net2820),
    .X(_00149_));
 sg13g2_mux2_1 _19995_ (.A0(net2531),
    .A1(net2500),
    .S(net2873),
    .X(_00150_));
 sg13g2_nor2_1 _19996_ (.A(net2527),
    .B(net2854),
    .Y(_00371_));
 sg13g2_a21oi_1 _19997_ (.A1(_05088_),
    .A2(net2854),
    .Y(_00151_),
    .B1(_00371_));
 sg13g2_nand2_1 _19998_ (.Y(_00372_),
    .A(net2497),
    .B(net2867));
 sg13g2_o21ai_1 _19999_ (.B1(_00372_),
    .Y(_00152_),
    .A1(net2183),
    .A2(net2883));
 sg13g2_nand2_1 _20000_ (.Y(_00373_),
    .A(net2887),
    .B(net277));
 sg13g2_o21ai_1 _20001_ (.B1(_00373_),
    .Y(_00153_),
    .A1(net2181),
    .A2(net2887));
 sg13g2_mux2_1 _20002_ (.A0(net2513),
    .A1(net2496),
    .S(net2825),
    .X(_00154_));
 sg13g2_mux2_1 _20003_ (.A0(net2509),
    .A1(net2492),
    .S(net2821),
    .X(_00155_));
 sg13g2_nor2_1 _20004_ (.A(net2505),
    .B(net2842),
    .Y(_00375_));
 sg13g2_a21oi_1 _20005_ (.A1(_05671_),
    .A2(net2842),
    .Y(_00156_),
    .B1(_00375_));
 sg13g2_mux2_1 _20006_ (.A0(net2502),
    .A1(net2484),
    .S(net2818),
    .X(_00157_));
 sg13g2_nor2_1 _20007_ (.A(net2501),
    .B(net2855),
    .Y(_00376_));
 sg13g2_a21oi_1 _20008_ (.A1(_05000_),
    .A2(net2855),
    .Y(_00158_),
    .B1(_00376_));
 sg13g2_nand2_1 _20009_ (.Y(_00377_),
    .A(net2480),
    .B(net2854));
 sg13g2_o21ai_1 _20010_ (.B1(_00377_),
    .Y(_00159_),
    .A1(_05088_),
    .A2(net2854));
 sg13g2_mux2_1 _20011_ (.A0(net2497),
    .A1(net2475),
    .S(net2876),
    .X(_00160_));
 sg13g2_nor2_1 _20012_ (.A(net2887),
    .B(net277),
    .Y(_00379_));
 sg13g2_a21oi_1 _20013_ (.A1(_05044_),
    .A2(net2888),
    .Y(_00161_),
    .B1(_00379_));
 sg13g2_nor2_1 _20014_ (.A(\net.in[129] ),
    .B(net2867),
    .Y(_00380_));
 sg13g2_a21oi_2 _20015_ (.B1(_00380_),
    .Y(_00162_),
    .A2(net2867),
    .A1(_05187_));
 sg13g2_nor2_1 _20016_ (.A(net2493),
    .B(net2848),
    .Y(_00381_));
 sg13g2_a21oi_1 _20017_ (.A1(net2179),
    .A2(net2848),
    .Y(_00163_),
    .B1(_00381_));
 sg13g2_nor2_1 _20018_ (.A(net2490),
    .B(net2852),
    .Y(_00382_));
 sg13g2_a21oi_1 _20019_ (.A1(_05440_),
    .A2(net2852),
    .Y(_00164_),
    .B1(_00382_));
 sg13g2_mux2_1 _20020_ (.A0(net2484),
    .A1(net2457),
    .S(net2825),
    .X(_00165_));
 sg13g2_nand2_1 _20021_ (.Y(_00383_),
    .A(net2455),
    .B(net2852));
 sg13g2_o21ai_1 _20022_ (.B1(_00383_),
    .Y(_00166_),
    .A1(_05000_),
    .A2(net2852));
 sg13g2_nor2_1 _20023_ (.A(net2478),
    .B(net2867),
    .Y(_00385_));
 sg13g2_a21oi_1 _20024_ (.A1(_05099_),
    .A2(net2866),
    .Y(_00167_),
    .B1(_00385_));
 sg13g2_mux2_1 _20025_ (.A0(net2473),
    .A1(net2448),
    .S(net2824),
    .X(_00168_));
 sg13g2_nand2_1 _20026_ (.Y(_00386_),
    .A(net284),
    .B(net2876));
 sg13g2_o21ai_1 _20027_ (.B1(_00386_),
    .Y(_00169_),
    .A1(_05044_),
    .A2(net2876));
 sg13g2_nand2_1 _20028_ (.Y(_00387_),
    .A(net331),
    .B(net2831));
 sg13g2_o21ai_1 _20029_ (.B1(_00387_),
    .Y(_00170_),
    .A1(_05187_),
    .A2(net2831));
 sg13g2_nor2_1 _20030_ (.A(net2463),
    .B(net2842),
    .Y(_00388_));
 sg13g2_a21oi_1 _20031_ (.A1(_05407_),
    .A2(net2842),
    .Y(_00171_),
    .B1(_00388_));
 sg13g2_nor2_1 _20032_ (.A(\net.in[139] ),
    .B(net2857),
    .Y(_00390_));
 sg13g2_a21oi_1 _20033_ (.A1(_05297_),
    .A2(net2858),
    .Y(_00172_),
    .B1(_00390_));
 sg13g2_nor2_1 _20034_ (.A(net2459),
    .B(net2874),
    .Y(_00391_));
 sg13g2_a21oi_1 _20035_ (.A1(_05418_),
    .A2(net2874),
    .Y(_00173_),
    .B1(_00391_));
 sg13g2_nor2_1 _20036_ (.A(net2455),
    .B(net2862),
    .Y(_00392_));
 sg13g2_a21oi_1 _20037_ (.A1(_05286_),
    .A2(net2862),
    .Y(_00174_),
    .B1(_00392_));
 sg13g2_nor2_1 _20038_ (.A(net2452),
    .B(net2833),
    .Y(_00393_));
 sg13g2_a21oi_1 _20039_ (.A1(_05022_),
    .A2(net2833),
    .Y(_00175_),
    .B1(_00393_));
 sg13g2_mux2_1 _20040_ (.A0(net2449),
    .A1(net2426),
    .S(net2824),
    .X(_00176_));
 sg13g2_nor2_1 _20041_ (.A(net284),
    .B(net2876),
    .Y(_00394_));
 sg13g2_a21oi_1 _20042_ (.A1(_05264_),
    .A2(net2875),
    .Y(_00177_),
    .B1(_00394_));
 sg13g2_mux2_1 _20043_ (.A0(\net.in[145] ),
    .A1(net2418),
    .S(net2836),
    .X(_00178_));
 sg13g2_nand2_1 _20044_ (.Y(_00396_),
    .A(net2415),
    .B(net2848));
 sg13g2_o21ai_1 _20045_ (.B1(_00396_),
    .Y(_00179_),
    .A1(_05407_),
    .A2(net2848));
 sg13g2_nor2_1 _20046_ (.A(net2443),
    .B(net2860),
    .Y(_00397_));
 sg13g2_a21oi_1 _20047_ (.A1(_05352_),
    .A2(net2860),
    .Y(_00180_),
    .B1(_00397_));
 sg13g2_nor2_1 _20048_ (.A(net2437),
    .B(net2820),
    .Y(_00398_));
 sg13g2_a21oi_1 _20049_ (.A1(_05968_),
    .A2(net2820),
    .Y(_00181_),
    .B1(_00398_));
 sg13g2_nand2_1 _20050_ (.Y(_00399_),
    .A(net2408),
    .B(net2862));
 sg13g2_o21ai_1 _20051_ (.B1(_00399_),
    .Y(_00182_),
    .A1(_05286_),
    .A2(net2862));
 sg13g2_nand2_1 _20052_ (.Y(_00401_),
    .A(net2405),
    .B(net2829));
 sg13g2_o21ai_1 _20053_ (.B1(_00401_),
    .Y(_00183_),
    .A1(_05022_),
    .A2(net2829));
 sg13g2_mux2_1 _20054_ (.A0(net2428),
    .A1(net2404),
    .S(net2864),
    .X(_00184_));
 sg13g2_nand2_1 _20055_ (.Y(_00402_),
    .A(net2863),
    .B(net278));
 sg13g2_o21ai_1 _20056_ (.B1(_00402_),
    .Y(_00185_),
    .A1(_05264_),
    .A2(net2863));
 sg13g2_mux2_1 _20057_ (.A0(net2419),
    .A1(\net.in[161] ),
    .S(net2887),
    .X(_00186_));
 sg13g2_mux2_1 _20058_ (.A0(net2417),
    .A1(net2401),
    .S(net2851),
    .X(_00187_));
 sg13g2_nand2_1 _20059_ (.Y(_00403_),
    .A(net2400),
    .B(net2857));
 sg13g2_o21ai_1 _20060_ (.B1(_00403_),
    .Y(_00188_),
    .A1(_05352_),
    .A2(net2857));
 sg13g2_nand2_1 _20061_ (.Y(_00404_),
    .A(net2393),
    .B(net2820));
 sg13g2_o21ai_1 _20062_ (.B1(_00404_),
    .Y(_00189_),
    .A1(_05968_),
    .A2(net2820));
 sg13g2_nor2_1 _20063_ (.A(net2408),
    .B(net2865),
    .Y(_00406_));
 sg13g2_a21oi_2 _20064_ (.B1(_00406_),
    .Y(_00190_),
    .A2(net2865),
    .A1(_05308_));
 sg13g2_nor2_1 _20065_ (.A(net2406),
    .B(net2863),
    .Y(_00407_));
 sg13g2_a21oi_1 _20066_ (.A1(_05539_),
    .A2(net2863),
    .Y(_00191_),
    .B1(_00407_));
 sg13g2_nor2_1 _20067_ (.A(net2404),
    .B(net2865),
    .Y(_00408_));
 sg13g2_a21oi_1 _20068_ (.A1(_05363_),
    .A2(net2866),
    .Y(_00192_),
    .B1(_00408_));
 sg13g2_nor2_1 _20069_ (.A(net2874),
    .B(net278),
    .Y(_00409_));
 sg13g2_a21oi_1 _20070_ (.A1(_05462_),
    .A2(net2875),
    .Y(_00193_),
    .B1(_00409_));
 sg13g2_nor2_1 _20071_ (.A(\net.in[161] ),
    .B(net2884),
    .Y(_00410_));
 sg13g2_a21oi_1 _20072_ (.A1(_05638_),
    .A2(net2883),
    .Y(_00194_),
    .B1(_00410_));
 sg13g2_mux2_1 _20073_ (.A0(net2403),
    .A1(net2371),
    .S(net2825),
    .X(_00195_));
 sg13g2_nor2_1 _20074_ (.A(net2400),
    .B(net2885),
    .Y(_00412_));
 sg13g2_a21oi_1 _20075_ (.A1(_05781_),
    .A2(net2885),
    .Y(_00196_),
    .B1(_00412_));
 sg13g2_mux2_1 _20076_ (.A0(net2393),
    .A1(net2364),
    .S(net2822),
    .X(_00197_));
 sg13g2_nand2_1 _20077_ (.Y(_00413_),
    .A(net2362),
    .B(net2826));
 sg13g2_o21ai_1 _20078_ (.B1(_00413_),
    .Y(_00198_),
    .A1(net2180),
    .A2(net2826));
 sg13g2_nand2_1 _20079_ (.Y(_00414_),
    .A(net2361),
    .B(net2863));
 sg13g2_o21ai_1 _20080_ (.B1(_00414_),
    .Y(_00199_),
    .A1(_05539_),
    .A2(net2863));
 sg13g2_nand2_1 _20081_ (.Y(_00415_),
    .A(\net.in[175] ),
    .B(net2855));
 sg13g2_o21ai_1 _20082_ (.B1(_00415_),
    .Y(_00200_),
    .A1(_05363_),
    .A2(net2855));
 sg13g2_nand2_1 _20083_ (.Y(_00417_),
    .A(net313),
    .B(net2875));
 sg13g2_o21ai_1 _20084_ (.B1(_00417_),
    .Y(_00201_),
    .A1(_05462_),
    .A2(net2875));
 sg13g2_nand2_1 _20085_ (.Y(_00418_),
    .A(net2360),
    .B(net2884));
 sg13g2_o21ai_1 _20086_ (.B1(_00418_),
    .Y(_00202_),
    .A1(_05638_),
    .A2(net2884));
 sg13g2_mux2_1 _20087_ (.A0(net2374),
    .A1(net2358),
    .S(net2853),
    .X(_00203_));
 sg13g2_nor2_1 _20088_ (.A(net2369),
    .B(net2876),
    .Y(_00419_));
 sg13g2_a21oi_1 _20089_ (.A1(_05473_),
    .A2(net2875),
    .Y(_00204_),
    .B1(_00419_));
 sg13g2_mux2_1 _20090_ (.A0(net2364),
    .A1(net2349),
    .S(net2822),
    .X(_00205_));
 sg13g2_nor2_1 _20091_ (.A(net2363),
    .B(net2861),
    .Y(_00420_));
 sg13g2_a21oi_1 _20092_ (.A1(_05121_),
    .A2(net2859),
    .Y(_00206_),
    .B1(_00420_));
 sg13g2_mux2_1 _20093_ (.A0(net2361),
    .A1(net2342),
    .S(net2851),
    .X(_00207_));
 sg13g2_nor2_1 _20094_ (.A(\net.in[175] ),
    .B(net2854),
    .Y(_00422_));
 sg13g2_a21oi_1 _20095_ (.A1(_05209_),
    .A2(net2854),
    .Y(_00208_),
    .B1(_00422_));
 sg13g2_mux2_1 _20096_ (.A0(net313),
    .A1(net2333),
    .S(net2877),
    .X(_00209_));
 sg13g2_nor2_1 _20097_ (.A(net2359),
    .B(net2828),
    .Y(_00423_));
 sg13g2_a21oi_1 _20098_ (.A1(_05803_),
    .A2(net2828),
    .Y(_00210_),
    .B1(_00423_));
 sg13g2_mux2_1 _20099_ (.A0(net2358),
    .A1(net2326),
    .S(net2873),
    .X(_00211_));
 sg13g2_nor2_1 _20100_ (.A(net2354),
    .B(net2832),
    .Y(_00424_));
 sg13g2_a21oi_1 _20101_ (.A1(_05275_),
    .A2(net2832),
    .Y(_00212_),
    .B1(_00424_));
 sg13g2_mux2_1 _20102_ (.A0(net2349),
    .A1(net2320),
    .S(net2825),
    .X(_00213_));
 sg13g2_nand2_1 _20103_ (.Y(_00426_),
    .A(net305),
    .B(net2867));
 sg13g2_o21ai_1 _20104_ (.B1(_00426_),
    .Y(_00214_),
    .A1(_05121_),
    .A2(net2867));
 sg13g2_mux2_1 _20105_ (.A0(net2342),
    .A1(net2316),
    .S(net2851),
    .X(_00215_));
 sg13g2_nand2_1 _20106_ (.Y(_00427_),
    .A(\net.in[191] ),
    .B(net2862));
 sg13g2_o21ai_1 _20107_ (.B1(_00427_),
    .Y(_00216_),
    .A1(_05209_),
    .A2(net2862));
 sg13g2_mux2_1 _20108_ (.A0(net2333),
    .A1(net329),
    .S(net2877),
    .X(_00217_));
 sg13g2_nand2_1 _20109_ (.Y(_00428_),
    .A(net2315),
    .B(net2829));
 sg13g2_o21ai_1 _20110_ (.B1(_00428_),
    .Y(_00218_),
    .A1(_05803_),
    .A2(net2829));
 sg13g2_nor2_1 _20111_ (.A(net2325),
    .B(net2836),
    .Y(_00429_));
 sg13g2_a21oi_1 _20112_ (.A1(_05319_),
    .A2(net2836),
    .Y(_00219_),
    .B1(_00429_));
 sg13g2_nand2_1 _20113_ (.Y(_00431_),
    .A(net2310),
    .B(net2833));
 sg13g2_o21ai_1 _20114_ (.B1(_00431_),
    .Y(_00220_),
    .A1(_05275_),
    .A2(net2833));
 sg13g2_nor2_1 _20115_ (.A(net2320),
    .B(net2833),
    .Y(_00432_));
 sg13g2_a21oi_1 _20116_ (.A1(_05066_),
    .A2(net2833),
    .Y(_00221_),
    .B1(_00432_));
 sg13g2_mux2_1 _20117_ (.A0(net2319),
    .A1(net2299),
    .S(net2818),
    .X(_00222_));
 sg13g2_nor2_1 _20118_ (.A(net2316),
    .B(net2832),
    .Y(_00433_));
 sg13g2_a21oi_1 _20119_ (.A1(_05077_),
    .A2(net2832),
    .Y(_00223_),
    .B1(_00433_));
 sg13g2_nor2_1 _20120_ (.A(\net.in[191] ),
    .B(net2855),
    .Y(_00434_));
 sg13g2_a21oi_1 _20121_ (.A1(_05484_),
    .A2(net2862),
    .Y(_00224_),
    .B1(_00434_));
 sg13g2_mux2_1 _20122_ (.A0(\net.in[192] ),
    .A1(net309),
    .S(net2877),
    .X(_00225_));
 sg13g2_mux2_1 _20123_ (.A0(net2315),
    .A1(net306),
    .S(net2872),
    .X(_00226_));
 sg13g2_nand2_1 _20124_ (.Y(_00436_),
    .A(net2286),
    .B(net2868));
 sg13g2_o21ai_1 _20125_ (.B1(_00436_),
    .Y(_00227_),
    .A1(_05319_),
    .A2(net2868));
 sg13g2_mux2_1 _20126_ (.A0(net2309),
    .A1(net2282),
    .S(net2819),
    .X(_00228_));
 sg13g2_nor2_1 _20127_ (.A(net2307),
    .B(net2860),
    .Y(_00437_));
 sg13g2_a21oi_1 _20128_ (.A1(_06056_),
    .A2(net2860),
    .Y(_00229_),
    .B1(_00437_));
 sg13g2_mux2_1 _20129_ (.A0(net2299),
    .A1(net2279),
    .S(net2819),
    .X(_00230_));
 sg13g2_nand2_1 _20130_ (.Y(_00438_),
    .A(net2277),
    .B(net2830));
 sg13g2_o21ai_1 _20131_ (.B1(_00438_),
    .Y(_00231_),
    .A1(_05077_),
    .A2(net2830));
 sg13g2_nand2_1 _20132_ (.Y(_00440_),
    .A(net2276),
    .B(net2865));
 sg13g2_o21ai_1 _20133_ (.B1(_00440_),
    .Y(_00232_),
    .A1(_05484_),
    .A2(net2865));
 sg13g2_mux2_1 _20134_ (.A0(net2290),
    .A1(net324),
    .S(net2833),
    .X(_00233_));
 sg13g2_mux2_1 _20135_ (.A0(net2287),
    .A1(\net.in[209] ),
    .S(net2834),
    .X(_00234_));
 sg13g2_nor2_1 _20136_ (.A(net2285),
    .B(net2827),
    .Y(_00441_));
 sg13g2_a21oi_2 _20137_ (.B1(_00441_),
    .Y(_00235_),
    .A2(net2834),
    .A1(_05935_));
 sg13g2_mux2_1 _20138_ (.A0(net2282),
    .A1(net2269),
    .S(net2821),
    .X(_00236_));
 sg13g2_nor2_1 _20139_ (.A(net2281),
    .B(net2881),
    .Y(_00442_));
 sg13g2_a21oi_1 _20140_ (.A1(_05528_),
    .A2(net2881),
    .Y(_00237_),
    .B1(_00442_));
 sg13g2_mux2_1 _20141_ (.A0(net2279),
    .A1(net2259),
    .S(net2821),
    .X(_00238_));
 sg13g2_mux2_1 _20142_ (.A0(net2277),
    .A1(net2256),
    .S(net2854),
    .X(_00239_));
 sg13g2_nor2_1 _20143_ (.A(net2276),
    .B(net2827),
    .Y(_00444_));
 sg13g2_a21oi_1 _20144_ (.A1(_05847_),
    .A2(net2827),
    .Y(_00240_),
    .B1(_00444_));
 sg13g2_mux2_1 _20145_ (.A0(net324),
    .A1(net2253),
    .S(net2833),
    .X(_00241_));
 sg13g2_mux2_1 _20146_ (.A0(\net.in[209] ),
    .A1(net2251),
    .S(net2860),
    .X(_00242_));
 sg13g2_nand2_1 _20147_ (.Y(_00445_),
    .A(net2249),
    .B(net2835));
 sg13g2_o21ai_1 _20148_ (.B1(_00445_),
    .Y(_00243_),
    .A1(_05935_),
    .A2(net2835));
 sg13g2_mux2_1 _20149_ (.A0(net2269),
    .A1(net2244),
    .S(net2823),
    .X(_00244_));
 sg13g2_nand2_1 _20150_ (.Y(_00446_),
    .A(net2242),
    .B(net2881));
 sg13g2_o21ai_1 _20151_ (.B1(_00446_),
    .Y(_00245_),
    .A1(_05528_),
    .A2(net2881));
 sg13g2_mux2_1 _20152_ (.A0(net2261),
    .A1(net2239),
    .S(net2862),
    .X(_00246_));
 sg13g2_mux2_1 _20153_ (.A0(net2256),
    .A1(\net.in[222] ),
    .S(net2835),
    .X(_00247_));
 sg13g2_nand2_1 _20154_ (.Y(_00448_),
    .A(\net.in[223] ),
    .B(net2826));
 sg13g2_o21ai_1 _20155_ (.B1(_00448_),
    .Y(_00248_),
    .A1(_05847_),
    .A2(net2826));
 sg13g2_mux2_1 _20156_ (.A0(net2254),
    .A1(net288),
    .S(net2874),
    .X(_00249_));
 sg13g2_mux2_1 _20157_ (.A0(net2251),
    .A1(net358),
    .S(net2868),
    .X(_00250_));
 sg13g2_mux2_1 _20158_ (.A0(net2248),
    .A1(net2237),
    .S(net2821),
    .X(_00251_));
 sg13g2_mux2_1 _20159_ (.A0(net2247),
    .A1(net2236),
    .S(net2863),
    .X(_00252_));
 sg13g2_mux2_1 _20160_ (.A0(net2241),
    .A1(net2233),
    .S(net2856),
    .X(_00253_));
 sg13g2_nor2_1 _20161_ (.A(net2240),
    .B(net2864),
    .Y(_00449_));
 sg13g2_a21oi_1 _20162_ (.A1(_05759_),
    .A2(net2863),
    .Y(_00254_),
    .B1(_00449_));
 sg13g2_mux2_1 _20163_ (.A0(net353),
    .A1(net2228),
    .S(net2858),
    .X(_00255_));
 sg13g2_nor2_1 _20164_ (.A(\net.in[223] ),
    .B(net2830),
    .Y(_00451_));
 sg13g2_a21oi_1 _20165_ (.A1(_05517_),
    .A2(net2830),
    .Y(_00256_),
    .B1(_00451_));
 sg13g2_nor2_1 _20166_ (.A(net2874),
    .B(net288),
    .Y(_00452_));
 sg13g2_a21oi_1 _20167_ (.A1(_05704_),
    .A2(net2874),
    .Y(_00257_),
    .B1(_00452_));
 sg13g2_mux2_1 _20168_ (.A0(net358),
    .A1(net2221),
    .S(net2866),
    .X(_00258_));
 sg13g2_nor2_1 _20169_ (.A(net2238),
    .B(net2851),
    .Y(_00453_));
 sg13g2_a21oi_1 _20170_ (.A1(_05132_),
    .A2(net2851),
    .Y(_00259_),
    .B1(_00453_));
 sg13g2_mux2_1 _20171_ (.A0(net2235),
    .A1(net2214),
    .S(net2819),
    .X(_00260_));
 sg13g2_mux2_1 _20172_ (.A0(net2232),
    .A1(net2212),
    .S(net2841),
    .X(_00261_));
 sg13g2_nor2_1 _20173_ (.A(net2230),
    .B(net2828),
    .Y(_00455_));
 sg13g2_a21oi_1 _20174_ (.A1(_05924_),
    .A2(net2828),
    .Y(_00262_),
    .B1(_00455_));
 sg13g2_mux2_1 _20175_ (.A0(net2226),
    .A1(net301),
    .S(net2829),
    .X(_00263_));
 sg13g2_nand2_1 _20176_ (.Y(_00456_),
    .A(net2830),
    .B(net283));
 sg13g2_o21ai_1 _20177_ (.B1(_00456_),
    .Y(_00264_),
    .A1(_05517_),
    .A2(net2830));
 sg13g2_nand2_1 _20178_ (.Y(_00457_),
    .A(net2878),
    .B(net281));
 sg13g2_o21ai_1 _20179_ (.B1(_00457_),
    .Y(_00265_),
    .A1(_05704_),
    .A2(net2878));
 sg13g2_nor2_1 _20180_ (.A(net2221),
    .B(net2865),
    .Y(_00458_));
 sg13g2_a21oi_2 _20181_ (.B1(_00458_),
    .Y(_00266_),
    .A2(net2865),
    .A1(_06034_));
 sg13g2_nand2_1 _20182_ (.Y(_00460_),
    .A(net2208),
    .B(net2851));
 sg13g2_o21ai_1 _20183_ (.B1(_00460_),
    .Y(_00267_),
    .A1(_05132_),
    .A2(net2851));
 sg13g2_mux2_1 _20184_ (.A0(net2216),
    .A1(net2207),
    .S(net2824),
    .X(_00268_));
 sg13g2_nor2_1 _20185_ (.A(net2212),
    .B(net2834),
    .Y(_00461_));
 sg13g2_a21oi_1 _20186_ (.A1(_05737_),
    .A2(net2834),
    .Y(_00269_),
    .B1(_00461_));
 sg13g2_nor2_1 _20187_ (.A(\net.in[237] ),
    .B(net2829),
    .Y(_00462_));
 sg13g2_a21oi_1 _20188_ (.A1(_05550_),
    .A2(net2824),
    .Y(_00270_),
    .B1(_00462_));
 sg13g2_mux2_1 _20189_ (.A0(net301),
    .A1(net2199),
    .S(net2829),
    .X(_00271_));
 sg13g2_nor2_1 _20190_ (.A(net2835),
    .B(net283),
    .Y(_00463_));
 sg13g2_a21oi_1 _20191_ (.A1(_06012_),
    .A2(net2834),
    .Y(_00272_),
    .B1(_00463_));
 sg13g2_nor2_1 _20192_ (.A(net2877),
    .B(net281),
    .Y(_00465_));
 sg13g2_a21oi_1 _20193_ (.A1(_05605_),
    .A2(net2878),
    .Y(_00273_),
    .B1(_00465_));
 sg13g2_nor2_1 _20194_ (.A(net2210),
    .B(net2885),
    .Y(_00466_));
 sg13g2_a21oi_1 _20195_ (.A1(_05396_),
    .A2(net2885),
    .Y(_00274_),
    .B1(_00466_));
 sg13g2_nor2_1 _20196_ (.A(net2208),
    .B(net2884),
    .Y(_00467_));
 sg13g2_a21oi_1 _20197_ (.A1(_05583_),
    .A2(net2884),
    .Y(_00275_),
    .B1(_00467_));
 sg13g2_nor2_1 _20198_ (.A(net2205),
    .B(net2873),
    .Y(_00468_));
 sg13g2_a21oi_1 _20199_ (.A1(_05253_),
    .A2(net2872),
    .Y(_00276_),
    .B1(_00468_));
 sg13g2_nand2_1 _20200_ (.Y(_00469_),
    .A(\net.in[252] ),
    .B(net2835));
 sg13g2_o21ai_1 _20201_ (.B1(_00469_),
    .Y(_00277_),
    .A1(_05737_),
    .A2(net2835));
 sg13g2_nand2_1 _20202_ (.Y(_00471_),
    .A(net300),
    .B(net2824));
 sg13g2_o21ai_1 _20203_ (.B1(_00471_),
    .Y(_00278_),
    .A1(_05550_),
    .A2(net2824));
 sg13g2_dfrbp_1 _20204_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net163),
    .D(_00025_),
    .Q_N(_10094_),
    .Q(\net.in[0] ));
 sg13g2_dfrbp_1 _20205_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net162),
    .D(_00026_),
    .Q_N(_10093_),
    .Q(\net.in[1] ));
 sg13g2_dfrbp_1 _20206_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net161),
    .D(_00027_),
    .Q_N(_10092_),
    .Q(\net.in[2] ));
 sg13g2_dfrbp_1 _20207_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net160),
    .D(_00028_),
    .Q_N(_10091_),
    .Q(\net.in[3] ));
 sg13g2_dfrbp_1 _20208_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net159),
    .D(_00029_),
    .Q_N(_10090_),
    .Q(\net.in[4] ));
 sg13g2_dfrbp_1 _20209_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net158),
    .D(_00030_),
    .Q_N(_10089_),
    .Q(\net.in[5] ));
 sg13g2_dfrbp_1 _20210_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net157),
    .D(_00031_),
    .Q_N(_10088_),
    .Q(\net.in[6] ));
 sg13g2_dfrbp_1 _20211_ (.CLK(clknet_4_5__leaf_clk),
    .RESET_B(net156),
    .D(_00032_),
    .Q_N(_10087_),
    .Q(\net.in[7] ));
 sg13g2_dfrbp_1 _20212_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net155),
    .D(_00033_),
    .Q_N(_10086_),
    .Q(\net.in[8] ));
 sg13g2_dfrbp_1 _20213_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net154),
    .D(_00034_),
    .Q_N(_00011_),
    .Q(\net.in[9] ));
 sg13g2_dfrbp_1 _20214_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net153),
    .D(_00035_),
    .Q_N(_10085_),
    .Q(\net.in[10] ));
 sg13g2_dfrbp_1 _20215_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net152),
    .D(_00036_),
    .Q_N(_10084_),
    .Q(\net.in[11] ));
 sg13g2_dfrbp_1 _20216_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net151),
    .D(_00037_),
    .Q_N(_10083_),
    .Q(\calc_categories[6].sum_bits.popcount128.ad0.genblk1[108].add3.a ));
 sg13g2_dfrbp_1 _20217_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net150),
    .D(_00038_),
    .Q_N(_10082_),
    .Q(\net.in[13] ));
 sg13g2_dfrbp_1 _20218_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net149),
    .D(_00039_),
    .Q_N(_10081_),
    .Q(\net.in[14] ));
 sg13g2_dfrbp_1 _20219_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(net287),
    .Q_N(_10080_),
    .Q(\net.in[15] ));
 sg13g2_dfrbp_1 _20220_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net147),
    .D(_00041_),
    .Q_N(_10079_),
    .Q(\net.in[16] ));
 sg13g2_dfrbp_1 _20221_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net146),
    .D(_00042_),
    .Q_N(_10078_),
    .Q(\net.in[17] ));
 sg13g2_dfrbp_1 _20222_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net145),
    .D(_00043_),
    .Q_N(_10077_),
    .Q(\net.in[18] ));
 sg13g2_dfrbp_1 _20223_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net144),
    .D(_00044_),
    .Q_N(_10076_),
    .Q(\net.in[19] ));
 sg13g2_dfrbp_1 _20224_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net143),
    .D(_00045_),
    .Q_N(_10075_),
    .Q(\net.in[20] ));
 sg13g2_dfrbp_1 _20225_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net142),
    .D(_00046_),
    .Q_N(_10074_),
    .Q(\net.in[21] ));
 sg13g2_dfrbp_1 _20226_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net141),
    .D(_00047_),
    .Q_N(_10073_),
    .Q(\net.in[22] ));
 sg13g2_dfrbp_1 _20227_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net140),
    .D(_00048_),
    .Q_N(_10072_),
    .Q(\net.in[23] ));
 sg13g2_dfrbp_1 _20228_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net139),
    .D(net274),
    .Q_N(_00024_),
    .Q(\net.in[24] ));
 sg13g2_dfrbp_1 _20229_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net138),
    .D(_00050_),
    .Q_N(_10071_),
    .Q(\net.in[25] ));
 sg13g2_dfrbp_1 _20230_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net137),
    .D(_00051_),
    .Q_N(_10070_),
    .Q(\net.in[26] ));
 sg13g2_dfrbp_1 _20231_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net136),
    .D(_00052_),
    .Q_N(_10069_),
    .Q(\net.in[27] ));
 sg13g2_dfrbp_1 _20232_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net135),
    .D(_00053_),
    .Q_N(_10068_),
    .Q(\net.in[28] ));
 sg13g2_dfrbp_1 _20233_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net134),
    .D(_00054_),
    .Q_N(_10067_),
    .Q(\net.in[29] ));
 sg13g2_dfrbp_1 _20234_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net133),
    .D(_00055_),
    .Q_N(_00020_),
    .Q(\net.in[30] ));
 sg13g2_dfrbp_1 _20235_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net132),
    .D(_00056_),
    .Q_N(_10066_),
    .Q(\net.in[31] ));
 sg13g2_dfrbp_1 _20236_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net131),
    .D(_00057_),
    .Q_N(_10065_),
    .Q(\net.in[32] ));
 sg13g2_dfrbp_1 _20237_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net130),
    .D(_00058_),
    .Q_N(_10064_),
    .Q(\net.in[33] ));
 sg13g2_dfrbp_1 _20238_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net129),
    .D(_00059_),
    .Q_N(_10063_),
    .Q(\net.in[34] ));
 sg13g2_dfrbp_1 _20239_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net128),
    .D(_00060_),
    .Q_N(_10062_),
    .Q(\net.in[35] ));
 sg13g2_dfrbp_1 _20240_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net127),
    .D(_00061_),
    .Q_N(_00019_),
    .Q(\net.in[36] ));
 sg13g2_dfrbp_1 _20241_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net126),
    .D(_00062_),
    .Q_N(_10061_),
    .Q(\net.in[37] ));
 sg13g2_dfrbp_1 _20242_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net125),
    .D(_00063_),
    .Q_N(_10060_),
    .Q(\net.in[38] ));
 sg13g2_dfrbp_1 _20243_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net124),
    .D(_00064_),
    .Q_N(_10059_),
    .Q(\net.in[39] ));
 sg13g2_dfrbp_1 _20244_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net123),
    .D(_00065_),
    .Q_N(_10058_),
    .Q(\net.in[40] ));
 sg13g2_dfrbp_1 _20245_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net122),
    .D(_00066_),
    .Q_N(_10057_),
    .Q(\net.in[41] ));
 sg13g2_dfrbp_1 _20246_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net121),
    .D(_00067_),
    .Q_N(_10056_),
    .Q(\net.in[42] ));
 sg13g2_dfrbp_1 _20247_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net120),
    .D(_00068_),
    .Q_N(_10055_),
    .Q(\net.in[43] ));
 sg13g2_dfrbp_1 _20248_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net119),
    .D(_00069_),
    .Q_N(_10054_),
    .Q(\net.in[44] ));
 sg13g2_dfrbp_1 _20249_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net118),
    .D(_00070_),
    .Q_N(_10053_),
    .Q(\net.in[45] ));
 sg13g2_dfrbp_1 _20250_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net117),
    .D(_00071_),
    .Q_N(_10052_),
    .Q(\net.in[46] ));
 sg13g2_dfrbp_1 _20251_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net116),
    .D(net303),
    .Q_N(_10051_),
    .Q(\net.in[47] ));
 sg13g2_dfrbp_1 _20252_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net115),
    .D(net276),
    .Q_N(_10050_),
    .Q(\net.in[48] ));
 sg13g2_dfrbp_1 _20253_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net114),
    .D(_00074_),
    .Q_N(_10049_),
    .Q(\net.in[49] ));
 sg13g2_dfrbp_1 _20254_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net113),
    .D(_00075_),
    .Q_N(_10048_),
    .Q(\net.in[50] ));
 sg13g2_dfrbp_1 _20255_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net112),
    .D(_00076_),
    .Q_N(_00000_),
    .Q(\net.in[51] ));
 sg13g2_dfrbp_1 _20256_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net111),
    .D(_00077_),
    .Q_N(_10047_),
    .Q(\net.in[52] ));
 sg13g2_dfrbp_1 _20257_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net110),
    .D(_00078_),
    .Q_N(_10046_),
    .Q(\net.in[53] ));
 sg13g2_dfrbp_1 _20258_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net109),
    .D(_00079_),
    .Q_N(_10045_),
    .Q(\net.in[54] ));
 sg13g2_dfrbp_1 _20259_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net108),
    .D(_00080_),
    .Q_N(_10044_),
    .Q(\net.in[55] ));
 sg13g2_dfrbp_1 _20260_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net107),
    .D(_00081_),
    .Q_N(_00015_),
    .Q(\net.in[56] ));
 sg13g2_dfrbp_1 _20261_ (.CLK(clknet_4_2__leaf_clk),
    .RESET_B(net106),
    .D(_00082_),
    .Q_N(_10043_),
    .Q(\net.in[57] ));
 sg13g2_dfrbp_1 _20262_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net105),
    .D(_00083_),
    .Q_N(_10042_),
    .Q(\net.in[58] ));
 sg13g2_dfrbp_1 _20263_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net104),
    .D(_00084_),
    .Q_N(_10041_),
    .Q(\net.in[59] ));
 sg13g2_dfrbp_1 _20264_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net103),
    .D(_00085_),
    .Q_N(_10040_),
    .Q(\net.in[60] ));
 sg13g2_dfrbp_1 _20265_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net102),
    .D(_00086_),
    .Q_N(_00008_),
    .Q(\net.in[61] ));
 sg13g2_dfrbp_1 _20266_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net101),
    .D(_00087_),
    .Q_N(_10039_),
    .Q(\net.in[62] ));
 sg13g2_dfrbp_1 _20267_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net100),
    .D(_00088_),
    .Q_N(_10038_),
    .Q(\net.in[63] ));
 sg13g2_dfrbp_1 _20268_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net99),
    .D(_00089_),
    .Q_N(_10037_),
    .Q(\net.in[64] ));
 sg13g2_dfrbp_1 _20269_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net98),
    .D(_00090_),
    .Q_N(_10036_),
    .Q(\net.in[65] ));
 sg13g2_dfrbp_1 _20270_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net97),
    .D(_00091_),
    .Q_N(_10035_),
    .Q(\net.in[66] ));
 sg13g2_dfrbp_1 _20271_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net96),
    .D(_00092_),
    .Q_N(_10034_),
    .Q(\net.in[67] ));
 sg13g2_dfrbp_1 _20272_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net95),
    .D(_00093_),
    .Q_N(_10033_),
    .Q(\net.in[68] ));
 sg13g2_dfrbp_1 _20273_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net94),
    .D(_00094_),
    .Q_N(_10032_),
    .Q(\net.in[69] ));
 sg13g2_dfrbp_1 _20274_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net93),
    .D(_00095_),
    .Q_N(_10031_),
    .Q(\net.in[70] ));
 sg13g2_dfrbp_1 _20275_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net92),
    .D(_00096_),
    .Q_N(_10030_),
    .Q(\net.in[71] ));
 sg13g2_dfrbp_1 _20276_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net91),
    .D(_00097_),
    .Q_N(_10029_),
    .Q(\net.in[72] ));
 sg13g2_dfrbp_1 _20277_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net90),
    .D(_00098_),
    .Q_N(_10028_),
    .Q(\net.in[73] ));
 sg13g2_dfrbp_1 _20278_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net89),
    .D(_00099_),
    .Q_N(_00022_),
    .Q(\net.in[74] ));
 sg13g2_dfrbp_1 _20279_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net88),
    .D(_00100_),
    .Q_N(_10027_),
    .Q(\net.in[75] ));
 sg13g2_dfrbp_1 _20280_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net87),
    .D(_00101_),
    .Q_N(_10026_),
    .Q(\net.in[76] ));
 sg13g2_dfrbp_1 _20281_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net86),
    .D(_00102_),
    .Q_N(_10025_),
    .Q(\net.in[77] ));
 sg13g2_dfrbp_1 _20282_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net85),
    .D(_00103_),
    .Q_N(_10024_),
    .Q(\net.in[78] ));
 sg13g2_dfrbp_1 _20283_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net84),
    .D(_00104_),
    .Q_N(_10023_),
    .Q(\net.in[79] ));
 sg13g2_dfrbp_1 _20284_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net83),
    .D(_00105_),
    .Q_N(_10022_),
    .Q(\net.in[80] ));
 sg13g2_dfrbp_1 _20285_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net82),
    .D(_00106_),
    .Q_N(_10021_),
    .Q(\net.in[81] ));
 sg13g2_dfrbp_1 _20286_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net81),
    .D(_00107_),
    .Q_N(_10020_),
    .Q(\net.in[82] ));
 sg13g2_dfrbp_1 _20287_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net80),
    .D(_00108_),
    .Q_N(_10019_),
    .Q(\net.in[83] ));
 sg13g2_dfrbp_1 _20288_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net79),
    .D(_00109_),
    .Q_N(_10018_),
    .Q(\net.in[84] ));
 sg13g2_dfrbp_1 _20289_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net78),
    .D(_00110_),
    .Q_N(_00003_),
    .Q(\net.in[85] ));
 sg13g2_dfrbp_1 _20290_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net77),
    .D(_00111_),
    .Q_N(_10017_),
    .Q(\net.in[86] ));
 sg13g2_dfrbp_1 _20291_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net76),
    .D(_00112_),
    .Q_N(_10016_),
    .Q(\net.in[87] ));
 sg13g2_dfrbp_1 _20292_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net75),
    .D(_00113_),
    .Q_N(_00001_),
    .Q(\net.in[88] ));
 sg13g2_dfrbp_1 _20293_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net74),
    .D(_00114_),
    .Q_N(_10015_),
    .Q(\net.in[89] ));
 sg13g2_dfrbp_1 _20294_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net73),
    .D(_00115_),
    .Q_N(_00010_),
    .Q(\net.in[90] ));
 sg13g2_dfrbp_1 _20295_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net72),
    .D(_00116_),
    .Q_N(_10014_),
    .Q(\net.in[91] ));
 sg13g2_dfrbp_1 _20296_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net71),
    .D(_00117_),
    .Q_N(_10013_),
    .Q(\net.in[92] ));
 sg13g2_dfrbp_1 _20297_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net70),
    .D(_00118_),
    .Q_N(_10012_),
    .Q(\net.in[93] ));
 sg13g2_dfrbp_1 _20298_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net69),
    .D(_00119_),
    .Q_N(_10011_),
    .Q(\net.in[94] ));
 sg13g2_dfrbp_1 _20299_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net68),
    .D(_00120_),
    .Q_N(_10010_),
    .Q(\net.in[95] ));
 sg13g2_dfrbp_1 _20300_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net67),
    .D(_00121_),
    .Q_N(_10009_),
    .Q(\net.in[96] ));
 sg13g2_dfrbp_1 _20301_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net66),
    .D(_00122_),
    .Q_N(_10008_),
    .Q(\net.in[97] ));
 sg13g2_dfrbp_1 _20302_ (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net65),
    .D(_00123_),
    .Q_N(_00006_),
    .Q(\net.in[98] ));
 sg13g2_dfrbp_1 _20303_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net64),
    .D(_00124_),
    .Q_N(_10007_),
    .Q(\net.in[99] ));
 sg13g2_dfrbp_1 _20304_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net63),
    .D(_00125_),
    .Q_N(_10006_),
    .Q(\net.in[100] ));
 sg13g2_dfrbp_1 _20305_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net62),
    .D(_00126_),
    .Q_N(_10005_),
    .Q(\net.in[101] ));
 sg13g2_dfrbp_1 _20306_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net61),
    .D(_00127_),
    .Q_N(_10004_),
    .Q(\net.in[102] ));
 sg13g2_dfrbp_1 _20307_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net60),
    .D(_00128_),
    .Q_N(_10003_),
    .Q(\net.in[103] ));
 sg13g2_dfrbp_1 _20308_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net59),
    .D(_00129_),
    .Q_N(_10002_),
    .Q(\net.in[104] ));
 sg13g2_dfrbp_1 _20309_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net58),
    .D(_00130_),
    .Q_N(_10001_),
    .Q(\net.in[105] ));
 sg13g2_dfrbp_1 _20310_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net57),
    .D(_00131_),
    .Q_N(_10000_),
    .Q(\net.in[106] ));
 sg13g2_dfrbp_1 _20311_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net56),
    .D(_00132_),
    .Q_N(_09999_),
    .Q(\net.in[107] ));
 sg13g2_dfrbp_1 _20312_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net55),
    .D(_00133_),
    .Q_N(_09998_),
    .Q(\net.in[108] ));
 sg13g2_dfrbp_1 _20313_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net54),
    .D(_00134_),
    .Q_N(_09997_),
    .Q(\net.in[109] ));
 sg13g2_dfrbp_1 _20314_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net53),
    .D(_00135_),
    .Q_N(_00005_),
    .Q(\net.in[110] ));
 sg13g2_dfrbp_1 _20315_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net52),
    .D(_00136_),
    .Q_N(_09996_),
    .Q(\net.in[111] ));
 sg13g2_dfrbp_1 _20316_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net51),
    .D(_00137_),
    .Q_N(_09995_),
    .Q(\net.in[112] ));
 sg13g2_dfrbp_1 _20317_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net50),
    .D(_00138_),
    .Q_N(_09994_),
    .Q(\net.in[113] ));
 sg13g2_dfrbp_1 _20318_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net49),
    .D(_00139_),
    .Q_N(_09993_),
    .Q(\net.in[114] ));
 sg13g2_dfrbp_1 _20319_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net48),
    .D(_00140_),
    .Q_N(_09992_),
    .Q(\net.in[115] ));
 sg13g2_dfrbp_1 _20320_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net47),
    .D(_00141_),
    .Q_N(_09991_),
    .Q(\net.in[116] ));
 sg13g2_dfrbp_1 _20321_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net46),
    .D(_00142_),
    .Q_N(_09990_),
    .Q(\net.in[117] ));
 sg13g2_dfrbp_1 _20322_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net45),
    .D(_00143_),
    .Q_N(_09989_),
    .Q(\net.in[118] ));
 sg13g2_dfrbp_1 _20323_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net44),
    .D(_00144_),
    .Q_N(_09988_),
    .Q(\net.in[119] ));
 sg13g2_dfrbp_1 _20324_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net43),
    .D(_00145_),
    .Q_N(_09987_),
    .Q(\net.in[120] ));
 sg13g2_dfrbp_1 _20325_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net42),
    .D(_00146_),
    .Q_N(_09986_),
    .Q(\net.in[121] ));
 sg13g2_dfrbp_1 _20326_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net41),
    .D(_00147_),
    .Q_N(_09985_),
    .Q(\net.in[122] ));
 sg13g2_dfrbp_1 _20327_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net40),
    .D(_00148_),
    .Q_N(_09984_),
    .Q(\net.in[123] ));
 sg13g2_dfrbp_1 _20328_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net39),
    .D(_00149_),
    .Q_N(_09983_),
    .Q(\net.in[124] ));
 sg13g2_dfrbp_1 _20329_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net38),
    .D(_00150_),
    .Q_N(_09982_),
    .Q(\net.in[125] ));
 sg13g2_dfrbp_1 _20330_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net37),
    .D(_00151_),
    .Q_N(_09981_),
    .Q(\net.in[126] ));
 sg13g2_dfrbp_1 _20331_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net36),
    .D(_00152_),
    .Q_N(_09980_),
    .Q(\net.in[127] ));
 sg13g2_dfrbp_1 _20332_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net35),
    .D(_00153_),
    .Q_N(_09979_),
    .Q(\net.in[128] ));
 sg13g2_dfrbp_1 _20333_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net34),
    .D(_00154_),
    .Q_N(_09978_),
    .Q(\net.in[129] ));
 sg13g2_dfrbp_1 _20334_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net33),
    .D(_00155_),
    .Q_N(_09977_),
    .Q(\net.in[130] ));
 sg13g2_dfrbp_1 _20335_ (.CLK(clknet_4_6__leaf_clk),
    .RESET_B(net32),
    .D(_00156_),
    .Q_N(_09976_),
    .Q(\net.in[131] ));
 sg13g2_dfrbp_1 _20336_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net31),
    .D(_00157_),
    .Q_N(_09975_),
    .Q(\net.in[132] ));
 sg13g2_dfrbp_1 _20337_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net30),
    .D(net327),
    .Q_N(_09974_),
    .Q(\net.in[133] ));
 sg13g2_dfrbp_1 _20338_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net29),
    .D(_00159_),
    .Q_N(_09973_),
    .Q(\net.in[134] ));
 sg13g2_dfrbp_1 _20339_ (.CLK(clknet_4_15__leaf_clk),
    .RESET_B(net28),
    .D(_00160_),
    .Q_N(_09972_),
    .Q(\net.in[135] ));
 sg13g2_dfrbp_1 _20340_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net27),
    .D(_00161_),
    .Q_N(_00004_),
    .Q(\net.in[136] ));
 sg13g2_dfrbp_1 _20341_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net26),
    .D(_00162_),
    .Q_N(_00018_),
    .Q(\net.in[137] ));
 sg13g2_dfrbp_1 _20342_ (.CLK(clknet_4_7__leaf_clk),
    .RESET_B(net25),
    .D(_00163_),
    .Q_N(_00023_),
    .Q(\net.in[138] ));
 sg13g2_dfrbp_1 _20343_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net24),
    .D(_00164_),
    .Q_N(_09971_),
    .Q(\net.in[139] ));
 sg13g2_dfrbp_1 _20344_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net23),
    .D(_00165_),
    .Q_N(_09970_),
    .Q(\net.in[140] ));
 sg13g2_dfrbp_1 _20345_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net22),
    .D(_00166_),
    .Q_N(_09969_),
    .Q(\net.in[141] ));
 sg13g2_dfrbp_1 _20346_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net21),
    .D(_00167_),
    .Q_N(_09968_),
    .Q(\calc_categories[0].sum_bits.popcount128.ad0.genblk1[105].add3.a ));
 sg13g2_dfrbp_1 _20347_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net20),
    .D(_00168_),
    .Q_N(_09967_),
    .Q(\net.in[143] ));
 sg13g2_dfrbp_1 _20348_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net19),
    .D(_00169_),
    .Q_N(_09966_),
    .Q(\net.in[144] ));
 sg13g2_dfrbp_1 _20349_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net18),
    .D(_00170_),
    .Q_N(_09965_),
    .Q(\net.in[145] ));
 sg13g2_dfrbp_1 _20350_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net17),
    .D(net317),
    .Q_N(_09964_),
    .Q(\net.in[146] ));
 sg13g2_dfrbp_1 _20351_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net16),
    .D(_00172_),
    .Q_N(_09963_),
    .Q(\net.in[147] ));
 sg13g2_dfrbp_1 _20352_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net15),
    .D(_00173_),
    .Q_N(_09962_),
    .Q(\net.in[148] ));
 sg13g2_dfrbp_1 _20353_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net14),
    .D(_00174_),
    .Q_N(_09961_),
    .Q(\net.in[149] ));
 sg13g2_dfrbp_1 _20354_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net13),
    .D(_00175_),
    .Q_N(_00002_),
    .Q(\net.in[150] ));
 sg13g2_dfrbp_1 _20355_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net12),
    .D(_00176_),
    .Q_N(_09960_),
    .Q(\net.in[151] ));
 sg13g2_dfrbp_1 _20356_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net265),
    .D(_00177_),
    .Q_N(_00012_),
    .Q(\net.in[152] ));
 sg13g2_dfrbp_1 _20357_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net264),
    .D(_00178_),
    .Q_N(_09959_),
    .Q(\calc_categories[4].sum_bits.popcount128.add3.genblk1[12].add3.c ));
 sg13g2_dfrbp_1 _20358_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net263),
    .D(_00179_),
    .Q_N(_00021_),
    .Q(\net.in[154] ));
 sg13g2_dfrbp_1 _20359_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net262),
    .D(_00180_),
    .Q_N(_09958_),
    .Q(\net.in[155] ));
 sg13g2_dfrbp_1 _20360_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net261),
    .D(_00181_),
    .Q_N(_09957_),
    .Q(\net.in[156] ));
 sg13g2_dfrbp_1 _20361_ (.CLK(clknet_4_9__leaf_clk),
    .RESET_B(net260),
    .D(_00182_),
    .Q_N(_09956_),
    .Q(\net.in[157] ));
 sg13g2_dfrbp_1 _20362_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net259),
    .D(_00183_),
    .Q_N(_09955_),
    .Q(\net.in[158] ));
 sg13g2_dfrbp_1 _20363_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net258),
    .D(_00184_),
    .Q_N(_09954_),
    .Q(\net.in[159] ));
 sg13g2_dfrbp_1 _20364_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net257),
    .D(_00185_),
    .Q_N(_09953_),
    .Q(\net.in[160] ));
 sg13g2_dfrbp_1 _20365_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net256),
    .D(_00186_),
    .Q_N(_09952_),
    .Q(\net.in[161] ));
 sg13g2_dfrbp_1 _20366_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net255),
    .D(_00187_),
    .Q_N(_09951_),
    .Q(\net.in[162] ));
 sg13g2_dfrbp_1 _20367_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net254),
    .D(_00188_),
    .Q_N(_00009_),
    .Q(\net.in[163] ));
 sg13g2_dfrbp_1 _20368_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net253),
    .D(_00189_),
    .Q_N(_09950_),
    .Q(\net.in[164] ));
 sg13g2_dfrbp_1 _20369_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net252),
    .D(_00190_),
    .Q_N(_09949_),
    .Q(\net.in[165] ));
 sg13g2_dfrbp_1 _20370_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net251),
    .D(_00191_),
    .Q_N(_09948_),
    .Q(\net.in[166] ));
 sg13g2_dfrbp_1 _20371_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net250),
    .D(_00192_),
    .Q_N(_09947_),
    .Q(\net.in[167] ));
 sg13g2_dfrbp_1 _20372_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net249),
    .D(_00193_),
    .Q_N(_09946_),
    .Q(\net.in[168] ));
 sg13g2_dfrbp_1 _20373_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net248),
    .D(_00194_),
    .Q_N(_09945_),
    .Q(\net.in[169] ));
 sg13g2_dfrbp_1 _20374_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net247),
    .D(_00195_),
    .Q_N(_09944_),
    .Q(\net.in[170] ));
 sg13g2_dfrbp_1 _20375_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net246),
    .D(_00196_),
    .Q_N(_09943_),
    .Q(\net.in[171] ));
 sg13g2_dfrbp_1 _20376_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net245),
    .D(_00197_),
    .Q_N(_09942_),
    .Q(\net.in[172] ));
 sg13g2_dfrbp_1 _20377_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net244),
    .D(_00198_),
    .Q_N(_09941_),
    .Q(\net.in[173] ));
 sg13g2_dfrbp_1 _20378_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net243),
    .D(_00199_),
    .Q_N(_09940_),
    .Q(\net.in[174] ));
 sg13g2_dfrbp_1 _20379_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net242),
    .D(_00200_),
    .Q_N(_09939_),
    .Q(\net.in[175] ));
 sg13g2_dfrbp_1 _20380_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net241),
    .D(_00201_),
    .Q_N(_09938_),
    .Q(\net.in[176] ));
 sg13g2_dfrbp_1 _20381_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net240),
    .D(_00202_),
    .Q_N(_09937_),
    .Q(\net.in[177] ));
 sg13g2_dfrbp_1 _20382_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net239),
    .D(_00203_),
    .Q_N(_00014_),
    .Q(\net.in[178] ));
 sg13g2_dfrbp_1 _20383_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net238),
    .D(net341),
    .Q_N(_09936_),
    .Q(\net.in[179] ));
 sg13g2_dfrbp_1 _20384_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net237),
    .D(_00205_),
    .Q_N(_09935_),
    .Q(\net.in[180] ));
 sg13g2_dfrbp_1 _20385_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net236),
    .D(_00206_),
    .Q_N(_09934_),
    .Q(\net.in[181] ));
 sg13g2_dfrbp_1 _20386_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net235),
    .D(_00207_),
    .Q_N(_09933_),
    .Q(\net.in[182] ));
 sg13g2_dfrbp_1 _20387_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net234),
    .D(_00208_),
    .Q_N(_09932_),
    .Q(\net.in[183] ));
 sg13g2_dfrbp_1 _20388_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net233),
    .D(_00209_),
    .Q_N(_09931_),
    .Q(\net.in[184] ));
 sg13g2_dfrbp_1 _20389_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net232),
    .D(_00210_),
    .Q_N(_09930_),
    .Q(\net.in[185] ));
 sg13g2_dfrbp_1 _20390_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net231),
    .D(_00211_),
    .Q_N(_09929_),
    .Q(\net.in[186] ));
 sg13g2_dfrbp_1 _20391_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net230),
    .D(_00212_),
    .Q_N(_09928_),
    .Q(\net.in[187] ));
 sg13g2_dfrbp_1 _20392_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net229),
    .D(_00213_),
    .Q_N(_09927_),
    .Q(\net.in[188] ));
 sg13g2_dfrbp_1 _20393_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net228),
    .D(_00214_),
    .Q_N(_09926_),
    .Q(\net.in[189] ));
 sg13g2_dfrbp_1 _20394_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net227),
    .D(_00215_),
    .Q_N(_09925_),
    .Q(\net.in[190] ));
 sg13g2_dfrbp_1 _20395_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net226),
    .D(_00216_),
    .Q_N(_09924_),
    .Q(\net.in[191] ));
 sg13g2_dfrbp_1 _20396_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net225),
    .D(_00217_),
    .Q_N(_09923_),
    .Q(\net.in[192] ));
 sg13g2_dfrbp_1 _20397_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net224),
    .D(_00218_),
    .Q_N(_09922_),
    .Q(\net.in[193] ));
 sg13g2_dfrbp_1 _20398_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net223),
    .D(_00219_),
    .Q_N(_09921_),
    .Q(\net.in[194] ));
 sg13g2_dfrbp_1 _20399_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net222),
    .D(net334),
    .Q_N(_09920_),
    .Q(\net.in[195] ));
 sg13g2_dfrbp_1 _20400_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net221),
    .D(_00221_),
    .Q_N(_09919_),
    .Q(\net.in[196] ));
 sg13g2_dfrbp_1 _20401_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net220),
    .D(_00222_),
    .Q_N(_09918_),
    .Q(\net.in[197] ));
 sg13g2_dfrbp_1 _20402_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net219),
    .D(_00223_),
    .Q_N(_09917_),
    .Q(\net.in[198] ));
 sg13g2_dfrbp_1 _20403_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net218),
    .D(_00224_),
    .Q_N(_09916_),
    .Q(\net.in[199] ));
 sg13g2_dfrbp_1 _20404_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net217),
    .D(net310),
    .Q_N(_09915_),
    .Q(\net.in[200] ));
 sg13g2_dfrbp_1 _20405_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net216),
    .D(net307),
    .Q_N(_09914_),
    .Q(\net.in[201] ));
 sg13g2_dfrbp_1 _20406_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net215),
    .D(_00227_),
    .Q_N(_09913_),
    .Q(\net.in[202] ));
 sg13g2_dfrbp_1 _20407_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net214),
    .D(_00228_),
    .Q_N(_09912_),
    .Q(\net.in[203] ));
 sg13g2_dfrbp_1 _20408_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net213),
    .D(_00229_),
    .Q_N(_09911_),
    .Q(\net.in[204] ));
 sg13g2_dfrbp_1 _20409_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net212),
    .D(_00230_),
    .Q_N(_09910_),
    .Q(\net.in[205] ));
 sg13g2_dfrbp_1 _20410_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net211),
    .D(_00231_),
    .Q_N(_09909_),
    .Q(\net.in[206] ));
 sg13g2_dfrbp_1 _20411_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net210),
    .D(_00232_),
    .Q_N(_09908_),
    .Q(\net.in[207] ));
 sg13g2_dfrbp_1 _20412_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net209),
    .D(_00233_),
    .Q_N(_09907_),
    .Q(\net.in[208] ));
 sg13g2_dfrbp_1 _20413_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net208),
    .D(_00234_),
    .Q_N(_09906_),
    .Q(\net.in[209] ));
 sg13g2_dfrbp_1 _20414_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net207),
    .D(_00235_),
    .Q_N(_00016_),
    .Q(\net.in[210] ));
 sg13g2_dfrbp_1 _20415_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net206),
    .D(_00236_),
    .Q_N(_09905_),
    .Q(\net.in[211] ));
 sg13g2_dfrbp_1 _20416_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net205),
    .D(_00237_),
    .Q_N(_09904_),
    .Q(\net.in[212] ));
 sg13g2_dfrbp_1 _20417_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net204),
    .D(_00238_),
    .Q_N(_09903_),
    .Q(\net.in[213] ));
 sg13g2_dfrbp_1 _20418_ (.CLK(clknet_4_13__leaf_clk),
    .RESET_B(net203),
    .D(_00239_),
    .Q_N(_09902_),
    .Q(\net.in[214] ));
 sg13g2_dfrbp_1 _20419_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net202),
    .D(_00240_),
    .Q_N(_09901_),
    .Q(\net.in[215] ));
 sg13g2_dfrbp_1 _20420_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net201),
    .D(_00241_),
    .Q_N(_09900_),
    .Q(\net.in[216] ));
 sg13g2_dfrbp_1 _20421_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net200),
    .D(_00242_),
    .Q_N(_09899_),
    .Q(\net.in[217] ));
 sg13g2_dfrbp_1 _20422_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net199),
    .D(_00243_),
    .Q_N(_09898_),
    .Q(\net.in[218] ));
 sg13g2_dfrbp_1 _20423_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net198),
    .D(_00244_),
    .Q_N(_09897_),
    .Q(\net.in[219] ));
 sg13g2_dfrbp_1 _20424_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net197),
    .D(_00245_),
    .Q_N(_09896_),
    .Q(\net.in[220] ));
 sg13g2_dfrbp_1 _20425_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net196),
    .D(_00246_),
    .Q_N(_09895_),
    .Q(\net.in[221] ));
 sg13g2_dfrbp_1 _20426_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net195),
    .D(net312),
    .Q_N(_09894_),
    .Q(\net.in[222] ));
 sg13g2_dfrbp_1 _20427_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net194),
    .D(_00248_),
    .Q_N(_09893_),
    .Q(\net.in[223] ));
 sg13g2_dfrbp_1 _20428_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net193),
    .D(_00249_),
    .Q_N(_09892_),
    .Q(\net.in[224] ));
 sg13g2_dfrbp_1 _20429_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net192),
    .D(_00250_),
    .Q_N(_09891_),
    .Q(\net.in[225] ));
 sg13g2_dfrbp_1 _20430_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net191),
    .D(_00251_),
    .Q_N(_09890_),
    .Q(\net.in[226] ));
 sg13g2_dfrbp_1 _20431_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net190),
    .D(net386),
    .Q_N(_00007_),
    .Q(\net.in[227] ));
 sg13g2_dfrbp_1 _20432_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net189),
    .D(_00253_),
    .Q_N(_09889_),
    .Q(\net.in[228] ));
 sg13g2_dfrbp_1 _20433_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net188),
    .D(_00254_),
    .Q_N(_09888_),
    .Q(\net.in[229] ));
 sg13g2_dfrbp_1 _20434_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net187),
    .D(_00255_),
    .Q_N(_09887_),
    .Q(\net.in[230] ));
 sg13g2_dfrbp_1 _20435_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net186),
    .D(_00256_),
    .Q_N(_09886_),
    .Q(\net.in[231] ));
 sg13g2_dfrbp_1 _20436_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net185),
    .D(net289),
    .Q_N(_09885_),
    .Q(\net.in[232] ));
 sg13g2_dfrbp_1 _20437_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net184),
    .D(_00258_),
    .Q_N(_09884_),
    .Q(\net.in[233] ));
 sg13g2_dfrbp_1 _20438_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net183),
    .D(_00259_),
    .Q_N(_09883_),
    .Q(\net.in[234] ));
 sg13g2_dfrbp_1 _20439_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net182),
    .D(_00260_),
    .Q_N(_09882_),
    .Q(\net.in[235] ));
 sg13g2_dfrbp_1 _20440_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net181),
    .D(_00261_),
    .Q_N(_09881_),
    .Q(\net.in[236] ));
 sg13g2_dfrbp_1 _20441_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net180),
    .D(_00262_),
    .Q_N(_09880_),
    .Q(\net.in[237] ));
 sg13g2_dfrbp_1 _20442_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net179),
    .D(_00263_),
    .Q_N(_09879_),
    .Q(\net.in[238] ));
 sg13g2_dfrbp_1 _20443_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net178),
    .D(_00264_),
    .Q_N(_09878_),
    .Q(\net.in[239] ));
 sg13g2_dfrbp_1 _20444_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net177),
    .D(_00265_),
    .Q_N(_09877_),
    .Q(\net.in[240] ));
 sg13g2_dfrbp_1 _20445_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net176),
    .D(_00266_),
    .Q_N(_09876_),
    .Q(\net.in[241] ));
 sg13g2_dfrbp_1 _20446_ (.CLK(clknet_4_8__leaf_clk),
    .RESET_B(net175),
    .D(_00267_),
    .Q_N(_09875_),
    .Q(\net.in[242] ));
 sg13g2_dfrbp_1 _20447_ (.CLK(clknet_4_1__leaf_clk),
    .RESET_B(net174),
    .D(_00268_),
    .Q_N(_09874_),
    .Q(\net.in[243] ));
 sg13g2_dfrbp_1 _20448_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net173),
    .D(_00269_),
    .Q_N(_09873_),
    .Q(\net.in[244] ));
 sg13g2_dfrbp_1 _20449_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net172),
    .D(_00270_),
    .Q_N(_00017_),
    .Q(\net.in[245] ));
 sg13g2_dfrbp_1 _20450_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net171),
    .D(_00271_),
    .Q_N(_09872_),
    .Q(\net.in[246] ));
 sg13g2_dfrbp_1 _20451_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net170),
    .D(_00272_),
    .Q_N(_00013_),
    .Q(\net.in[247] ));
 sg13g2_dfrbp_1 _20452_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net169),
    .D(_00273_),
    .Q_N(_09871_),
    .Q(\net.in[248] ));
 sg13g2_dfrbp_1 _20453_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net168),
    .D(_00274_),
    .Q_N(_09870_),
    .Q(\net.in[249] ));
 sg13g2_dfrbp_1 _20454_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net167),
    .D(_00275_),
    .Q_N(_09869_),
    .Q(\net.in[250] ));
 sg13g2_dfrbp_1 _20455_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net166),
    .D(_00276_),
    .Q_N(_09868_),
    .Q(\net.in[251] ));
 sg13g2_dfrbp_1 _20456_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net165),
    .D(_00277_),
    .Q_N(_09867_),
    .Q(\net.in[252] ));
 sg13g2_dfrbp_1 _20457_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net164),
    .D(_00278_),
    .Q_N(_09866_),
    .Q(\net.in[253] ));
 sg13g2_tiehi _20354__13 (.L_HI(net13));
 sg13g2_tiehi _20353__14 (.L_HI(net14));
 sg13g2_tiehi _20352__15 (.L_HI(net15));
 sg13g2_tiehi _20351__16 (.L_HI(net16));
 sg13g2_tiehi _20350__17 (.L_HI(net17));
 sg13g2_tiehi _20349__18 (.L_HI(net18));
 sg13g2_tiehi _20348__19 (.L_HI(net19));
 sg13g2_tiehi _20347__20 (.L_HI(net20));
 sg13g2_tiehi _20346__21 (.L_HI(net21));
 sg13g2_tiehi _20345__22 (.L_HI(net22));
 sg13g2_tiehi _20344__23 (.L_HI(net23));
 sg13g2_tiehi _20343__24 (.L_HI(net24));
 sg13g2_tiehi _20342__25 (.L_HI(net25));
 sg13g2_tiehi _20341__26 (.L_HI(net26));
 sg13g2_tiehi _20340__27 (.L_HI(net27));
 sg13g2_tiehi _20339__28 (.L_HI(net28));
 sg13g2_tiehi _20338__29 (.L_HI(net29));
 sg13g2_tiehi _20337__30 (.L_HI(net30));
 sg13g2_tiehi _20336__31 (.L_HI(net31));
 sg13g2_tiehi _20335__32 (.L_HI(net32));
 sg13g2_tiehi _20334__33 (.L_HI(net33));
 sg13g2_tiehi _20333__34 (.L_HI(net34));
 sg13g2_tiehi _20332__35 (.L_HI(net35));
 sg13g2_tiehi _20331__36 (.L_HI(net36));
 sg13g2_tiehi _20330__37 (.L_HI(net37));
 sg13g2_tiehi _20329__38 (.L_HI(net38));
 sg13g2_tiehi _20328__39 (.L_HI(net39));
 sg13g2_tiehi _20327__40 (.L_HI(net40));
 sg13g2_tiehi _20326__41 (.L_HI(net41));
 sg13g2_tiehi _20325__42 (.L_HI(net42));
 sg13g2_tiehi _20324__43 (.L_HI(net43));
 sg13g2_tiehi _20323__44 (.L_HI(net44));
 sg13g2_tiehi _20322__45 (.L_HI(net45));
 sg13g2_tiehi _20321__46 (.L_HI(net46));
 sg13g2_tiehi _20320__47 (.L_HI(net47));
 sg13g2_tiehi _20319__48 (.L_HI(net48));
 sg13g2_tiehi _20318__49 (.L_HI(net49));
 sg13g2_tiehi _20317__50 (.L_HI(net50));
 sg13g2_tiehi _20316__51 (.L_HI(net51));
 sg13g2_tiehi _20315__52 (.L_HI(net52));
 sg13g2_tiehi _20314__53 (.L_HI(net53));
 sg13g2_tiehi _20313__54 (.L_HI(net54));
 sg13g2_tiehi _20312__55 (.L_HI(net55));
 sg13g2_tiehi _20311__56 (.L_HI(net56));
 sg13g2_tiehi _20310__57 (.L_HI(net57));
 sg13g2_tiehi _20309__58 (.L_HI(net58));
 sg13g2_tiehi _20308__59 (.L_HI(net59));
 sg13g2_tiehi _20307__60 (.L_HI(net60));
 sg13g2_tiehi _20306__61 (.L_HI(net61));
 sg13g2_tiehi _20305__62 (.L_HI(net62));
 sg13g2_tiehi _20304__63 (.L_HI(net63));
 sg13g2_tiehi _20303__64 (.L_HI(net64));
 sg13g2_tiehi _20302__65 (.L_HI(net65));
 sg13g2_tiehi _20301__66 (.L_HI(net66));
 sg13g2_tiehi _20300__67 (.L_HI(net67));
 sg13g2_tiehi _20299__68 (.L_HI(net68));
 sg13g2_tiehi _20298__69 (.L_HI(net69));
 sg13g2_tiehi _20297__70 (.L_HI(net70));
 sg13g2_tiehi _20296__71 (.L_HI(net71));
 sg13g2_tiehi _20295__72 (.L_HI(net72));
 sg13g2_tiehi _20294__73 (.L_HI(net73));
 sg13g2_tiehi _20293__74 (.L_HI(net74));
 sg13g2_tiehi _20292__75 (.L_HI(net75));
 sg13g2_tiehi _20291__76 (.L_HI(net76));
 sg13g2_tiehi _20290__77 (.L_HI(net77));
 sg13g2_tiehi _20289__78 (.L_HI(net78));
 sg13g2_tiehi _20288__79 (.L_HI(net79));
 sg13g2_tiehi _20287__80 (.L_HI(net80));
 sg13g2_tiehi _20286__81 (.L_HI(net81));
 sg13g2_tiehi _20285__82 (.L_HI(net82));
 sg13g2_tiehi _20284__83 (.L_HI(net83));
 sg13g2_tiehi _20283__84 (.L_HI(net84));
 sg13g2_tiehi _20282__85 (.L_HI(net85));
 sg13g2_tiehi _20281__86 (.L_HI(net86));
 sg13g2_tiehi _20280__87 (.L_HI(net87));
 sg13g2_tiehi _20279__88 (.L_HI(net88));
 sg13g2_tiehi _20278__89 (.L_HI(net89));
 sg13g2_tiehi _20277__90 (.L_HI(net90));
 sg13g2_tiehi _20276__91 (.L_HI(net91));
 sg13g2_tiehi _20275__92 (.L_HI(net92));
 sg13g2_tiehi _20274__93 (.L_HI(net93));
 sg13g2_tiehi _20273__94 (.L_HI(net94));
 sg13g2_tiehi _20272__95 (.L_HI(net95));
 sg13g2_tiehi _20271__96 (.L_HI(net96));
 sg13g2_tiehi _20270__97 (.L_HI(net97));
 sg13g2_tiehi _20269__98 (.L_HI(net98));
 sg13g2_tiehi _20268__99 (.L_HI(net99));
 sg13g2_tiehi _20267__100 (.L_HI(net100));
 sg13g2_tiehi _20266__101 (.L_HI(net101));
 sg13g2_tiehi _20265__102 (.L_HI(net102));
 sg13g2_tiehi _20264__103 (.L_HI(net103));
 sg13g2_tiehi _20263__104 (.L_HI(net104));
 sg13g2_tiehi _20262__105 (.L_HI(net105));
 sg13g2_tiehi _20261__106 (.L_HI(net106));
 sg13g2_tiehi _20260__107 (.L_HI(net107));
 sg13g2_tiehi _20259__108 (.L_HI(net108));
 sg13g2_tiehi _20258__109 (.L_HI(net109));
 sg13g2_tiehi _20257__110 (.L_HI(net110));
 sg13g2_tiehi _20256__111 (.L_HI(net111));
 sg13g2_tiehi _20255__112 (.L_HI(net112));
 sg13g2_tiehi _20254__113 (.L_HI(net113));
 sg13g2_tiehi _20253__114 (.L_HI(net114));
 sg13g2_tiehi _20252__115 (.L_HI(net115));
 sg13g2_tiehi _20251__116 (.L_HI(net116));
 sg13g2_tiehi _20250__117 (.L_HI(net117));
 sg13g2_tiehi _20249__118 (.L_HI(net118));
 sg13g2_tiehi _20248__119 (.L_HI(net119));
 sg13g2_tiehi _20247__120 (.L_HI(net120));
 sg13g2_tiehi _20246__121 (.L_HI(net121));
 sg13g2_tiehi _20245__122 (.L_HI(net122));
 sg13g2_tiehi _20244__123 (.L_HI(net123));
 sg13g2_tiehi _20243__124 (.L_HI(net124));
 sg13g2_tiehi _20242__125 (.L_HI(net125));
 sg13g2_tiehi _20241__126 (.L_HI(net126));
 sg13g2_tiehi _20240__127 (.L_HI(net127));
 sg13g2_tiehi _20239__128 (.L_HI(net128));
 sg13g2_tiehi _20238__129 (.L_HI(net129));
 sg13g2_tiehi _20237__130 (.L_HI(net130));
 sg13g2_tiehi _20236__131 (.L_HI(net131));
 sg13g2_tiehi _20235__132 (.L_HI(net132));
 sg13g2_tiehi _20234__133 (.L_HI(net133));
 sg13g2_tiehi _20233__134 (.L_HI(net134));
 sg13g2_tiehi _20232__135 (.L_HI(net135));
 sg13g2_tiehi _20231__136 (.L_HI(net136));
 sg13g2_tiehi _20230__137 (.L_HI(net137));
 sg13g2_tiehi _20229__138 (.L_HI(net138));
 sg13g2_tiehi _20228__139 (.L_HI(net139));
 sg13g2_tiehi _20227__140 (.L_HI(net140));
 sg13g2_tiehi _20226__141 (.L_HI(net141));
 sg13g2_tiehi _20225__142 (.L_HI(net142));
 sg13g2_tiehi _20224__143 (.L_HI(net143));
 sg13g2_tiehi _20223__144 (.L_HI(net144));
 sg13g2_tiehi _20222__145 (.L_HI(net145));
 sg13g2_tiehi _20221__146 (.L_HI(net146));
 sg13g2_tiehi _20220__147 (.L_HI(net147));
 sg13g2_tiehi _20219__148 (.L_HI(net148));
 sg13g2_tiehi _20218__149 (.L_HI(net149));
 sg13g2_tiehi _20217__150 (.L_HI(net150));
 sg13g2_tiehi _20216__151 (.L_HI(net151));
 sg13g2_tiehi _20215__152 (.L_HI(net152));
 sg13g2_tiehi _20214__153 (.L_HI(net153));
 sg13g2_tiehi _20213__154 (.L_HI(net154));
 sg13g2_tiehi _20212__155 (.L_HI(net155));
 sg13g2_tiehi _20211__156 (.L_HI(net156));
 sg13g2_tiehi _20210__157 (.L_HI(net157));
 sg13g2_tiehi _20209__158 (.L_HI(net158));
 sg13g2_tiehi _20208__159 (.L_HI(net159));
 sg13g2_tiehi _20207__160 (.L_HI(net160));
 sg13g2_tiehi _20206__161 (.L_HI(net161));
 sg13g2_tiehi _20205__162 (.L_HI(net162));
 sg13g2_tiehi _20204__163 (.L_HI(net163));
 sg13g2_tiehi _20457__164 (.L_HI(net164));
 sg13g2_tiehi _20456__165 (.L_HI(net165));
 sg13g2_tiehi _20455__166 (.L_HI(net166));
 sg13g2_tiehi _20454__167 (.L_HI(net167));
 sg13g2_tiehi _20453__168 (.L_HI(net168));
 sg13g2_tiehi _20452__169 (.L_HI(net169));
 sg13g2_tiehi _20451__170 (.L_HI(net170));
 sg13g2_tiehi _20450__171 (.L_HI(net171));
 sg13g2_tiehi _20449__172 (.L_HI(net172));
 sg13g2_tiehi _20448__173 (.L_HI(net173));
 sg13g2_tiehi _20447__174 (.L_HI(net174));
 sg13g2_tiehi _20446__175 (.L_HI(net175));
 sg13g2_tiehi _20445__176 (.L_HI(net176));
 sg13g2_tiehi _20444__177 (.L_HI(net177));
 sg13g2_tiehi _20443__178 (.L_HI(net178));
 sg13g2_tiehi _20442__179 (.L_HI(net179));
 sg13g2_tiehi _20441__180 (.L_HI(net180));
 sg13g2_tiehi _20440__181 (.L_HI(net181));
 sg13g2_tiehi _20439__182 (.L_HI(net182));
 sg13g2_tiehi _20438__183 (.L_HI(net183));
 sg13g2_tiehi _20437__184 (.L_HI(net184));
 sg13g2_tiehi _20436__185 (.L_HI(net185));
 sg13g2_tiehi _20435__186 (.L_HI(net186));
 sg13g2_tiehi _20434__187 (.L_HI(net187));
 sg13g2_tiehi _20433__188 (.L_HI(net188));
 sg13g2_tiehi _20432__189 (.L_HI(net189));
 sg13g2_tiehi _20431__190 (.L_HI(net190));
 sg13g2_tiehi _20430__191 (.L_HI(net191));
 sg13g2_tiehi _20429__192 (.L_HI(net192));
 sg13g2_tiehi _20428__193 (.L_HI(net193));
 sg13g2_tiehi _20427__194 (.L_HI(net194));
 sg13g2_tiehi _20426__195 (.L_HI(net195));
 sg13g2_tiehi _20425__196 (.L_HI(net196));
 sg13g2_tiehi _20424__197 (.L_HI(net197));
 sg13g2_tiehi _20423__198 (.L_HI(net198));
 sg13g2_tiehi _20422__199 (.L_HI(net199));
 sg13g2_tiehi _20421__200 (.L_HI(net200));
 sg13g2_tiehi _20420__201 (.L_HI(net201));
 sg13g2_tiehi _20419__202 (.L_HI(net202));
 sg13g2_tiehi _20418__203 (.L_HI(net203));
 sg13g2_tiehi _20417__204 (.L_HI(net204));
 sg13g2_tiehi _20416__205 (.L_HI(net205));
 sg13g2_tiehi _20415__206 (.L_HI(net206));
 sg13g2_tiehi _20414__207 (.L_HI(net207));
 sg13g2_tiehi _20413__208 (.L_HI(net208));
 sg13g2_tiehi _20412__209 (.L_HI(net209));
 sg13g2_tiehi _20411__210 (.L_HI(net210));
 sg13g2_tiehi _20410__211 (.L_HI(net211));
 sg13g2_tiehi _20409__212 (.L_HI(net212));
 sg13g2_tiehi _20408__213 (.L_HI(net213));
 sg13g2_tiehi _20407__214 (.L_HI(net214));
 sg13g2_tiehi _20406__215 (.L_HI(net215));
 sg13g2_tiehi _20405__216 (.L_HI(net216));
 sg13g2_tiehi _20404__217 (.L_HI(net217));
 sg13g2_tiehi _20403__218 (.L_HI(net218));
 sg13g2_tiehi _20402__219 (.L_HI(net219));
 sg13g2_tiehi _20401__220 (.L_HI(net220));
 sg13g2_tiehi _20400__221 (.L_HI(net221));
 sg13g2_tiehi _20399__222 (.L_HI(net222));
 sg13g2_tiehi _20398__223 (.L_HI(net223));
 sg13g2_tiehi _20397__224 (.L_HI(net224));
 sg13g2_tiehi _20396__225 (.L_HI(net225));
 sg13g2_tiehi _20395__226 (.L_HI(net226));
 sg13g2_tiehi _20394__227 (.L_HI(net227));
 sg13g2_tiehi _20393__228 (.L_HI(net228));
 sg13g2_tiehi _20392__229 (.L_HI(net229));
 sg13g2_tiehi _20391__230 (.L_HI(net230));
 sg13g2_tiehi _20390__231 (.L_HI(net231));
 sg13g2_tiehi _20389__232 (.L_HI(net232));
 sg13g2_tiehi _20388__233 (.L_HI(net233));
 sg13g2_tiehi _20387__234 (.L_HI(net234));
 sg13g2_tiehi _20386__235 (.L_HI(net235));
 sg13g2_tiehi _20385__236 (.L_HI(net236));
 sg13g2_tiehi _20384__237 (.L_HI(net237));
 sg13g2_tiehi _20383__238 (.L_HI(net238));
 sg13g2_tiehi _20382__239 (.L_HI(net239));
 sg13g2_tiehi _20381__240 (.L_HI(net240));
 sg13g2_tiehi _20380__241 (.L_HI(net241));
 sg13g2_tiehi _20379__242 (.L_HI(net242));
 sg13g2_tiehi _20378__243 (.L_HI(net243));
 sg13g2_tiehi _20377__244 (.L_HI(net244));
 sg13g2_tiehi _20376__245 (.L_HI(net245));
 sg13g2_tiehi _20375__246 (.L_HI(net246));
 sg13g2_tiehi _20374__247 (.L_HI(net247));
 sg13g2_tiehi _20373__248 (.L_HI(net248));
 sg13g2_tiehi _20372__249 (.L_HI(net249));
 sg13g2_tiehi _20371__250 (.L_HI(net250));
 sg13g2_tiehi _20370__251 (.L_HI(net251));
 sg13g2_tiehi _20369__252 (.L_HI(net252));
 sg13g2_tiehi _20368__253 (.L_HI(net253));
 sg13g2_tiehi _20367__254 (.L_HI(net254));
 sg13g2_tiehi _20366__255 (.L_HI(net255));
 sg13g2_tiehi _20365__256 (.L_HI(net256));
 sg13g2_tiehi _20364__257 (.L_HI(net257));
 sg13g2_tiehi _20363__258 (.L_HI(net258));
 sg13g2_tiehi _20362__259 (.L_HI(net259));
 sg13g2_tiehi _20361__260 (.L_HI(net260));
 sg13g2_tiehi _20360__261 (.L_HI(net261));
 sg13g2_tiehi _20359__262 (.L_HI(net262));
 sg13g2_tiehi _20358__263 (.L_HI(net263));
 sg13g2_tiehi _20357__264 (.L_HI(net264));
 sg13g2_tiehi _20356__265 (.L_HI(net265));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_266 (.L_HI(net266));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_267 (.L_HI(net267));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_268 (.L_HI(net268));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_269 (.L_HI(net269));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_270 (.L_HI(net270));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_271 (.L_HI(net271));
 sg13g2_tiehi tt_um_rejunity_lgn_mnist_272 (.L_HI(net272));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_rejunity_lgn_mnist_11 (.L_LO(net11));
 sg13g2_tiehi _20355__12 (.L_HI(net12));
 sg13g2_buf_1 _20721_ (.A(net2846),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout2166 (.A(net2167),
    .X(net2166));
 sg13g2_buf_2 fanout2167 (.A(_09827_),
    .X(net2167));
 sg13g2_buf_4 fanout2168 (.X(net2168),
    .A(_09692_));
 sg13g2_buf_2 fanout2169 (.A(_07719_),
    .X(net2169));
 sg13g2_buf_1 fanout2170 (.A(_07719_),
    .X(net2170));
 sg13g2_buf_2 fanout2171 (.A(_07683_),
    .X(net2171));
 sg13g2_buf_1 fanout2172 (.A(_07683_),
    .X(net2172));
 sg13g2_buf_2 fanout2173 (.A(net2174),
    .X(net2173));
 sg13g2_buf_2 fanout2174 (.A(_03801_),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(net2176),
    .X(net2175));
 sg13g2_buf_2 fanout2176 (.A(_03764_),
    .X(net2176));
 sg13g2_buf_16 fanout2177 (.X(net2177),
    .A(_05792_));
 sg13g2_buf_8 fanout2178 (.A(_05385_),
    .X(net2178));
 sg13g2_buf_8 fanout2179 (.A(_05374_),
    .X(net2179));
 sg13g2_buf_8 fanout2180 (.A(_05308_),
    .X(net2180));
 sg13g2_buf_8 fanout2181 (.A(net2182),
    .X(net2181));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(_05198_));
 sg13g2_buf_8 fanout2183 (.A(_05033_),
    .X(net2183));
 sg13g2_buf_8 fanout2184 (.A(_05000_),
    .X(net2184));
 sg13g2_buf_8 fanout2185 (.A(\net.in[251] ),
    .X(net2185));
 sg13g2_buf_8 fanout2186 (.A(net2187),
    .X(net2186));
 sg13g2_buf_16 fanout2187 (.X(net2187),
    .A(\net.in[251] ));
 sg13g2_buf_8 fanout2188 (.A(net2189),
    .X(net2188));
 sg13g2_buf_8 fanout2189 (.A(net349),
    .X(net2189));
 sg13g2_buf_8 fanout2190 (.A(net2193),
    .X(net2190));
 sg13g2_buf_8 fanout2191 (.A(net2193),
    .X(net2191));
 sg13g2_buf_2 fanout2192 (.A(net2193),
    .X(net2192));
 sg13g2_buf_4 fanout2193 (.X(net2193),
    .A(\net.in[249] ));
 sg13g2_buf_8 fanout2194 (.A(net2196),
    .X(net2194));
 sg13g2_buf_4 fanout2195 (.X(net2195),
    .A(net2196));
 sg13g2_buf_8 fanout2196 (.A(net285),
    .X(net2196));
 sg13g2_buf_8 fanout2197 (.A(net2198),
    .X(net2197));
 sg13g2_buf_8 fanout2198 (.A(\net.in[247] ),
    .X(net2198));
 sg13g2_buf_16 fanout2199 (.X(net2199),
    .A(\net.in[246] ));
 sg13g2_buf_8 fanout2200 (.A(net2202),
    .X(net2200));
 sg13g2_buf_8 fanout2201 (.A(net2202),
    .X(net2201));
 sg13g2_buf_8 fanout2202 (.A(\net.in[245] ),
    .X(net2202));
 sg13g2_buf_8 fanout2203 (.A(\net.in[244] ),
    .X(net2203));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(\net.in[244] ));
 sg13g2_buf_4 fanout2205 (.X(net2205),
    .A(net2206));
 sg13g2_buf_4 fanout2206 (.X(net2206),
    .A(net2207));
 sg13g2_buf_8 fanout2207 (.A(net342),
    .X(net2207));
 sg13g2_buf_8 fanout2208 (.A(net2209),
    .X(net2208));
 sg13g2_buf_8 fanout2209 (.A(\net.in[242] ),
    .X(net2209));
 sg13g2_buf_8 fanout2210 (.A(net2211),
    .X(net2210));
 sg13g2_buf_8 fanout2211 (.A(\net.in[241] ),
    .X(net2211));
 sg13g2_buf_8 fanout2212 (.A(net378),
    .X(net2212));
 sg13g2_buf_8 fanout2213 (.A(\net.in[236] ),
    .X(net2213));
 sg13g2_buf_8 fanout2214 (.A(net2216),
    .X(net2214));
 sg13g2_buf_2 fanout2215 (.A(net2216),
    .X(net2215));
 sg13g2_buf_8 fanout2216 (.A(net2217),
    .X(net2216));
 sg13g2_buf_16 fanout2217 (.X(net2217),
    .A(\net.in[235] ));
 sg13g2_buf_16 fanout2218 (.X(net2218),
    .A(\net.in[234] ));
 sg13g2_buf_8 fanout2219 (.A(\net.in[234] ),
    .X(net2219));
 sg13g2_buf_8 fanout2220 (.A(net2221),
    .X(net2220));
 sg13g2_buf_8 fanout2221 (.A(net347),
    .X(net2221));
 sg13g2_buf_8 fanout2222 (.A(net2223),
    .X(net2222));
 sg13g2_buf_8 fanout2223 (.A(\net.in[232] ),
    .X(net2223));
 sg13g2_buf_16 fanout2224 (.X(net2224),
    .A(\net.in[231] ));
 sg13g2_buf_4 fanout2225 (.X(net2225),
    .A(\net.in[231] ));
 sg13g2_buf_8 fanout2226 (.A(net2229),
    .X(net2226));
 sg13g2_buf_8 fanout2227 (.A(net2229),
    .X(net2227));
 sg13g2_buf_4 fanout2228 (.X(net2228),
    .A(net2229));
 sg13g2_buf_2 fanout2229 (.A(\net.in[230] ),
    .X(net2229));
 sg13g2_buf_8 fanout2230 (.A(\net.in[229] ),
    .X(net2230));
 sg13g2_buf_8 fanout2231 (.A(net2234),
    .X(net2231));
 sg13g2_buf_4 fanout2232 (.X(net2232),
    .A(net2234));
 sg13g2_buf_8 fanout2233 (.A(net2234),
    .X(net2233));
 sg13g2_buf_8 fanout2234 (.A(\net.in[228] ),
    .X(net2234));
 sg13g2_buf_8 fanout2235 (.A(\net.in[227] ),
    .X(net2235));
 sg13g2_buf_8 fanout2236 (.A(\net.in[227] ),
    .X(net2236));
 sg13g2_buf_8 fanout2237 (.A(net370),
    .X(net2237));
 sg13g2_buf_8 fanout2238 (.A(net392),
    .X(net2238));
 sg13g2_buf_8 fanout2239 (.A(net348),
    .X(net2239));
 sg13g2_buf_4 fanout2240 (.X(net2240),
    .A(net348));
 sg13g2_buf_8 fanout2241 (.A(net2242),
    .X(net2241));
 sg13g2_buf_8 fanout2242 (.A(net2243),
    .X(net2242));
 sg13g2_buf_4 fanout2243 (.X(net2243),
    .A(\net.in[220] ));
 sg13g2_buf_4 fanout2244 (.X(net2244),
    .A(net2246));
 sg13g2_buf_4 fanout2245 (.X(net2245),
    .A(net2246));
 sg13g2_buf_2 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_16 fanout2247 (.X(net2247),
    .A(net385));
 sg13g2_buf_8 fanout2248 (.A(net2250),
    .X(net2248));
 sg13g2_buf_4 fanout2249 (.X(net2249),
    .A(net2250));
 sg13g2_buf_8 fanout2250 (.A(\net.in[218] ),
    .X(net2250));
 sg13g2_buf_8 fanout2251 (.A(net2252),
    .X(net2251));
 sg13g2_buf_16 fanout2252 (.X(net2252),
    .A(\net.in[217] ));
 sg13g2_buf_8 fanout2253 (.A(net296),
    .X(net2253));
 sg13g2_buf_8 fanout2254 (.A(net296),
    .X(net2254));
 sg13g2_buf_8 fanout2255 (.A(net367),
    .X(net2255));
 sg13g2_buf_8 fanout2256 (.A(net2258),
    .X(net2256));
 sg13g2_buf_8 fanout2257 (.A(net2258),
    .X(net2257));
 sg13g2_buf_8 fanout2258 (.A(net311),
    .X(net2258));
 sg13g2_buf_8 fanout2259 (.A(net2263),
    .X(net2259));
 sg13g2_buf_2 fanout2260 (.A(net2263),
    .X(net2260));
 sg13g2_buf_8 fanout2261 (.A(net2263),
    .X(net2261));
 sg13g2_buf_4 fanout2262 (.X(net2262),
    .A(net2263));
 sg13g2_buf_8 fanout2263 (.A(\net.in[213] ),
    .X(net2263));
 sg13g2_buf_8 fanout2264 (.A(net2268),
    .X(net2264));
 sg13g2_buf_4 fanout2265 (.X(net2265),
    .A(net2268));
 sg13g2_buf_8 fanout2266 (.A(net2268),
    .X(net2266));
 sg13g2_buf_4 fanout2267 (.X(net2267),
    .A(net2268));
 sg13g2_buf_4 fanout2268 (.X(net2268),
    .A(\net.in[212] ));
 sg13g2_buf_4 fanout2269 (.X(net2269),
    .A(net2270));
 sg13g2_buf_8 fanout2270 (.A(net2271),
    .X(net2270));
 sg13g2_buf_8 fanout2271 (.A(\net.in[211] ),
    .X(net2271));
 sg13g2_buf_8 fanout2272 (.A(\net.in[211] ),
    .X(net2272));
 sg13g2_buf_4 fanout2273 (.X(net2273),
    .A(\net.in[211] ));
 sg13g2_buf_8 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_8 fanout2275 (.A(net376),
    .X(net2275));
 sg13g2_buf_8 fanout2276 (.A(net344),
    .X(net2276));
 sg13g2_buf_16 fanout2277 (.X(net2277),
    .A(net374));
 sg13g2_buf_8 fanout2278 (.A(\net.in[206] ),
    .X(net2278));
 sg13g2_buf_16 fanout2279 (.X(net2279),
    .A(\net.in[205] ));
 sg13g2_buf_8 fanout2280 (.A(\net.in[205] ),
    .X(net2280));
 sg13g2_buf_16 fanout2281 (.X(net2281),
    .A(\net.in[204] ));
 sg13g2_buf_8 fanout2282 (.A(net2284),
    .X(net2282));
 sg13g2_buf_8 fanout2283 (.A(net2284),
    .X(net2283));
 sg13g2_buf_8 fanout2284 (.A(\net.in[203] ),
    .X(net2284));
 sg13g2_buf_8 fanout2285 (.A(\net.in[202] ),
    .X(net2285));
 sg13g2_buf_8 fanout2286 (.A(net388),
    .X(net2286));
 sg13g2_buf_8 fanout2287 (.A(net2288),
    .X(net2287));
 sg13g2_buf_8 fanout2288 (.A(\net.in[201] ),
    .X(net2288));
 sg13g2_buf_8 fanout2289 (.A(net2290),
    .X(net2289));
 sg13g2_buf_16 fanout2290 (.X(net2290),
    .A(net309));
 sg13g2_buf_8 fanout2291 (.A(net2294),
    .X(net2291));
 sg13g2_buf_4 fanout2292 (.X(net2292),
    .A(net2294));
 sg13g2_buf_8 fanout2293 (.A(net2294),
    .X(net2293));
 sg13g2_buf_8 fanout2294 (.A(\net.in[199] ),
    .X(net2294));
 sg13g2_buf_8 fanout2295 (.A(\net.in[198] ),
    .X(net2295));
 sg13g2_buf_8 fanout2296 (.A(\net.in[198] ),
    .X(net2296));
 sg13g2_buf_8 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_8 fanout2298 (.A(\net.in[198] ),
    .X(net2298));
 sg13g2_buf_8 fanout2299 (.A(net2301),
    .X(net2299));
 sg13g2_buf_8 fanout2300 (.A(net2301),
    .X(net2300));
 sg13g2_buf_8 fanout2301 (.A(\net.in[197] ),
    .X(net2301));
 sg13g2_buf_8 fanout2302 (.A(net2303),
    .X(net2302));
 sg13g2_buf_8 fanout2303 (.A(\net.in[197] ),
    .X(net2303));
 sg13g2_buf_8 fanout2304 (.A(net2306),
    .X(net2304));
 sg13g2_buf_4 fanout2305 (.X(net2305),
    .A(net2306));
 sg13g2_buf_8 fanout2306 (.A(\net.in[196] ),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(\net.in[196] ),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(\net.in[196] ),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(net333),
    .X(net2309));
 sg13g2_buf_8 fanout2310 (.A(net333),
    .X(net2310));
 sg13g2_buf_4 fanout2311 (.X(net2311),
    .A(net2312));
 sg13g2_buf_2 fanout2312 (.A(net2313),
    .X(net2312));
 sg13g2_buf_8 fanout2313 (.A(\net.in[194] ),
    .X(net2313));
 sg13g2_buf_8 fanout2314 (.A(net2315),
    .X(net2314));
 sg13g2_buf_8 fanout2315 (.A(net319),
    .X(net2315));
 sg13g2_buf_8 fanout2316 (.A(net339),
    .X(net2316));
 sg13g2_buf_4 fanout2317 (.X(net2317),
    .A(\net.in[190] ));
 sg13g2_buf_8 fanout2318 (.A(net2319),
    .X(net2318));
 sg13g2_buf_16 fanout2319 (.X(net2319),
    .A(net305));
 sg13g2_buf_8 fanout2320 (.A(net2321),
    .X(net2320));
 sg13g2_buf_8 fanout2321 (.A(\net.in[188] ),
    .X(net2321));
 sg13g2_buf_8 fanout2322 (.A(net2323),
    .X(net2322));
 sg13g2_buf_16 fanout2323 (.X(net2323),
    .A(\net.in[187] ));
 sg13g2_buf_8 fanout2324 (.A(net2325),
    .X(net2324));
 sg13g2_buf_8 fanout2325 (.A(net2327),
    .X(net2325));
 sg13g2_buf_8 fanout2326 (.A(net2327),
    .X(net2326));
 sg13g2_buf_8 fanout2327 (.A(\net.in[186] ),
    .X(net2327));
 sg13g2_buf_8 fanout2328 (.A(net2329),
    .X(net2328));
 sg13g2_buf_8 fanout2329 (.A(net2331),
    .X(net2329));
 sg13g2_buf_8 fanout2330 (.A(net2331),
    .X(net2330));
 sg13g2_buf_4 fanout2331 (.X(net2331),
    .A(\net.in[185] ));
 sg13g2_buf_8 fanout2332 (.A(net2335),
    .X(net2332));
 sg13g2_buf_8 fanout2333 (.A(net2335),
    .X(net2333));
 sg13g2_buf_2 fanout2334 (.A(net2335),
    .X(net2334));
 sg13g2_buf_8 fanout2335 (.A(\net.in[184] ),
    .X(net2335));
 sg13g2_buf_8 fanout2336 (.A(net2340),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(net2338),
    .X(net2337));
 sg13g2_buf_8 fanout2338 (.A(net2339),
    .X(net2338));
 sg13g2_buf_8 fanout2339 (.A(net2340),
    .X(net2339));
 sg13g2_buf_8 fanout2340 (.A(net366),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(net2344),
    .X(net2341));
 sg13g2_buf_8 fanout2342 (.A(net2343),
    .X(net2342));
 sg13g2_buf_8 fanout2343 (.A(net2344),
    .X(net2343));
 sg13g2_buf_8 fanout2344 (.A(\net.in[182] ),
    .X(net2344));
 sg13g2_buf_8 fanout2345 (.A(net2348),
    .X(net2345));
 sg13g2_buf_8 fanout2346 (.A(net2348),
    .X(net2346));
 sg13g2_buf_4 fanout2347 (.X(net2347),
    .A(net2348));
 sg13g2_buf_8 fanout2348 (.A(\net.in[181] ),
    .X(net2348));
 sg13g2_buf_8 fanout2349 (.A(net2353),
    .X(net2349));
 sg13g2_buf_8 fanout2350 (.A(net2352),
    .X(net2350));
 sg13g2_buf_2 fanout2351 (.A(net2352),
    .X(net2351));
 sg13g2_buf_8 fanout2352 (.A(net2353),
    .X(net2352));
 sg13g2_buf_8 fanout2353 (.A(\net.in[180] ),
    .X(net2353));
 sg13g2_buf_8 fanout2354 (.A(net2355),
    .X(net2354));
 sg13g2_buf_8 fanout2355 (.A(\net.in[179] ),
    .X(net2355));
 sg13g2_buf_8 fanout2356 (.A(\net.in[179] ),
    .X(net2356));
 sg13g2_buf_8 fanout2357 (.A(\net.in[178] ),
    .X(net2357));
 sg13g2_buf_8 fanout2358 (.A(net372),
    .X(net2358));
 sg13g2_buf_4 fanout2359 (.X(net2359),
    .A(net2360));
 sg13g2_buf_8 fanout2360 (.A(\net.in[177] ),
    .X(net2360));
 sg13g2_buf_8 fanout2361 (.A(net322),
    .X(net2361));
 sg13g2_buf_8 fanout2362 (.A(net365),
    .X(net2362));
 sg13g2_buf_8 fanout2363 (.A(net365),
    .X(net2363));
 sg13g2_buf_4 fanout2364 (.X(net2364),
    .A(net2365));
 sg13g2_buf_8 fanout2365 (.A(net2366),
    .X(net2365));
 sg13g2_buf_8 fanout2366 (.A(\net.in[172] ),
    .X(net2366));
 sg13g2_buf_4 fanout2367 (.X(net2367),
    .A(net2368));
 sg13g2_buf_8 fanout2368 (.A(net2369),
    .X(net2368));
 sg13g2_buf_8 fanout2369 (.A(net340),
    .X(net2369));
 sg13g2_buf_8 fanout2370 (.A(net2373),
    .X(net2370));
 sg13g2_buf_2 fanout2371 (.A(net2373),
    .X(net2371));
 sg13g2_buf_8 fanout2372 (.A(net2373),
    .X(net2372));
 sg13g2_buf_8 fanout2373 (.A(\net.in[170] ),
    .X(net2373));
 sg13g2_buf_4 fanout2374 (.X(net2374),
    .A(\net.in[170] ));
 sg13g2_buf_4 fanout2375 (.X(net2375),
    .A(\net.in[170] ));
 sg13g2_buf_16 fanout2376 (.X(net2376),
    .A(\net.in[169] ));
 sg13g2_buf_8 fanout2377 (.A(\net.in[169] ),
    .X(net2377));
 sg13g2_buf_8 fanout2378 (.A(net2379),
    .X(net2378));
 sg13g2_buf_8 fanout2379 (.A(net2380),
    .X(net2379));
 sg13g2_buf_8 fanout2380 (.A(\net.in[168] ),
    .X(net2380));
 sg13g2_buf_4 fanout2381 (.X(net2381),
    .A(net2382));
 sg13g2_buf_8 fanout2382 (.A(\net.in[167] ),
    .X(net2382));
 sg13g2_buf_8 fanout2383 (.A(\net.in[167] ),
    .X(net2383));
 sg13g2_buf_8 fanout2384 (.A(\net.in[167] ),
    .X(net2384));
 sg13g2_buf_4 fanout2385 (.X(net2385),
    .A(net2386));
 sg13g2_buf_4 fanout2386 (.X(net2386),
    .A(net2387));
 sg13g2_buf_4 fanout2387 (.X(net2387),
    .A(net2388));
 sg13g2_buf_8 fanout2388 (.A(\net.in[166] ),
    .X(net2388));
 sg13g2_buf_8 fanout2389 (.A(net2392),
    .X(net2389));
 sg13g2_buf_8 fanout2390 (.A(net2392),
    .X(net2390));
 sg13g2_buf_8 fanout2391 (.A(net2392),
    .X(net2391));
 sg13g2_buf_8 fanout2392 (.A(\net.in[165] ),
    .X(net2392));
 sg13g2_buf_8 fanout2393 (.A(net2396),
    .X(net2393));
 sg13g2_buf_4 fanout2394 (.X(net2394),
    .A(net2396));
 sg13g2_buf_8 fanout2395 (.A(net2396),
    .X(net2395));
 sg13g2_buf_16 fanout2396 (.X(net2396),
    .A(\net.in[164] ));
 sg13g2_buf_8 fanout2397 (.A(\net.in[163] ),
    .X(net2397));
 sg13g2_buf_4 fanout2398 (.X(net2398),
    .A(\net.in[163] ));
 sg13g2_buf_8 fanout2399 (.A(net2400),
    .X(net2399));
 sg13g2_buf_8 fanout2400 (.A(net351),
    .X(net2400));
 sg13g2_buf_8 fanout2401 (.A(net2403),
    .X(net2401));
 sg13g2_buf_4 fanout2402 (.X(net2402),
    .A(net2403));
 sg13g2_buf_16 fanout2403 (.X(net2403),
    .A(net360));
 sg13g2_buf_8 fanout2404 (.A(net379),
    .X(net2404));
 sg13g2_buf_8 fanout2405 (.A(net2406),
    .X(net2405));
 sg13g2_buf_8 fanout2406 (.A(net328),
    .X(net2406));
 sg13g2_buf_4 fanout2407 (.X(net2407),
    .A(net2408));
 sg13g2_buf_16 fanout2408 (.X(net2408),
    .A(net314));
 sg13g2_buf_8 fanout2409 (.A(net2411),
    .X(net2409));
 sg13g2_buf_2 fanout2410 (.A(net2411),
    .X(net2410));
 sg13g2_buf_8 fanout2411 (.A(\net.in[156] ),
    .X(net2411));
 sg13g2_buf_8 fanout2412 (.A(net2414),
    .X(net2412));
 sg13g2_buf_2 fanout2413 (.A(net2414),
    .X(net2413));
 sg13g2_buf_16 fanout2414 (.X(net2414),
    .A(net377));
 sg13g2_buf_4 fanout2415 (.X(net2415),
    .A(net2416));
 sg13g2_buf_8 fanout2416 (.A(\net.in[154] ),
    .X(net2416));
 sg13g2_buf_8 fanout2417 (.A(\net.in[154] ),
    .X(net2417));
 sg13g2_buf_8 fanout2418 (.A(net2421),
    .X(net2418));
 sg13g2_buf_8 fanout2419 (.A(net2421),
    .X(net2419));
 sg13g2_buf_4 fanout2420 (.X(net2420),
    .A(net2421));
 sg13g2_buf_8 fanout2421 (.A(\calc_categories[4].sum_bits.popcount128.add3.genblk1[12].add3.c ),
    .X(net2421));
 sg13g2_buf_8 fanout2422 (.A(\net.in[152] ),
    .X(net2422));
 sg13g2_buf_4 fanout2423 (.X(net2423),
    .A(net2424));
 sg13g2_buf_8 fanout2424 (.A(\net.in[152] ),
    .X(net2424));
 sg13g2_buf_8 fanout2425 (.A(net2426),
    .X(net2425));
 sg13g2_buf_8 fanout2426 (.A(net2429),
    .X(net2426));
 sg13g2_buf_8 fanout2427 (.A(net2429),
    .X(net2427));
 sg13g2_buf_8 fanout2428 (.A(net2429),
    .X(net2428));
 sg13g2_buf_8 fanout2429 (.A(\net.in[151] ),
    .X(net2429));
 sg13g2_buf_8 fanout2430 (.A(net2433),
    .X(net2430));
 sg13g2_buf_4 fanout2431 (.X(net2431),
    .A(net2433));
 sg13g2_buf_8 fanout2432 (.A(net2433),
    .X(net2432));
 sg13g2_buf_8 fanout2433 (.A(\net.in[150] ),
    .X(net2433));
 sg13g2_buf_8 fanout2434 (.A(net2436),
    .X(net2434));
 sg13g2_buf_4 fanout2435 (.X(net2435),
    .A(net2436));
 sg13g2_buf_16 fanout2436 (.X(net2436),
    .A(\net.in[149] ));
 sg13g2_buf_8 fanout2437 (.A(net2441),
    .X(net2437));
 sg13g2_buf_4 fanout2438 (.X(net2438),
    .A(net2441));
 sg13g2_buf_8 fanout2439 (.A(net2441),
    .X(net2439));
 sg13g2_buf_4 fanout2440 (.X(net2440),
    .A(net2441));
 sg13g2_buf_8 fanout2441 (.A(\net.in[148] ),
    .X(net2441));
 sg13g2_buf_16 fanout2442 (.X(net2442),
    .A(net2444));
 sg13g2_buf_8 fanout2443 (.A(net2444),
    .X(net2443));
 sg13g2_buf_4 fanout2444 (.X(net2444),
    .A(\net.in[147] ));
 sg13g2_buf_4 fanout2445 (.X(net2445),
    .A(net2447));
 sg13g2_buf_4 fanout2446 (.X(net2446),
    .A(net2447));
 sg13g2_buf_16 fanout2447 (.X(net2447),
    .A(\net.in[146] ));
 sg13g2_buf_8 fanout2448 (.A(net2450),
    .X(net2448));
 sg13g2_buf_2 fanout2449 (.A(net2450),
    .X(net2449));
 sg13g2_buf_4 fanout2450 (.X(net2450),
    .A(net2451));
 sg13g2_buf_8 fanout2451 (.A(\net.in[143] ),
    .X(net2451));
 sg13g2_buf_8 fanout2452 (.A(net389),
    .X(net2452));
 sg13g2_buf_4 fanout2453 (.X(net2453),
    .A(net2454));
 sg13g2_buf_8 fanout2454 (.A(net2456),
    .X(net2454));
 sg13g2_buf_8 fanout2455 (.A(net2456),
    .X(net2455));
 sg13g2_buf_8 fanout2456 (.A(\net.in[141] ),
    .X(net2456));
 sg13g2_buf_8 fanout2457 (.A(net2458),
    .X(net2457));
 sg13g2_buf_8 fanout2458 (.A(\net.in[140] ),
    .X(net2458));
 sg13g2_buf_8 fanout2459 (.A(\net.in[140] ),
    .X(net2459));
 sg13g2_buf_8 fanout2460 (.A(net2462),
    .X(net2460));
 sg13g2_buf_2 fanout2461 (.A(net2462),
    .X(net2461));
 sg13g2_buf_8 fanout2462 (.A(\net.in[139] ),
    .X(net2462));
 sg13g2_buf_8 fanout2463 (.A(net2466),
    .X(net2463));
 sg13g2_buf_8 fanout2464 (.A(net2465),
    .X(net2464));
 sg13g2_buf_8 fanout2465 (.A(net2466),
    .X(net2465));
 sg13g2_buf_4 fanout2466 (.X(net2466),
    .A(net316));
 sg13g2_buf_8 fanout2467 (.A(\net.in[137] ),
    .X(net2467));
 sg13g2_buf_4 fanout2468 (.X(net2468),
    .A(\net.in[137] ));
 sg13g2_buf_8 fanout2469 (.A(net2470),
    .X(net2469));
 sg13g2_buf_8 fanout2470 (.A(\net.in[137] ),
    .X(net2470));
 sg13g2_buf_16 fanout2471 (.X(net2471),
    .A(\net.in[136] ));
 sg13g2_buf_8 fanout2472 (.A(\net.in[136] ),
    .X(net2472));
 sg13g2_buf_8 fanout2473 (.A(net2477),
    .X(net2473));
 sg13g2_buf_8 fanout2474 (.A(net2476),
    .X(net2474));
 sg13g2_buf_8 fanout2475 (.A(net2476),
    .X(net2475));
 sg13g2_buf_8 fanout2476 (.A(net2477),
    .X(net2476));
 sg13g2_buf_8 fanout2477 (.A(net373),
    .X(net2477));
 sg13g2_buf_8 fanout2478 (.A(net2479),
    .X(net2478));
 sg13g2_buf_4 fanout2479 (.X(net2479),
    .A(net2480));
 sg13g2_buf_8 fanout2480 (.A(net355),
    .X(net2480));
 sg13g2_buf_8 fanout2481 (.A(\net.in[134] ),
    .X(net2481));
 sg13g2_buf_8 fanout2482 (.A(net2483),
    .X(net2482));
 sg13g2_buf_8 fanout2483 (.A(\net.in[133] ),
    .X(net2483));
 sg13g2_buf_8 fanout2484 (.A(\net.in[132] ),
    .X(net2484));
 sg13g2_buf_4 fanout2485 (.X(net2485),
    .A(\net.in[132] ));
 sg13g2_buf_8 fanout2486 (.A(net2487),
    .X(net2486));
 sg13g2_buf_16 fanout2487 (.X(net2487),
    .A(\net.in[132] ));
 sg13g2_buf_8 fanout2488 (.A(net2491),
    .X(net2488));
 sg13g2_buf_4 fanout2489 (.X(net2489),
    .A(net2491));
 sg13g2_buf_8 fanout2490 (.A(net2491),
    .X(net2490));
 sg13g2_buf_8 fanout2491 (.A(net308),
    .X(net2491));
 sg13g2_buf_8 fanout2492 (.A(\net.in[130] ),
    .X(net2492));
 sg13g2_buf_4 fanout2493 (.X(net2493),
    .A(\net.in[130] ));
 sg13g2_buf_8 fanout2494 (.A(net2495),
    .X(net2494));
 sg13g2_buf_8 fanout2495 (.A(\net.in[130] ),
    .X(net2495));
 sg13g2_buf_16 fanout2496 (.X(net2496),
    .A(\net.in[129] ));
 sg13g2_buf_8 fanout2497 (.A(net343),
    .X(net2497));
 sg13g2_buf_8 fanout2498 (.A(\net.in[126] ),
    .X(net2498));
 sg13g2_buf_8 fanout2499 (.A(\net.in[126] ),
    .X(net2499));
 sg13g2_buf_8 fanout2500 (.A(net2501),
    .X(net2500));
 sg13g2_buf_16 fanout2501 (.X(net2501),
    .A(net326));
 sg13g2_buf_4 fanout2502 (.X(net2502),
    .A(net2504));
 sg13g2_buf_2 fanout2503 (.A(net2504),
    .X(net2503));
 sg13g2_buf_16 fanout2504 (.X(net2504),
    .A(\net.in[124] ));
 sg13g2_buf_4 fanout2505 (.X(net2505),
    .A(\net.in[123] ));
 sg13g2_buf_4 fanout2506 (.X(net2506),
    .A(\net.in[123] ));
 sg13g2_buf_8 fanout2507 (.A(net2508),
    .X(net2507));
 sg13g2_buf_8 fanout2508 (.A(\net.in[123] ),
    .X(net2508));
 sg13g2_buf_8 fanout2509 (.A(\net.in[122] ),
    .X(net2509));
 sg13g2_buf_2 fanout2510 (.A(\net.in[122] ),
    .X(net2510));
 sg13g2_buf_4 fanout2511 (.X(net2511),
    .A(net2512));
 sg13g2_buf_8 fanout2512 (.A(\net.in[122] ),
    .X(net2512));
 sg13g2_buf_8 fanout2513 (.A(net2516),
    .X(net2513));
 sg13g2_buf_8 fanout2514 (.A(net2515),
    .X(net2514));
 sg13g2_buf_8 fanout2515 (.A(net2516),
    .X(net2515));
 sg13g2_buf_8 fanout2516 (.A(net387),
    .X(net2516));
 sg13g2_buf_8 fanout2517 (.A(net2520),
    .X(net2517));
 sg13g2_buf_8 fanout2518 (.A(net2519),
    .X(net2518));
 sg13g2_buf_8 fanout2519 (.A(net2520),
    .X(net2519));
 sg13g2_buf_8 fanout2520 (.A(\net.in[120] ),
    .X(net2520));
 sg13g2_buf_16 fanout2521 (.X(net2521),
    .A(net2524));
 sg13g2_buf_8 fanout2522 (.A(net2523),
    .X(net2522));
 sg13g2_buf_8 fanout2523 (.A(net2524),
    .X(net2523));
 sg13g2_buf_8 fanout2524 (.A(\net.in[119] ),
    .X(net2524));
 sg13g2_buf_4 fanout2525 (.X(net2525),
    .A(net2526));
 sg13g2_buf_8 fanout2526 (.A(\net.in[118] ),
    .X(net2526));
 sg13g2_buf_8 fanout2527 (.A(net2529),
    .X(net2527));
 sg13g2_buf_4 fanout2528 (.X(net2528),
    .A(net2529));
 sg13g2_buf_8 fanout2529 (.A(\net.in[118] ),
    .X(net2529));
 sg13g2_buf_8 fanout2530 (.A(net2533),
    .X(net2530));
 sg13g2_buf_8 fanout2531 (.A(net2532),
    .X(net2531));
 sg13g2_buf_8 fanout2532 (.A(net2533),
    .X(net2532));
 sg13g2_buf_8 fanout2533 (.A(\net.in[117] ),
    .X(net2533));
 sg13g2_buf_8 fanout2534 (.A(net2535),
    .X(net2534));
 sg13g2_buf_8 fanout2535 (.A(\net.in[116] ),
    .X(net2535));
 sg13g2_buf_8 fanout2536 (.A(net2538),
    .X(net2536));
 sg13g2_buf_2 fanout2537 (.A(net2538),
    .X(net2537));
 sg13g2_buf_8 fanout2538 (.A(\net.in[116] ),
    .X(net2538));
 sg13g2_buf_8 fanout2539 (.A(net2543),
    .X(net2539));
 sg13g2_buf_4 fanout2540 (.X(net2540),
    .A(net2541));
 sg13g2_buf_2 fanout2541 (.A(net2542),
    .X(net2541));
 sg13g2_buf_4 fanout2542 (.X(net2542),
    .A(net2543));
 sg13g2_buf_4 fanout2543 (.X(net2543),
    .A(\net.in[115] ));
 sg13g2_buf_4 fanout2544 (.X(net2544),
    .A(net2546));
 sg13g2_buf_4 fanout2545 (.X(net2545),
    .A(net2546));
 sg13g2_buf_8 fanout2546 (.A(net323),
    .X(net2546));
 sg13g2_buf_8 fanout2547 (.A(net391),
    .X(net2547));
 sg13g2_buf_8 fanout2548 (.A(net2549),
    .X(net2548));
 sg13g2_buf_8 fanout2549 (.A(\net.in[113] ),
    .X(net2549));
 sg13g2_buf_16 fanout2550 (.X(net2550),
    .A(net364));
 sg13g2_buf_4 fanout2551 (.X(net2551),
    .A(net390));
 sg13g2_buf_8 fanout2552 (.A(\net.in[110] ),
    .X(net2552));
 sg13g2_buf_8 fanout2553 (.A(net2555),
    .X(net2553));
 sg13g2_buf_8 fanout2554 (.A(net2555),
    .X(net2554));
 sg13g2_buf_8 fanout2555 (.A(\net.in[109] ),
    .X(net2555));
 sg13g2_buf_8 fanout2556 (.A(net2557),
    .X(net2556));
 sg13g2_buf_8 fanout2557 (.A(\net.in[108] ),
    .X(net2557));
 sg13g2_buf_8 fanout2558 (.A(net2561),
    .X(net2558));
 sg13g2_buf_2 fanout2559 (.A(net2561),
    .X(net2559));
 sg13g2_buf_8 fanout2560 (.A(net2561),
    .X(net2560));
 sg13g2_buf_8 fanout2561 (.A(\net.in[107] ),
    .X(net2561));
 sg13g2_buf_8 fanout2562 (.A(net2565),
    .X(net2562));
 sg13g2_buf_8 fanout2563 (.A(net2565),
    .X(net2563));
 sg13g2_buf_4 fanout2564 (.X(net2564),
    .A(net2565));
 sg13g2_buf_8 fanout2565 (.A(\net.in[106] ),
    .X(net2565));
 sg13g2_buf_8 fanout2566 (.A(net2569),
    .X(net2566));
 sg13g2_buf_4 fanout2567 (.X(net2567),
    .A(net2569));
 sg13g2_buf_8 fanout2568 (.A(net2569),
    .X(net2568));
 sg13g2_buf_8 fanout2569 (.A(\net.in[105] ),
    .X(net2569));
 sg13g2_buf_4 fanout2570 (.X(net2570),
    .A(net2571));
 sg13g2_buf_8 fanout2571 (.A(net2572),
    .X(net2571));
 sg13g2_buf_8 fanout2572 (.A(net2574),
    .X(net2572));
 sg13g2_buf_8 fanout2573 (.A(net2574),
    .X(net2573));
 sg13g2_buf_4 fanout2574 (.X(net2574),
    .A(\net.in[104] ));
 sg13g2_buf_8 fanout2575 (.A(\net.in[103] ),
    .X(net2575));
 sg13g2_buf_8 fanout2576 (.A(\net.in[103] ),
    .X(net2576));
 sg13g2_buf_8 fanout2577 (.A(net2580),
    .X(net2577));
 sg13g2_buf_8 fanout2578 (.A(net2580),
    .X(net2578));
 sg13g2_buf_4 fanout2579 (.X(net2579),
    .A(net2580));
 sg13g2_buf_2 fanout2580 (.A(\net.in[103] ),
    .X(net2580));
 sg13g2_buf_8 fanout2581 (.A(net2585),
    .X(net2581));
 sg13g2_buf_4 fanout2582 (.X(net2582),
    .A(net2585));
 sg13g2_buf_8 fanout2583 (.A(net2585),
    .X(net2583));
 sg13g2_buf_4 fanout2584 (.X(net2584),
    .A(net2585));
 sg13g2_buf_8 fanout2585 (.A(\net.in[102] ),
    .X(net2585));
 sg13g2_buf_8 fanout2586 (.A(net2591),
    .X(net2586));
 sg13g2_buf_4 fanout2587 (.X(net2587),
    .A(net2588));
 sg13g2_buf_4 fanout2588 (.X(net2588),
    .A(net2591));
 sg13g2_buf_8 fanout2589 (.A(net2590),
    .X(net2589));
 sg13g2_buf_8 fanout2590 (.A(net2591),
    .X(net2590));
 sg13g2_buf_8 fanout2591 (.A(\net.in[101] ),
    .X(net2591));
 sg13g2_buf_16 fanout2592 (.X(net2592),
    .A(net2595));
 sg13g2_buf_4 fanout2593 (.X(net2593),
    .A(net2594));
 sg13g2_buf_8 fanout2594 (.A(net2595),
    .X(net2594));
 sg13g2_buf_8 fanout2595 (.A(net362),
    .X(net2595));
 sg13g2_buf_8 fanout2596 (.A(\net.in[99] ),
    .X(net2596));
 sg13g2_buf_8 fanout2597 (.A(\net.in[99] ),
    .X(net2597));
 sg13g2_buf_8 fanout2598 (.A(net2599),
    .X(net2598));
 sg13g2_buf_16 fanout2599 (.X(net2599),
    .A(\net.in[99] ));
 sg13g2_buf_8 fanout2600 (.A(\net.in[98] ),
    .X(net2600));
 sg13g2_buf_2 fanout2601 (.A(\net.in[98] ),
    .X(net2601));
 sg13g2_buf_8 fanout2602 (.A(\net.in[98] ),
    .X(net2602));
 sg13g2_buf_8 fanout2603 (.A(net368),
    .X(net2603));
 sg13g2_buf_4 fanout2604 (.X(net2604),
    .A(net2605));
 sg13g2_buf_16 fanout2605 (.X(net2605),
    .A(\net.in[95] ));
 sg13g2_buf_8 fanout2606 (.A(net2608),
    .X(net2606));
 sg13g2_buf_8 fanout2607 (.A(net2608),
    .X(net2607));
 sg13g2_buf_8 fanout2608 (.A(net336),
    .X(net2608));
 sg13g2_buf_8 fanout2609 (.A(net2613),
    .X(net2609));
 sg13g2_buf_4 fanout2610 (.X(net2610),
    .A(net2611));
 sg13g2_buf_2 fanout2611 (.A(net2612),
    .X(net2611));
 sg13g2_buf_4 fanout2612 (.X(net2612),
    .A(net2613));
 sg13g2_buf_2 fanout2613 (.A(net350),
    .X(net2613));
 sg13g2_buf_8 fanout2614 (.A(net2615),
    .X(net2614));
 sg13g2_buf_4 fanout2615 (.X(net2615),
    .A(net375));
 sg13g2_buf_8 fanout2616 (.A(net2617),
    .X(net2616));
 sg13g2_buf_8 fanout2617 (.A(\net.in[92] ),
    .X(net2617));
 sg13g2_buf_16 fanout2618 (.X(net2618),
    .A(net2622));
 sg13g2_buf_8 fanout2619 (.A(net2621),
    .X(net2619));
 sg13g2_buf_2 fanout2620 (.A(net2621),
    .X(net2620));
 sg13g2_buf_8 fanout2621 (.A(net2622),
    .X(net2621));
 sg13g2_buf_4 fanout2622 (.X(net2622),
    .A(\net.in[91] ));
 sg13g2_buf_8 fanout2623 (.A(net2625),
    .X(net2623));
 sg13g2_buf_4 fanout2624 (.X(net2624),
    .A(net2625));
 sg13g2_buf_4 fanout2625 (.X(net2625),
    .A(\net.in[90] ));
 sg13g2_buf_4 fanout2626 (.X(net2626),
    .A(net2627));
 sg13g2_buf_4 fanout2627 (.X(net2627),
    .A(net2628));
 sg13g2_buf_8 fanout2628 (.A(net356),
    .X(net2628));
 sg13g2_buf_8 fanout2629 (.A(net2633),
    .X(net2629));
 sg13g2_buf_8 fanout2630 (.A(net2633),
    .X(net2630));
 sg13g2_buf_8 fanout2631 (.A(net2633),
    .X(net2631));
 sg13g2_buf_4 fanout2632 (.X(net2632),
    .A(net2633));
 sg13g2_buf_4 fanout2633 (.X(net2633),
    .A(\net.in[89] ));
 sg13g2_buf_8 fanout2634 (.A(net2637),
    .X(net2634));
 sg13g2_buf_8 fanout2635 (.A(net2637),
    .X(net2635));
 sg13g2_buf_8 fanout2636 (.A(net2637),
    .X(net2636));
 sg13g2_buf_8 fanout2637 (.A(\net.in[88] ),
    .X(net2637));
 sg13g2_buf_8 fanout2638 (.A(net2641),
    .X(net2638));
 sg13g2_buf_4 fanout2639 (.X(net2639),
    .A(net2641));
 sg13g2_buf_8 fanout2640 (.A(net2641),
    .X(net2640));
 sg13g2_buf_8 fanout2641 (.A(\net.in[87] ),
    .X(net2641));
 sg13g2_buf_8 fanout2642 (.A(net2645),
    .X(net2642));
 sg13g2_buf_4 fanout2643 (.X(net2643),
    .A(net2645));
 sg13g2_buf_8 fanout2644 (.A(net2645),
    .X(net2644));
 sg13g2_buf_8 fanout2645 (.A(\net.in[86] ),
    .X(net2645));
 sg13g2_buf_8 fanout2646 (.A(\net.in[85] ),
    .X(net2646));
 sg13g2_buf_4 fanout2647 (.X(net2647),
    .A(\net.in[85] ));
 sg13g2_buf_8 fanout2648 (.A(net2649),
    .X(net2648));
 sg13g2_buf_8 fanout2649 (.A(\net.in[85] ),
    .X(net2649));
 sg13g2_buf_8 fanout2650 (.A(net2651),
    .X(net2650));
 sg13g2_buf_16 fanout2651 (.X(net2651),
    .A(\net.in[84] ));
 sg13g2_buf_8 fanout2652 (.A(net2655),
    .X(net2652));
 sg13g2_buf_8 fanout2653 (.A(net2654),
    .X(net2653));
 sg13g2_buf_8 fanout2654 (.A(net2655),
    .X(net2654));
 sg13g2_buf_8 fanout2655 (.A(\net.in[83] ),
    .X(net2655));
 sg13g2_buf_8 fanout2656 (.A(net2658),
    .X(net2656));
 sg13g2_buf_8 fanout2657 (.A(net2658),
    .X(net2657));
 sg13g2_buf_8 fanout2658 (.A(\net.in[82] ),
    .X(net2658));
 sg13g2_buf_4 fanout2659 (.X(net2659),
    .A(net2660));
 sg13g2_buf_16 fanout2660 (.X(net2660),
    .A(\net.in[79] ));
 sg13g2_buf_4 fanout2661 (.X(net2661),
    .A(net2665));
 sg13g2_buf_8 fanout2662 (.A(net2665),
    .X(net2662));
 sg13g2_buf_8 fanout2663 (.A(net2665),
    .X(net2663));
 sg13g2_buf_8 fanout2664 (.A(net2665),
    .X(net2664));
 sg13g2_buf_8 fanout2665 (.A(\net.in[78] ),
    .X(net2665));
 sg13g2_buf_8 fanout2666 (.A(net2667),
    .X(net2666));
 sg13g2_buf_8 fanout2667 (.A(net352),
    .X(net2667));
 sg13g2_buf_8 fanout2668 (.A(net2671),
    .X(net2668));
 sg13g2_buf_4 fanout2669 (.X(net2669),
    .A(net2671));
 sg13g2_buf_8 fanout2670 (.A(net2671),
    .X(net2670));
 sg13g2_buf_8 fanout2671 (.A(\net.in[76] ),
    .X(net2671));
 sg13g2_buf_8 fanout2672 (.A(\net.in[75] ),
    .X(net2672));
 sg13g2_buf_8 fanout2673 (.A(\net.in[75] ),
    .X(net2673));
 sg13g2_buf_8 fanout2674 (.A(net2675),
    .X(net2674));
 sg13g2_buf_8 fanout2675 (.A(net383),
    .X(net2675));
 sg13g2_buf_8 fanout2676 (.A(\net.in[74] ),
    .X(net2676));
 sg13g2_buf_8 fanout2677 (.A(net2681),
    .X(net2677));
 sg13g2_buf_8 fanout2678 (.A(net2680),
    .X(net2678));
 sg13g2_buf_8 fanout2679 (.A(net2680),
    .X(net2679));
 sg13g2_buf_8 fanout2680 (.A(net2681),
    .X(net2680));
 sg13g2_buf_8 fanout2681 (.A(\net.in[73] ),
    .X(net2681));
 sg13g2_buf_8 fanout2682 (.A(net2685),
    .X(net2682));
 sg13g2_buf_8 fanout2683 (.A(net2685),
    .X(net2683));
 sg13g2_buf_2 fanout2684 (.A(net2685),
    .X(net2684));
 sg13g2_buf_8 fanout2685 (.A(\net.in[72] ),
    .X(net2685));
 sg13g2_buf_8 fanout2686 (.A(net2689),
    .X(net2686));
 sg13g2_buf_16 fanout2687 (.X(net2687),
    .A(net2689));
 sg13g2_buf_8 fanout2688 (.A(net2689),
    .X(net2688));
 sg13g2_buf_8 fanout2689 (.A(\net.in[71] ),
    .X(net2689));
 sg13g2_buf_4 fanout2690 (.X(net2690),
    .A(net2691));
 sg13g2_buf_8 fanout2691 (.A(\net.in[70] ),
    .X(net2691));
 sg13g2_buf_8 fanout2692 (.A(\net.in[70] ),
    .X(net2692));
 sg13g2_buf_4 fanout2693 (.X(net2693),
    .A(\net.in[70] ));
 sg13g2_buf_8 fanout2694 (.A(net2696),
    .X(net2694));
 sg13g2_buf_2 fanout2695 (.A(net2696),
    .X(net2695));
 sg13g2_buf_8 fanout2696 (.A(net2697),
    .X(net2696));
 sg13g2_buf_8 fanout2697 (.A(\net.in[69] ),
    .X(net2697));
 sg13g2_buf_8 fanout2698 (.A(net2699),
    .X(net2698));
 sg13g2_buf_16 fanout2699 (.X(net2699),
    .A(net369));
 sg13g2_buf_8 fanout2700 (.A(net338),
    .X(net2700));
 sg13g2_buf_4 fanout2701 (.X(net2701),
    .A(net338));
 sg13g2_buf_8 fanout2702 (.A(net363),
    .X(net2702));
 sg13g2_buf_4 fanout2703 (.X(net2703),
    .A(\net.in[66] ));
 sg13g2_buf_8 fanout2704 (.A(\net.in[65] ),
    .X(net2704));
 sg13g2_buf_16 fanout2705 (.X(net2705),
    .A(net345));
 sg13g2_buf_4 fanout2706 (.X(net2706),
    .A(\net.in[63] ));
 sg13g2_buf_16 fanout2707 (.X(net2707),
    .A(\net.in[62] ));
 sg13g2_buf_8 fanout2708 (.A(\net.in[62] ),
    .X(net2708));
 sg13g2_buf_4 fanout2709 (.X(net2709),
    .A(net2710));
 sg13g2_buf_16 fanout2710 (.X(net2710),
    .A(net382));
 sg13g2_buf_8 fanout2711 (.A(net2713),
    .X(net2711));
 sg13g2_buf_8 fanout2712 (.A(net2713),
    .X(net2712));
 sg13g2_buf_8 fanout2713 (.A(\net.in[60] ),
    .X(net2713));
 sg13g2_buf_8 fanout2714 (.A(net2715),
    .X(net2714));
 sg13g2_buf_8 fanout2715 (.A(\net.in[59] ),
    .X(net2715));
 sg13g2_buf_8 fanout2716 (.A(net2717),
    .X(net2716));
 sg13g2_buf_8 fanout2717 (.A(net2719),
    .X(net2717));
 sg13g2_buf_8 fanout2718 (.A(net2719),
    .X(net2718));
 sg13g2_buf_8 fanout2719 (.A(\net.in[58] ),
    .X(net2719));
 sg13g2_buf_4 fanout2720 (.X(net2720),
    .A(net2721));
 sg13g2_buf_8 fanout2721 (.A(net2724),
    .X(net2721));
 sg13g2_buf_8 fanout2722 (.A(net2724),
    .X(net2722));
 sg13g2_buf_8 fanout2723 (.A(net2724),
    .X(net2723));
 sg13g2_buf_8 fanout2724 (.A(net371),
    .X(net2724));
 sg13g2_buf_8 fanout2725 (.A(net2727),
    .X(net2725));
 sg13g2_buf_4 fanout2726 (.X(net2726),
    .A(net2727));
 sg13g2_buf_8 fanout2727 (.A(\net.in[56] ),
    .X(net2727));
 sg13g2_buf_8 fanout2728 (.A(net2730),
    .X(net2728));
 sg13g2_buf_8 fanout2729 (.A(net2730),
    .X(net2729));
 sg13g2_buf_8 fanout2730 (.A(\net.in[55] ),
    .X(net2730));
 sg13g2_buf_8 fanout2731 (.A(net2732),
    .X(net2731));
 sg13g2_buf_8 fanout2732 (.A(\net.in[54] ),
    .X(net2732));
 sg13g2_buf_16 fanout2733 (.X(net2733),
    .A(\net.in[54] ));
 sg13g2_buf_8 fanout2734 (.A(net2737),
    .X(net2734));
 sg13g2_buf_8 fanout2735 (.A(net2736),
    .X(net2735));
 sg13g2_buf_8 fanout2736 (.A(net2737),
    .X(net2736));
 sg13g2_buf_4 fanout2737 (.X(net2737),
    .A(\net.in[53] ));
 sg13g2_buf_8 fanout2738 (.A(\net.in[52] ),
    .X(net2738));
 sg13g2_buf_8 fanout2739 (.A(\net.in[52] ),
    .X(net2739));
 sg13g2_buf_8 fanout2740 (.A(net2742),
    .X(net2740));
 sg13g2_buf_8 fanout2741 (.A(net2742),
    .X(net2741));
 sg13g2_buf_4 fanout2742 (.X(net2742),
    .A(net325));
 sg13g2_buf_8 fanout2743 (.A(\net.in[50] ),
    .X(net2743));
 sg13g2_buf_4 fanout2744 (.X(net2744),
    .A(\net.in[50] ));
 sg13g2_buf_8 fanout2745 (.A(net302),
    .X(net2745));
 sg13g2_buf_8 fanout2746 (.A(net2747),
    .X(net2746));
 sg13g2_buf_8 fanout2747 (.A(\net.in[46] ),
    .X(net2747));
 sg13g2_buf_8 fanout2748 (.A(\net.in[45] ),
    .X(net2748));
 sg13g2_buf_4 fanout2749 (.X(net2749),
    .A(\net.in[45] ));
 sg13g2_buf_8 fanout2750 (.A(net2751),
    .X(net2750));
 sg13g2_buf_8 fanout2751 (.A(\net.in[44] ),
    .X(net2751));
 sg13g2_buf_8 fanout2752 (.A(net2753),
    .X(net2752));
 sg13g2_buf_8 fanout2753 (.A(net384),
    .X(net2753));
 sg13g2_buf_8 fanout2754 (.A(\net.in[42] ),
    .X(net2754));
 sg13g2_buf_8 fanout2755 (.A(net361),
    .X(net2755));
 sg13g2_buf_8 fanout2756 (.A(net2757),
    .X(net2756));
 sg13g2_buf_8 fanout2757 (.A(net2759),
    .X(net2757));
 sg13g2_buf_8 fanout2758 (.A(net2759),
    .X(net2758));
 sg13g2_buf_8 fanout2759 (.A(\net.in[41] ),
    .X(net2759));
 sg13g2_buf_8 fanout2760 (.A(\net.in[40] ),
    .X(net2760));
 sg13g2_buf_8 fanout2761 (.A(\net.in[40] ),
    .X(net2761));
 sg13g2_buf_8 fanout2762 (.A(net2763),
    .X(net2762));
 sg13g2_buf_8 fanout2763 (.A(\net.in[39] ),
    .X(net2763));
 sg13g2_buf_8 fanout2764 (.A(net2765),
    .X(net2764));
 sg13g2_buf_8 fanout2765 (.A(net315),
    .X(net2765));
 sg13g2_buf_8 fanout2766 (.A(net2768),
    .X(net2766));
 sg13g2_buf_8 fanout2767 (.A(net2768),
    .X(net2767));
 sg13g2_buf_8 fanout2768 (.A(\net.in[37] ),
    .X(net2768));
 sg13g2_buf_8 fanout2769 (.A(net2770),
    .X(net2769));
 sg13g2_buf_8 fanout2770 (.A(\net.in[36] ),
    .X(net2770));
 sg13g2_buf_4 fanout2771 (.X(net2771),
    .A(\net.in[36] ));
 sg13g2_buf_16 fanout2772 (.X(net2772),
    .A(\net.in[35] ));
 sg13g2_buf_16 fanout2773 (.X(net2773),
    .A(\net.in[34] ));
 sg13g2_buf_8 fanout2774 (.A(\net.in[30] ),
    .X(net2774));
 sg13g2_buf_2 fanout2775 (.A(net335),
    .X(net2775));
 sg13g2_buf_8 fanout2776 (.A(net2777),
    .X(net2776));
 sg13g2_buf_8 fanout2777 (.A(\net.in[29] ),
    .X(net2777));
 sg13g2_buf_8 fanout2778 (.A(net2780),
    .X(net2778));
 sg13g2_buf_4 fanout2779 (.X(net2779),
    .A(net2780));
 sg13g2_buf_8 fanout2780 (.A(\net.in[28] ),
    .X(net2780));
 sg13g2_buf_8 fanout2781 (.A(net2782),
    .X(net2781));
 sg13g2_buf_16 fanout2782 (.X(net2782),
    .A(net359));
 sg13g2_buf_4 fanout2783 (.X(net2783),
    .A(net359));
 sg13g2_buf_8 fanout2784 (.A(\net.in[26] ),
    .X(net2784));
 sg13g2_buf_4 fanout2785 (.X(net2785),
    .A(net2786));
 sg13g2_buf_16 fanout2786 (.X(net2786),
    .A(\net.in[26] ));
 sg13g2_buf_8 fanout2787 (.A(net2789),
    .X(net2787));
 sg13g2_buf_8 fanout2788 (.A(net2789),
    .X(net2788));
 sg13g2_buf_16 fanout2789 (.X(net2789),
    .A(\net.in[25] ));
 sg13g2_buf_8 fanout2790 (.A(net2791),
    .X(net2790));
 sg13g2_buf_16 fanout2791 (.X(net2791),
    .A(\net.in[24] ));
 sg13g2_buf_8 fanout2792 (.A(net2794),
    .X(net2792));
 sg13g2_buf_4 fanout2793 (.X(net2793),
    .A(net2794));
 sg13g2_buf_16 fanout2794 (.X(net2794),
    .A(\net.in[23] ));
 sg13g2_buf_8 fanout2795 (.A(net2796),
    .X(net2795));
 sg13g2_buf_16 fanout2796 (.X(net2796),
    .A(\net.in[22] ));
 sg13g2_buf_8 fanout2797 (.A(\net.in[21] ),
    .X(net2797));
 sg13g2_buf_4 fanout2798 (.X(net2798),
    .A(\net.in[21] ));
 sg13g2_buf_8 fanout2799 (.A(\net.in[21] ),
    .X(net2799));
 sg13g2_buf_8 fanout2800 (.A(net2801),
    .X(net2800));
 sg13g2_buf_8 fanout2801 (.A(net297),
    .X(net2801));
 sg13g2_buf_8 fanout2802 (.A(net346),
    .X(net2802));
 sg13g2_buf_8 fanout2803 (.A(\calc_categories[6].sum_bits.popcount128.ad0.genblk1[108].add3.a ),
    .X(net2803));
 sg13g2_buf_2 fanout2804 (.A(net332),
    .X(net2804));
 sg13g2_buf_8 fanout2805 (.A(net2806),
    .X(net2805));
 sg13g2_buf_16 fanout2806 (.X(net2806),
    .A(\net.in[11] ));
 sg13g2_buf_16 fanout2807 (.X(net2807),
    .A(\net.in[9] ));
 sg13g2_buf_16 fanout2808 (.X(net2808),
    .A(\net.in[9] ));
 sg13g2_buf_8 fanout2809 (.A(net2811),
    .X(net2809));
 sg13g2_buf_8 fanout2810 (.A(net2811),
    .X(net2810));
 sg13g2_buf_8 fanout2811 (.A(net298),
    .X(net2811));
 sg13g2_buf_8 fanout2812 (.A(\net.in[7] ),
    .X(net2812));
 sg13g2_buf_4 fanout2813 (.X(net2813),
    .A(\net.in[7] ));
 sg13g2_buf_16 fanout2814 (.X(net2814),
    .A(net2815));
 sg13g2_buf_16 fanout2815 (.X(net2815),
    .A(\net.in[6] ));
 sg13g2_buf_8 fanout2816 (.A(net2817),
    .X(net2816));
 sg13g2_buf_16 fanout2817 (.X(net2817),
    .A(\net.in[5] ));
 sg13g2_buf_4 fanout2818 (.X(net2818),
    .A(net2820));
 sg13g2_buf_2 fanout2819 (.A(net2820),
    .X(net2819));
 sg13g2_buf_4 fanout2820 (.X(net2820),
    .A(net2821));
 sg13g2_buf_2 fanout2821 (.A(net2822),
    .X(net2821));
 sg13g2_buf_2 fanout2822 (.A(net2823),
    .X(net2822));
 sg13g2_buf_4 fanout2823 (.X(net2823),
    .A(net2850));
 sg13g2_buf_4 fanout2824 (.X(net2824),
    .A(net2837));
 sg13g2_buf_4 fanout2825 (.X(net2825),
    .A(net2837));
 sg13g2_buf_2 fanout2826 (.A(net2828),
    .X(net2826));
 sg13g2_buf_2 fanout2827 (.A(net2828),
    .X(net2827));
 sg13g2_buf_2 fanout2828 (.A(net2829),
    .X(net2828));
 sg13g2_buf_4 fanout2829 (.X(net2829),
    .A(net2837));
 sg13g2_buf_2 fanout2830 (.A(net2832),
    .X(net2830));
 sg13g2_buf_1 fanout2831 (.A(net2832),
    .X(net2831));
 sg13g2_buf_2 fanout2832 (.A(net2836),
    .X(net2832));
 sg13g2_buf_2 fanout2833 (.A(net2836),
    .X(net2833));
 sg13g2_buf_4 fanout2834 (.X(net2834),
    .A(net2835));
 sg13g2_buf_4 fanout2835 (.X(net2835),
    .A(net2836));
 sg13g2_buf_4 fanout2836 (.X(net2836),
    .A(net2837));
 sg13g2_buf_2 fanout2837 (.A(net2850),
    .X(net2837));
 sg13g2_buf_2 fanout2838 (.A(net2841),
    .X(net2838));
 sg13g2_buf_2 fanout2839 (.A(net2840),
    .X(net2839));
 sg13g2_buf_2 fanout2840 (.A(net2841),
    .X(net2840));
 sg13g2_buf_2 fanout2841 (.A(net2843),
    .X(net2841));
 sg13g2_buf_4 fanout2842 (.X(net2842),
    .A(net2843));
 sg13g2_buf_2 fanout2843 (.A(net2847),
    .X(net2843));
 sg13g2_buf_2 fanout2844 (.A(net2845),
    .X(net2844));
 sg13g2_buf_2 fanout2845 (.A(net2846),
    .X(net2845));
 sg13g2_buf_4 fanout2846 (.X(net2846),
    .A(net2847));
 sg13g2_buf_2 fanout2847 (.A(net2850),
    .X(net2847));
 sg13g2_buf_2 fanout2848 (.A(net2850),
    .X(net2848));
 sg13g2_buf_2 fanout2849 (.A(net2850),
    .X(net2849));
 sg13g2_buf_8 fanout2850 (.A(net2888),
    .X(net2850));
 sg13g2_buf_4 fanout2851 (.X(net2851),
    .A(net2852));
 sg13g2_buf_4 fanout2852 (.X(net2852),
    .A(net2853));
 sg13g2_buf_4 fanout2853 (.X(net2853),
    .A(net2880));
 sg13g2_buf_4 fanout2854 (.X(net2854),
    .A(net2856));
 sg13g2_buf_4 fanout2855 (.X(net2855),
    .A(net2856));
 sg13g2_buf_2 fanout2856 (.A(net2869),
    .X(net2856));
 sg13g2_buf_2 fanout2857 (.A(net2858),
    .X(net2857));
 sg13g2_buf_4 fanout2858 (.X(net2858),
    .A(net2861));
 sg13g2_buf_2 fanout2859 (.A(net2860),
    .X(net2859));
 sg13g2_buf_4 fanout2860 (.X(net2860),
    .A(net2861));
 sg13g2_buf_2 fanout2861 (.A(net2869),
    .X(net2861));
 sg13g2_buf_4 fanout2862 (.X(net2862),
    .A(net2864));
 sg13g2_buf_4 fanout2863 (.X(net2863),
    .A(net2864));
 sg13g2_buf_2 fanout2864 (.A(net2869),
    .X(net2864));
 sg13g2_buf_4 fanout2865 (.X(net2865),
    .A(net2868));
 sg13g2_buf_4 fanout2866 (.X(net2866),
    .A(net2867));
 sg13g2_buf_4 fanout2867 (.X(net2867),
    .A(net2868));
 sg13g2_buf_2 fanout2868 (.A(net2869),
    .X(net2868));
 sg13g2_buf_2 fanout2869 (.A(net2880),
    .X(net2869));
 sg13g2_buf_4 fanout2870 (.X(net2870),
    .A(net2871));
 sg13g2_buf_4 fanout2871 (.X(net2871),
    .A(net2872));
 sg13g2_buf_2 fanout2872 (.A(net2873),
    .X(net2872));
 sg13g2_buf_4 fanout2873 (.X(net2873),
    .A(net2880));
 sg13g2_buf_2 fanout2874 (.A(net2875),
    .X(net2874));
 sg13g2_buf_2 fanout2875 (.A(net2876),
    .X(net2875));
 sg13g2_buf_4 fanout2876 (.X(net2876),
    .A(net2879));
 sg13g2_buf_4 fanout2877 (.X(net2877),
    .A(net2878));
 sg13g2_buf_2 fanout2878 (.A(net2879),
    .X(net2878));
 sg13g2_buf_2 fanout2879 (.A(net2880),
    .X(net2879));
 sg13g2_buf_4 fanout2880 (.X(net2880),
    .A(net2888));
 sg13g2_buf_2 fanout2881 (.A(net2882),
    .X(net2881));
 sg13g2_buf_2 fanout2882 (.A(net2886),
    .X(net2882));
 sg13g2_buf_4 fanout2883 (.X(net2883),
    .A(net2886));
 sg13g2_buf_2 fanout2884 (.A(net2885),
    .X(net2884));
 sg13g2_buf_4 fanout2885 (.X(net2885),
    .A(net2886));
 sg13g2_buf_2 fanout2886 (.A(net2887),
    .X(net2886));
 sg13g2_buf_8 fanout2887 (.A(net2888),
    .X(net2887));
 sg13g2_buf_8 fanout2888 (.A(uio_in[7]),
    .X(net2888));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_16 wire9 (.X(net9),
    .A(_07681_));
 sg13g2_tielo tt_um_rejunity_lgn_mnist_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sg13g2_buf_2 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sg13g2_buf_2 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2__leaf_clk));
 sg13g2_buf_2 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3__leaf_clk));
 sg13g2_buf_2 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4__leaf_clk));
 sg13g2_buf_2 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5__leaf_clk));
 sg13g2_buf_2 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6__leaf_clk));
 sg13g2_buf_2 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7__leaf_clk));
 sg13g2_buf_2 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8__leaf_clk));
 sg13g2_buf_2 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9__leaf_clk));
 sg13g2_buf_2 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10__leaf_clk));
 sg13g2_buf_2 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11__leaf_clk));
 sg13g2_buf_2 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12__leaf_clk));
 sg13g2_buf_2 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13__leaf_clk));
 sg13g2_buf_2 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14__leaf_clk));
 sg13g2_buf_2 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_3__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_4__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_6__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_11__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_12__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_15__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_77_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_78_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_71_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_76_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_68_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_73_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_74_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_67_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_14_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_59_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_62_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_63_clk));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_48_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_51_clk));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_46_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload38 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload39 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_61_clk));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload42 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload43 (.A(clknet_leaf_39_clk));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_40_clk));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_60_clk));
 sg13g2_inv_2 clkload46 (.A(clknet_leaf_32_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\net.in[16] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00049_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold3 (.A(\net.in[48] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00073_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold5 (.A(\net.in[128] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold6 (.A(\net.in[160] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold7 (.A(\net.in[2] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold8 (.A(\net.in[18] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold9 (.A(\net.in[240] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold10 (.A(\net.in[32] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold11 (.A(\net.in[239] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold12 (.A(\net.in[144] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold13 (.A(\net.in[248] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold14 (.A(\net.in[15] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold15 (.A(_00040_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold16 (.A(\net.in[224] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold17 (.A(_00257_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold18 (.A(\net.in[14] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold19 (.A(\net.in[64] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold20 (.A(\net.in[0] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold21 (.A(\net.in[33] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold22 (.A(\net.in[1] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold23 (.A(\net.in[17] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold24 (.A(\net.in[216] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold25 (.A(\net.in[20] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold26 (.A(\net.in[8] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold27 (.A(\net.in[3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold28 (.A(\net.in[253] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold29 (.A(\net.in[238] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold30 (.A(\net.in[47] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold31 (.A(_00072_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold32 (.A(\net.in[81] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold33 (.A(\net.in[189] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold34 (.A(\net.in[201] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold35 (.A(_00226_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold36 (.A(\net.in[131] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold37 (.A(\net.in[200] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold38 (.A(_00225_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold39 (.A(\net.in[214] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold40 (.A(_00247_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold41 (.A(\net.in[176] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold42 (.A(\net.in[157] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold43 (.A(\net.in[38] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold44 (.A(\net.in[138] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00171_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold46 (.A(\calc_categories[0].sum_bits.popcount128.ad0.genblk1[105].add3.a ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold47 (.A(\net.in[193] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold48 (.A(\net.in[98] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold49 (.A(\net.in[96] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold50 (.A(\net.in[174] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold51 (.A(\net.in[114] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold52 (.A(\net.in[208] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold53 (.A(\net.in[51] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold54 (.A(\net.in[125] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold55 (.A(_00158_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold56 (.A(\net.in[158] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold57 (.A(\net.in[192] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold58 (.A(\net.in[31] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold59 (.A(\net.in[145] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold60 (.A(\calc_categories[6].sum_bits.popcount128.ad0.genblk1[108].add3.a ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold61 (.A(\net.in[195] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00220_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold63 (.A(\net.in[30] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold64 (.A(\net.in[94] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold65 (.A(\net.in[55] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold66 (.A(\net.in[67] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold67 (.A(\net.in[190] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold68 (.A(\net.in[171] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold69 (.A(_00204_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold70 (.A(\net.in[243] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold71 (.A(\net.in[127] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold72 (.A(\net.in[207] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold73 (.A(\net.in[63] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold74 (.A(\net.in[19] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold75 (.A(\net.in[233] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold76 (.A(\net.in[221] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold77 (.A(\net.in[250] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold78 (.A(\net.in[93] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold79 (.A(\net.in[163] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold80 (.A(\net.in[77] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold81 (.A(\net.in[222] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold82 (.A(\net.in[187] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold83 (.A(\net.in[134] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold84 (.A(\net.in[90] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold85 (.A(\net.in[204] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold86 (.A(\net.in[225] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold87 (.A(\net.in[27] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold88 (.A(\net.in[162] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold89 (.A(\net.in[42] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold90 (.A(\net.in[100] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold91 (.A(\net.in[66] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold92 (.A(\net.in[111] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold93 (.A(\net.in[173] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold94 (.A(\net.in[183] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold95 (.A(\net.in[215] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold96 (.A(\net.in[97] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold97 (.A(\net.in[68] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold98 (.A(\net.in[226] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold99 (.A(\net.in[57] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold100 (.A(\net.in[178] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold101 (.A(\net.in[135] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold102 (.A(\net.in[206] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold103 (.A(\net.in[92] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold104 (.A(\net.in[210] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold105 (.A(\net.in[155] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold106 (.A(\net.in[236] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold107 (.A(\net.in[159] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold108 (.A(\net.in[13] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold109 (.A(\net.in[112] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold110 (.A(\net.in[61] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold111 (.A(\net.in[74] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold112 (.A(\net.in[43] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold113 (.A(\net.in[219] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold114 (.A(_00252_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold115 (.A(\net.in[121] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold116 (.A(\net.in[202] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold117 (.A(\calc_categories[0].sum_bits.popcount128.ad0.genblk1[105].add3.a ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold118 (.A(\net.in[111] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold119 (.A(\net.in[114] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold120 (.A(\net.in[226] ),
    .X(net392));
 sg13g2_antennanp ANTENNA_1 (.A(_00472_));
 sg13g2_antennanp ANTENNA_2 (.A(_00472_));
 sg13g2_antennanp ANTENNA_3 (.A(_05176_));
 sg13g2_antennanp ANTENNA_4 (.A(_05176_));
 sg13g2_antennanp ANTENNA_5 (.A(_05176_));
 sg13g2_antennanp ANTENNA_6 (.A(_05176_));
 sg13g2_antennanp ANTENNA_7 (.A(_05176_));
 sg13g2_antennanp ANTENNA_8 (.A(_05176_));
 sg13g2_antennanp ANTENNA_9 (.A(_05176_));
 sg13g2_antennanp ANTENNA_10 (.A(_05176_));
 sg13g2_antennanp ANTENNA_11 (.A(_05176_));
 sg13g2_antennanp ANTENNA_12 (.A(_05176_));
 sg13g2_antennanp ANTENNA_13 (.A(_05176_));
 sg13g2_antennanp ANTENNA_14 (.A(_05561_));
 sg13g2_antennanp ANTENNA_15 (.A(_05561_));
 sg13g2_antennanp ANTENNA_16 (.A(_05561_));
 sg13g2_antennanp ANTENNA_17 (.A(_05561_));
 sg13g2_antennanp ANTENNA_18 (.A(_05561_));
 sg13g2_antennanp ANTENNA_19 (.A(_05561_));
 sg13g2_antennanp ANTENNA_20 (.A(_05561_));
 sg13g2_antennanp ANTENNA_21 (.A(_05561_));
 sg13g2_antennanp ANTENNA_22 (.A(_05561_));
 sg13g2_antennanp ANTENNA_23 (.A(_05561_));
 sg13g2_antennanp ANTENNA_24 (.A(_05561_));
 sg13g2_antennanp ANTENNA_25 (.A(_05561_));
 sg13g2_antennanp ANTENNA_26 (.A(_05561_));
 sg13g2_antennanp ANTENNA_27 (.A(_05561_));
 sg13g2_antennanp ANTENNA_28 (.A(_05561_));
 sg13g2_antennanp ANTENNA_29 (.A(_05561_));
 sg13g2_antennanp ANTENNA_30 (.A(_05847_));
 sg13g2_antennanp ANTENNA_31 (.A(_05847_));
 sg13g2_antennanp ANTENNA_32 (.A(_05847_));
 sg13g2_antennanp ANTENNA_33 (.A(_05847_));
 sg13g2_antennanp ANTENNA_34 (.A(_05847_));
 sg13g2_antennanp ANTENNA_35 (.A(_05847_));
 sg13g2_antennanp ANTENNA_36 (.A(_05847_));
 sg13g2_antennanp ANTENNA_37 (.A(_05847_));
 sg13g2_antennanp ANTENNA_38 (.A(_05847_));
 sg13g2_antennanp ANTENNA_39 (.A(_05847_));
 sg13g2_antennanp ANTENNA_40 (.A(_05847_));
 sg13g2_antennanp ANTENNA_41 (.A(_05847_));
 sg13g2_antennanp ANTENNA_42 (.A(_05847_));
 sg13g2_antennanp ANTENNA_43 (.A(_05847_));
 sg13g2_antennanp ANTENNA_44 (.A(_05847_));
 sg13g2_antennanp ANTENNA_45 (.A(_05847_));
 sg13g2_antennanp ANTENNA_46 (.A(_05858_));
 sg13g2_antennanp ANTENNA_47 (.A(_05858_));
 sg13g2_antennanp ANTENNA_48 (.A(_05858_));
 sg13g2_antennanp ANTENNA_49 (.A(_07984_));
 sg13g2_antennanp ANTENNA_50 (.A(_07984_));
 sg13g2_antennanp ANTENNA_51 (.A(_07984_));
 sg13g2_antennanp ANTENNA_52 (.A(_07984_));
 sg13g2_antennanp ANTENNA_53 (.A(_07984_));
 sg13g2_antennanp ANTENNA_54 (.A(_07984_));
 sg13g2_antennanp ANTENNA_55 (.A(_08349_));
 sg13g2_antennanp ANTENNA_56 (.A(_08349_));
 sg13g2_antennanp ANTENNA_57 (.A(clk));
 sg13g2_antennanp ANTENNA_58 (.A(clk));
 sg13g2_antennanp ANTENNA_59 (.A(\net.in[112] ));
 sg13g2_antennanp ANTENNA_60 (.A(\net.in[112] ));
 sg13g2_antennanp ANTENNA_61 (.A(\net.in[112] ));
 sg13g2_antennanp ANTENNA_62 (.A(\net.in[112] ));
 sg13g2_antennanp ANTENNA_63 (.A(\net.in[112] ));
 sg13g2_antennanp ANTENNA_64 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_65 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_66 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_67 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_68 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_69 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_70 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_71 (.A(\net.in[209] ));
 sg13g2_antennanp ANTENNA_72 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_73 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_74 (.A(net2199));
 sg13g2_antennanp ANTENNA_75 (.A(net2199));
 sg13g2_antennanp ANTENNA_76 (.A(net2199));
 sg13g2_antennanp ANTENNA_77 (.A(net2199));
 sg13g2_antennanp ANTENNA_78 (.A(net2199));
 sg13g2_antennanp ANTENNA_79 (.A(net2199));
 sg13g2_antennanp ANTENNA_80 (.A(net2199));
 sg13g2_antennanp ANTENNA_81 (.A(net2199));
 sg13g2_antennanp ANTENNA_82 (.A(net2199));
 sg13g2_antennanp ANTENNA_83 (.A(net2199));
 sg13g2_antennanp ANTENNA_84 (.A(net2199));
 sg13g2_antennanp ANTENNA_85 (.A(net2199));
 sg13g2_antennanp ANTENNA_86 (.A(net2199));
 sg13g2_antennanp ANTENNA_87 (.A(net2199));
 sg13g2_antennanp ANTENNA_88 (.A(net2199));
 sg13g2_antennanp ANTENNA_89 (.A(net2199));
 sg13g2_antennanp ANTENNA_90 (.A(net2221));
 sg13g2_antennanp ANTENNA_91 (.A(net2221));
 sg13g2_antennanp ANTENNA_92 (.A(net2221));
 sg13g2_antennanp ANTENNA_93 (.A(net2221));
 sg13g2_antennanp ANTENNA_94 (.A(net2221));
 sg13g2_antennanp ANTENNA_95 (.A(net2221));
 sg13g2_antennanp ANTENNA_96 (.A(net2221));
 sg13g2_antennanp ANTENNA_97 (.A(net2221));
 sg13g2_antennanp ANTENNA_98 (.A(net2221));
 sg13g2_antennanp ANTENNA_99 (.A(net2221));
 sg13g2_antennanp ANTENNA_100 (.A(net2221));
 sg13g2_antennanp ANTENNA_101 (.A(net2221));
 sg13g2_antennanp ANTENNA_102 (.A(net2221));
 sg13g2_antennanp ANTENNA_103 (.A(net2221));
 sg13g2_antennanp ANTENNA_104 (.A(net2221));
 sg13g2_antennanp ANTENNA_105 (.A(net2221));
 sg13g2_antennanp ANTENNA_106 (.A(net2238));
 sg13g2_antennanp ANTENNA_107 (.A(net2238));
 sg13g2_antennanp ANTENNA_108 (.A(net2238));
 sg13g2_antennanp ANTENNA_109 (.A(net2238));
 sg13g2_antennanp ANTENNA_110 (.A(net2238));
 sg13g2_antennanp ANTENNA_111 (.A(net2266));
 sg13g2_antennanp ANTENNA_112 (.A(net2266));
 sg13g2_antennanp ANTENNA_113 (.A(net2266));
 sg13g2_antennanp ANTENNA_114 (.A(net2266));
 sg13g2_antennanp ANTENNA_115 (.A(net2266));
 sg13g2_antennanp ANTENNA_116 (.A(net2266));
 sg13g2_antennanp ANTENNA_117 (.A(net2266));
 sg13g2_antennanp ANTENNA_118 (.A(net2266));
 sg13g2_antennanp ANTENNA_119 (.A(net2266));
 sg13g2_antennanp ANTENNA_120 (.A(net2266));
 sg13g2_antennanp ANTENNA_121 (.A(net2266));
 sg13g2_antennanp ANTENNA_122 (.A(net2266));
 sg13g2_antennanp ANTENNA_123 (.A(net2277));
 sg13g2_antennanp ANTENNA_124 (.A(net2277));
 sg13g2_antennanp ANTENNA_125 (.A(net2277));
 sg13g2_antennanp ANTENNA_126 (.A(net2277));
 sg13g2_antennanp ANTENNA_127 (.A(net2277));
 sg13g2_antennanp ANTENNA_128 (.A(net2277));
 sg13g2_antennanp ANTENNA_129 (.A(net2277));
 sg13g2_antennanp ANTENNA_130 (.A(net2277));
 sg13g2_antennanp ANTENNA_131 (.A(net2277));
 sg13g2_antennanp ANTENNA_132 (.A(net2277));
 sg13g2_antennanp ANTENNA_133 (.A(net2277));
 sg13g2_antennanp ANTENNA_134 (.A(net2277));
 sg13g2_antennanp ANTENNA_135 (.A(net2277));
 sg13g2_antennanp ANTENNA_136 (.A(net2277));
 sg13g2_antennanp ANTENNA_137 (.A(net2277));
 sg13g2_antennanp ANTENNA_138 (.A(net2277));
 sg13g2_antennanp ANTENNA_139 (.A(net2277));
 sg13g2_antennanp ANTENNA_140 (.A(net2277));
 sg13g2_antennanp ANTENNA_141 (.A(net2277));
 sg13g2_antennanp ANTENNA_142 (.A(net2277));
 sg13g2_antennanp ANTENNA_143 (.A(net2281));
 sg13g2_antennanp ANTENNA_144 (.A(net2281));
 sg13g2_antennanp ANTENNA_145 (.A(net2281));
 sg13g2_antennanp ANTENNA_146 (.A(net2281));
 sg13g2_antennanp ANTENNA_147 (.A(net2281));
 sg13g2_antennanp ANTENNA_148 (.A(net2281));
 sg13g2_antennanp ANTENNA_149 (.A(net2281));
 sg13g2_antennanp ANTENNA_150 (.A(net2281));
 sg13g2_antennanp ANTENNA_151 (.A(net2281));
 sg13g2_antennanp ANTENNA_152 (.A(net2281));
 sg13g2_antennanp ANTENNA_153 (.A(net2281));
 sg13g2_antennanp ANTENNA_154 (.A(net2281));
 sg13g2_antennanp ANTENNA_155 (.A(net2281));
 sg13g2_antennanp ANTENNA_156 (.A(net2281));
 sg13g2_antennanp ANTENNA_157 (.A(net2284));
 sg13g2_antennanp ANTENNA_158 (.A(net2284));
 sg13g2_antennanp ANTENNA_159 (.A(net2284));
 sg13g2_antennanp ANTENNA_160 (.A(net2284));
 sg13g2_antennanp ANTENNA_161 (.A(net2284));
 sg13g2_antennanp ANTENNA_162 (.A(net2403));
 sg13g2_antennanp ANTENNA_163 (.A(net2403));
 sg13g2_antennanp ANTENNA_164 (.A(net2403));
 sg13g2_antennanp ANTENNA_165 (.A(net2403));
 sg13g2_antennanp ANTENNA_166 (.A(net2403));
 sg13g2_antennanp ANTENNA_167 (.A(net2403));
 sg13g2_antennanp ANTENNA_168 (.A(net2403));
 sg13g2_antennanp ANTENNA_169 (.A(net2403));
 sg13g2_antennanp ANTENNA_170 (.A(net2403));
 sg13g2_antennanp ANTENNA_171 (.A(net2403));
 sg13g2_antennanp ANTENNA_172 (.A(net2403));
 sg13g2_antennanp ANTENNA_173 (.A(net2403));
 sg13g2_antennanp ANTENNA_174 (.A(net2403));
 sg13g2_antennanp ANTENNA_175 (.A(net2403));
 sg13g2_antennanp ANTENNA_176 (.A(net2403));
 sg13g2_antennanp ANTENNA_177 (.A(net2403));
 sg13g2_antennanp ANTENNA_178 (.A(net2403));
 sg13g2_antennanp ANTENNA_179 (.A(net2403));
 sg13g2_antennanp ANTENNA_180 (.A(net2403));
 sg13g2_antennanp ANTENNA_181 (.A(net2403));
 sg13g2_antennanp ANTENNA_182 (.A(net2411));
 sg13g2_antennanp ANTENNA_183 (.A(net2411));
 sg13g2_antennanp ANTENNA_184 (.A(net2411));
 sg13g2_antennanp ANTENNA_185 (.A(net2411));
 sg13g2_antennanp ANTENNA_186 (.A(net2411));
 sg13g2_antennanp ANTENNA_187 (.A(net2463));
 sg13g2_antennanp ANTENNA_188 (.A(net2463));
 sg13g2_antennanp ANTENNA_189 (.A(net2463));
 sg13g2_antennanp ANTENNA_190 (.A(net2463));
 sg13g2_antennanp ANTENNA_191 (.A(net2463));
 sg13g2_antennanp ANTENNA_192 (.A(net2463));
 sg13g2_antennanp ANTENNA_193 (.A(net2463));
 sg13g2_antennanp ANTENNA_194 (.A(net2463));
 sg13g2_antennanp ANTENNA_195 (.A(net2463));
 sg13g2_antennanp ANTENNA_196 (.A(net2463));
 sg13g2_antennanp ANTENNA_197 (.A(net2463));
 sg13g2_antennanp ANTENNA_198 (.A(net2463));
 sg13g2_antennanp ANTENNA_199 (.A(net2463));
 sg13g2_antennanp ANTENNA_200 (.A(net2463));
 sg13g2_antennanp ANTENNA_201 (.A(net2465));
 sg13g2_antennanp ANTENNA_202 (.A(net2465));
 sg13g2_antennanp ANTENNA_203 (.A(net2465));
 sg13g2_antennanp ANTENNA_204 (.A(net2465));
 sg13g2_antennanp ANTENNA_205 (.A(net2497));
 sg13g2_antennanp ANTENNA_206 (.A(net2497));
 sg13g2_antennanp ANTENNA_207 (.A(net2497));
 sg13g2_antennanp ANTENNA_208 (.A(net2497));
 sg13g2_antennanp ANTENNA_209 (.A(net2497));
 sg13g2_antennanp ANTENNA_210 (.A(net2497));
 sg13g2_antennanp ANTENNA_211 (.A(net2497));
 sg13g2_antennanp ANTENNA_212 (.A(net2497));
 sg13g2_antennanp ANTENNA_213 (.A(net2497));
 sg13g2_antennanp ANTENNA_214 (.A(net2497));
 sg13g2_antennanp ANTENNA_215 (.A(net2497));
 sg13g2_antennanp ANTENNA_216 (.A(net2497));
 sg13g2_antennanp ANTENNA_217 (.A(net2497));
 sg13g2_antennanp ANTENNA_218 (.A(net2497));
 sg13g2_antennanp ANTENNA_219 (.A(net2497));
 sg13g2_antennanp ANTENNA_220 (.A(net2497));
 sg13g2_antennanp ANTENNA_221 (.A(net2497));
 sg13g2_antennanp ANTENNA_222 (.A(net2497));
 sg13g2_antennanp ANTENNA_223 (.A(net2501));
 sg13g2_antennanp ANTENNA_224 (.A(net2501));
 sg13g2_antennanp ANTENNA_225 (.A(net2501));
 sg13g2_antennanp ANTENNA_226 (.A(net2501));
 sg13g2_antennanp ANTENNA_227 (.A(net2501));
 sg13g2_antennanp ANTENNA_228 (.A(net2501));
 sg13g2_antennanp ANTENNA_229 (.A(net2501));
 sg13g2_antennanp ANTENNA_230 (.A(net2501));
 sg13g2_antennanp ANTENNA_231 (.A(net2501));
 sg13g2_antennanp ANTENNA_232 (.A(net2501));
 sg13g2_antennanp ANTENNA_233 (.A(net2501));
 sg13g2_antennanp ANTENNA_234 (.A(net2501));
 sg13g2_antennanp ANTENNA_235 (.A(net2501));
 sg13g2_antennanp ANTENNA_236 (.A(net2501));
 sg13g2_antennanp ANTENNA_237 (.A(net2501));
 sg13g2_antennanp ANTENNA_238 (.A(net2501));
 sg13g2_antennanp ANTENNA_239 (.A(net2501));
 sg13g2_antennanp ANTENNA_240 (.A(net2501));
 sg13g2_antennanp ANTENNA_241 (.A(net2501));
 sg13g2_antennanp ANTENNA_242 (.A(net2501));
 sg13g2_antennanp ANTENNA_243 (.A(net2501));
 sg13g2_antennanp ANTENNA_244 (.A(net2552));
 sg13g2_antennanp ANTENNA_245 (.A(net2552));
 sg13g2_antennanp ANTENNA_246 (.A(net2552));
 sg13g2_antennanp ANTENNA_247 (.A(net2552));
 sg13g2_antennanp ANTENNA_248 (.A(net2552));
 sg13g2_antennanp ANTENNA_249 (.A(net2552));
 sg13g2_antennanp ANTENNA_250 (.A(net2552));
 sg13g2_antennanp ANTENNA_251 (.A(net2552));
 sg13g2_antennanp ANTENNA_252 (.A(net2552));
 sg13g2_antennanp ANTENNA_253 (.A(net2552));
 sg13g2_antennanp ANTENNA_254 (.A(net2552));
 sg13g2_antennanp ANTENNA_255 (.A(net2552));
 sg13g2_antennanp ANTENNA_256 (.A(net2552));
 sg13g2_antennanp ANTENNA_257 (.A(net2552));
 sg13g2_antennanp ANTENNA_258 (.A(net2552));
 sg13g2_antennanp ANTENNA_259 (.A(net2585));
 sg13g2_antennanp ANTENNA_260 (.A(net2585));
 sg13g2_antennanp ANTENNA_261 (.A(net2585));
 sg13g2_antennanp ANTENNA_262 (.A(net2585));
 sg13g2_antennanp ANTENNA_263 (.A(net2585));
 sg13g2_antennanp ANTENNA_264 (.A(net2585));
 sg13g2_antennanp ANTENNA_265 (.A(net2585));
 sg13g2_antennanp ANTENNA_266 (.A(net2585));
 sg13g2_antennanp ANTENNA_267 (.A(net2585));
 sg13g2_antennanp ANTENNA_268 (.A(net2585));
 sg13g2_antennanp ANTENNA_269 (.A(net2651));
 sg13g2_antennanp ANTENNA_270 (.A(net2651));
 sg13g2_antennanp ANTENNA_271 (.A(net2651));
 sg13g2_antennanp ANTENNA_272 (.A(net2651));
 sg13g2_antennanp ANTENNA_273 (.A(net2651));
 sg13g2_antennanp ANTENNA_274 (.A(net2651));
 sg13g2_antennanp ANTENNA_275 (.A(net2651));
 sg13g2_antennanp ANTENNA_276 (.A(net2651));
 sg13g2_antennanp ANTENNA_277 (.A(net2651));
 sg13g2_antennanp ANTENNA_278 (.A(net2651));
 sg13g2_antennanp ANTENNA_279 (.A(net2651));
 sg13g2_antennanp ANTENNA_280 (.A(net2651));
 sg13g2_antennanp ANTENNA_281 (.A(net2651));
 sg13g2_antennanp ANTENNA_282 (.A(net2651));
 sg13g2_antennanp ANTENNA_283 (.A(net2683));
 sg13g2_antennanp ANTENNA_284 (.A(net2683));
 sg13g2_antennanp ANTENNA_285 (.A(net2683));
 sg13g2_antennanp ANTENNA_286 (.A(net2683));
 sg13g2_antennanp ANTENNA_287 (.A(net2683));
 sg13g2_antennanp ANTENNA_288 (.A(net2683));
 sg13g2_antennanp ANTENNA_289 (.A(net2683));
 sg13g2_antennanp ANTENNA_290 (.A(net2683));
 sg13g2_antennanp ANTENNA_291 (.A(net2683));
 sg13g2_antennanp ANTENNA_292 (.A(net2683));
 sg13g2_antennanp ANTENNA_293 (.A(net2683));
 sg13g2_antennanp ANTENNA_294 (.A(net2701));
 sg13g2_antennanp ANTENNA_295 (.A(net2701));
 sg13g2_antennanp ANTENNA_296 (.A(net2701));
 sg13g2_antennanp ANTENNA_297 (.A(net2701));
 sg13g2_antennanp ANTENNA_298 (.A(net2761));
 sg13g2_antennanp ANTENNA_299 (.A(net2761));
 sg13g2_antennanp ANTENNA_300 (.A(net2761));
 sg13g2_antennanp ANTENNA_301 (.A(net2761));
 sg13g2_antennanp ANTENNA_302 (.A(net2761));
 sg13g2_antennanp ANTENNA_303 (.A(net2761));
 sg13g2_antennanp ANTENNA_304 (.A(net2761));
 sg13g2_antennanp ANTENNA_305 (.A(net2761));
 sg13g2_antennanp ANTENNA_306 (.A(net2761));
 sg13g2_antennanp ANTENNA_307 (.A(net2761));
 sg13g2_antennanp ANTENNA_308 (.A(net2761));
 sg13g2_antennanp ANTENNA_309 (.A(net2761));
 sg13g2_antennanp ANTENNA_310 (.A(net2772));
 sg13g2_antennanp ANTENNA_311 (.A(net2772));
 sg13g2_antennanp ANTENNA_312 (.A(net2772));
 sg13g2_antennanp ANTENNA_313 (.A(net2772));
 sg13g2_antennanp ANTENNA_314 (.A(net2772));
 sg13g2_antennanp ANTENNA_315 (.A(net2772));
 sg13g2_antennanp ANTENNA_316 (.A(net2772));
 sg13g2_antennanp ANTENNA_317 (.A(net2772));
 sg13g2_antennanp ANTENNA_318 (.A(net2772));
 sg13g2_antennanp ANTENNA_319 (.A(net2772));
 sg13g2_antennanp ANTENNA_320 (.A(net2802));
 sg13g2_antennanp ANTENNA_321 (.A(net2802));
 sg13g2_antennanp ANTENNA_322 (.A(net2802));
 sg13g2_antennanp ANTENNA_323 (.A(net2802));
 sg13g2_antennanp ANTENNA_324 (.A(net2802));
 sg13g2_antennanp ANTENNA_325 (.A(net2802));
 sg13g2_antennanp ANTENNA_326 (.A(net2802));
 sg13g2_antennanp ANTENNA_327 (.A(net2802));
 sg13g2_antennanp ANTENNA_328 (.A(net2802));
 sg13g2_antennanp ANTENNA_329 (.A(net2802));
 sg13g2_antennanp ANTENNA_330 (.A(net2802));
 sg13g2_antennanp ANTENNA_331 (.A(net2802));
 sg13g2_antennanp ANTENNA_332 (.A(net2802));
 sg13g2_antennanp ANTENNA_333 (.A(net2802));
 sg13g2_antennanp ANTENNA_334 (.A(net2802));
 sg13g2_antennanp ANTENNA_335 (.A(net2802));
 sg13g2_antennanp ANTENNA_336 (.A(net2802));
 sg13g2_antennanp ANTENNA_337 (.A(net2802));
 sg13g2_antennanp ANTENNA_338 (.A(net2802));
 sg13g2_antennanp ANTENNA_339 (.A(net2802));
 sg13g2_antennanp ANTENNA_340 (.A(net2802));
 sg13g2_antennanp ANTENNA_341 (.A(net2802));
 sg13g2_antennanp ANTENNA_342 (.A(net2802));
 sg13g2_antennanp ANTENNA_343 (.A(net2802));
 sg13g2_antennanp ANTENNA_344 (.A(net2802));
 sg13g2_antennanp ANTENNA_345 (.A(net2802));
 sg13g2_antennanp ANTENNA_346 (.A(net2802));
 sg13g2_antennanp ANTENNA_347 (.A(net2802));
 sg13g2_antennanp ANTENNA_348 (.A(net2802));
 sg13g2_antennanp ANTENNA_349 (.A(net2802));
 sg13g2_antennanp ANTENNA_350 (.A(net2802));
 sg13g2_antennanp ANTENNA_351 (.A(net2802));
 sg13g2_antennanp ANTENNA_352 (.A(net2802));
 sg13g2_antennanp ANTENNA_353 (.A(net2802));
 sg13g2_antennanp ANTENNA_354 (.A(net2802));
 sg13g2_antennanp ANTENNA_355 (.A(net2802));
 sg13g2_antennanp ANTENNA_356 (.A(net2802));
 sg13g2_antennanp ANTENNA_357 (.A(net2802));
 sg13g2_antennanp ANTENNA_358 (.A(net2802));
 sg13g2_antennanp ANTENNA_359 (.A(net2802));
 sg13g2_antennanp ANTENNA_360 (.A(net2802));
 sg13g2_antennanp ANTENNA_361 (.A(net2802));
 sg13g2_antennanp ANTENNA_362 (.A(net2802));
 sg13g2_antennanp ANTENNA_363 (.A(net2802));
 sg13g2_antennanp ANTENNA_364 (.A(net2817));
 sg13g2_antennanp ANTENNA_365 (.A(net2817));
 sg13g2_antennanp ANTENNA_366 (.A(net2817));
 sg13g2_antennanp ANTENNA_367 (.A(net2817));
 sg13g2_antennanp ANTENNA_368 (.A(net2817));
 sg13g2_antennanp ANTENNA_369 (.A(net2817));
 sg13g2_antennanp ANTENNA_370 (.A(net2817));
 sg13g2_antennanp ANTENNA_371 (.A(net2817));
 sg13g2_antennanp ANTENNA_372 (.A(net2850));
 sg13g2_antennanp ANTENNA_373 (.A(net2850));
 sg13g2_antennanp ANTENNA_374 (.A(net2850));
 sg13g2_antennanp ANTENNA_375 (.A(net2850));
 sg13g2_antennanp ANTENNA_376 (.A(net2850));
 sg13g2_antennanp ANTENNA_377 (.A(net2850));
 sg13g2_antennanp ANTENNA_378 (.A(net2850));
 sg13g2_antennanp ANTENNA_379 (.A(net2850));
 sg13g2_antennanp ANTENNA_380 (.A(net2880));
 sg13g2_antennanp ANTENNA_381 (.A(net2880));
 sg13g2_antennanp ANTENNA_382 (.A(net2880));
 sg13g2_antennanp ANTENNA_383 (.A(net2880));
 sg13g2_antennanp ANTENNA_384 (.A(net2880));
 sg13g2_antennanp ANTENNA_385 (.A(net2880));
 sg13g2_antennanp ANTENNA_386 (.A(net2880));
 sg13g2_antennanp ANTENNA_387 (.A(net2880));
 sg13g2_antennanp ANTENNA_388 (.A(net2880));
 sg13g2_antennanp ANTENNA_389 (.A(net2880));
 sg13g2_antennanp ANTENNA_390 (.A(_00472_));
 sg13g2_antennanp ANTENNA_391 (.A(_00472_));
 sg13g2_antennanp ANTENNA_392 (.A(_05847_));
 sg13g2_antennanp ANTENNA_393 (.A(_05847_));
 sg13g2_antennanp ANTENNA_394 (.A(_05847_));
 sg13g2_antennanp ANTENNA_395 (.A(_05847_));
 sg13g2_antennanp ANTENNA_396 (.A(_05847_));
 sg13g2_antennanp ANTENNA_397 (.A(_05847_));
 sg13g2_antennanp ANTENNA_398 (.A(_05847_));
 sg13g2_antennanp ANTENNA_399 (.A(_05847_));
 sg13g2_antennanp ANTENNA_400 (.A(_05847_));
 sg13g2_antennanp ANTENNA_401 (.A(_05847_));
 sg13g2_antennanp ANTENNA_402 (.A(_05847_));
 sg13g2_antennanp ANTENNA_403 (.A(_05847_));
 sg13g2_antennanp ANTENNA_404 (.A(_05847_));
 sg13g2_antennanp ANTENNA_405 (.A(_05858_));
 sg13g2_antennanp ANTENNA_406 (.A(_05858_));
 sg13g2_antennanp ANTENNA_407 (.A(_05858_));
 sg13g2_antennanp ANTENNA_408 (.A(clk));
 sg13g2_antennanp ANTENNA_409 (.A(clk));
 sg13g2_antennanp ANTENNA_410 (.A(\net.in[70] ));
 sg13g2_antennanp ANTENNA_411 (.A(\net.in[70] ));
 sg13g2_antennanp ANTENNA_412 (.A(\net.in[70] ));
 sg13g2_antennanp ANTENNA_413 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_414 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_415 (.A(net2199));
 sg13g2_antennanp ANTENNA_416 (.A(net2199));
 sg13g2_antennanp ANTENNA_417 (.A(net2199));
 sg13g2_antennanp ANTENNA_418 (.A(net2199));
 sg13g2_antennanp ANTENNA_419 (.A(net2199));
 sg13g2_antennanp ANTENNA_420 (.A(net2199));
 sg13g2_antennanp ANTENNA_421 (.A(net2199));
 sg13g2_antennanp ANTENNA_422 (.A(net2199));
 sg13g2_antennanp ANTENNA_423 (.A(net2199));
 sg13g2_antennanp ANTENNA_424 (.A(net2199));
 sg13g2_antennanp ANTENNA_425 (.A(net2199));
 sg13g2_antennanp ANTENNA_426 (.A(net2199));
 sg13g2_antennanp ANTENNA_427 (.A(net2199));
 sg13g2_antennanp ANTENNA_428 (.A(net2199));
 sg13g2_antennanp ANTENNA_429 (.A(net2199));
 sg13g2_antennanp ANTENNA_430 (.A(net2199));
 sg13g2_antennanp ANTENNA_431 (.A(net2199));
 sg13g2_antennanp ANTENNA_432 (.A(net2199));
 sg13g2_antennanp ANTENNA_433 (.A(net2199));
 sg13g2_antennanp ANTENNA_434 (.A(net2199));
 sg13g2_antennanp ANTENNA_435 (.A(net2199));
 sg13g2_antennanp ANTENNA_436 (.A(net2199));
 sg13g2_antennanp ANTENNA_437 (.A(net2199));
 sg13g2_antennanp ANTENNA_438 (.A(net2199));
 sg13g2_antennanp ANTENNA_439 (.A(net2199));
 sg13g2_antennanp ANTENNA_440 (.A(net2199));
 sg13g2_antennanp ANTENNA_441 (.A(net2199));
 sg13g2_antennanp ANTENNA_442 (.A(net2199));
 sg13g2_antennanp ANTENNA_443 (.A(net2199));
 sg13g2_antennanp ANTENNA_444 (.A(net2199));
 sg13g2_antennanp ANTENNA_445 (.A(net2199));
 sg13g2_antennanp ANTENNA_446 (.A(net2199));
 sg13g2_antennanp ANTENNA_447 (.A(net2199));
 sg13g2_antennanp ANTENNA_448 (.A(net2199));
 sg13g2_antennanp ANTENNA_449 (.A(net2199));
 sg13g2_antennanp ANTENNA_450 (.A(net2199));
 sg13g2_antennanp ANTENNA_451 (.A(net2221));
 sg13g2_antennanp ANTENNA_452 (.A(net2221));
 sg13g2_antennanp ANTENNA_453 (.A(net2221));
 sg13g2_antennanp ANTENNA_454 (.A(net2221));
 sg13g2_antennanp ANTENNA_455 (.A(net2221));
 sg13g2_antennanp ANTENNA_456 (.A(net2221));
 sg13g2_antennanp ANTENNA_457 (.A(net2221));
 sg13g2_antennanp ANTENNA_458 (.A(net2221));
 sg13g2_antennanp ANTENNA_459 (.A(net2221));
 sg13g2_antennanp ANTENNA_460 (.A(net2221));
 sg13g2_antennanp ANTENNA_461 (.A(net2221));
 sg13g2_antennanp ANTENNA_462 (.A(net2221));
 sg13g2_antennanp ANTENNA_463 (.A(net2221));
 sg13g2_antennanp ANTENNA_464 (.A(net2221));
 sg13g2_antennanp ANTENNA_465 (.A(net2221));
 sg13g2_antennanp ANTENNA_466 (.A(net2239));
 sg13g2_antennanp ANTENNA_467 (.A(net2239));
 sg13g2_antennanp ANTENNA_468 (.A(net2239));
 sg13g2_antennanp ANTENNA_469 (.A(net2239));
 sg13g2_antennanp ANTENNA_470 (.A(net2239));
 sg13g2_antennanp ANTENNA_471 (.A(net2239));
 sg13g2_antennanp ANTENNA_472 (.A(net2239));
 sg13g2_antennanp ANTENNA_473 (.A(net2239));
 sg13g2_antennanp ANTENNA_474 (.A(net2239));
 sg13g2_antennanp ANTENNA_475 (.A(net2239));
 sg13g2_antennanp ANTENNA_476 (.A(net2239));
 sg13g2_antennanp ANTENNA_477 (.A(net2239));
 sg13g2_antennanp ANTENNA_478 (.A(net2239));
 sg13g2_antennanp ANTENNA_479 (.A(net2239));
 sg13g2_antennanp ANTENNA_480 (.A(net2266));
 sg13g2_antennanp ANTENNA_481 (.A(net2266));
 sg13g2_antennanp ANTENNA_482 (.A(net2266));
 sg13g2_antennanp ANTENNA_483 (.A(net2266));
 sg13g2_antennanp ANTENNA_484 (.A(net2266));
 sg13g2_antennanp ANTENNA_485 (.A(net2266));
 sg13g2_antennanp ANTENNA_486 (.A(net2266));
 sg13g2_antennanp ANTENNA_487 (.A(net2266));
 sg13g2_antennanp ANTENNA_488 (.A(net2266));
 sg13g2_antennanp ANTENNA_489 (.A(net2266));
 sg13g2_antennanp ANTENNA_490 (.A(net2266));
 sg13g2_antennanp ANTENNA_491 (.A(net2266));
 sg13g2_antennanp ANTENNA_492 (.A(net2281));
 sg13g2_antennanp ANTENNA_493 (.A(net2281));
 sg13g2_antennanp ANTENNA_494 (.A(net2281));
 sg13g2_antennanp ANTENNA_495 (.A(net2281));
 sg13g2_antennanp ANTENNA_496 (.A(net2281));
 sg13g2_antennanp ANTENNA_497 (.A(net2281));
 sg13g2_antennanp ANTENNA_498 (.A(net2281));
 sg13g2_antennanp ANTENNA_499 (.A(net2281));
 sg13g2_antennanp ANTENNA_500 (.A(net2281));
 sg13g2_antennanp ANTENNA_501 (.A(net2281));
 sg13g2_antennanp ANTENNA_502 (.A(net2281));
 sg13g2_antennanp ANTENNA_503 (.A(net2281));
 sg13g2_antennanp ANTENNA_504 (.A(net2281));
 sg13g2_antennanp ANTENNA_505 (.A(net2281));
 sg13g2_antennanp ANTENNA_506 (.A(net2284));
 sg13g2_antennanp ANTENNA_507 (.A(net2284));
 sg13g2_antennanp ANTENNA_508 (.A(net2284));
 sg13g2_antennanp ANTENNA_509 (.A(net2284));
 sg13g2_antennanp ANTENNA_510 (.A(net2284));
 sg13g2_antennanp ANTENNA_511 (.A(net2403));
 sg13g2_antennanp ANTENNA_512 (.A(net2403));
 sg13g2_antennanp ANTENNA_513 (.A(net2403));
 sg13g2_antennanp ANTENNA_514 (.A(net2403));
 sg13g2_antennanp ANTENNA_515 (.A(net2403));
 sg13g2_antennanp ANTENNA_516 (.A(net2403));
 sg13g2_antennanp ANTENNA_517 (.A(net2403));
 sg13g2_antennanp ANTENNA_518 (.A(net2403));
 sg13g2_antennanp ANTENNA_519 (.A(net2403));
 sg13g2_antennanp ANTENNA_520 (.A(net2403));
 sg13g2_antennanp ANTENNA_521 (.A(net2403));
 sg13g2_antennanp ANTENNA_522 (.A(net2403));
 sg13g2_antennanp ANTENNA_523 (.A(net2403));
 sg13g2_antennanp ANTENNA_524 (.A(net2403));
 sg13g2_antennanp ANTENNA_525 (.A(net2403));
 sg13g2_antennanp ANTENNA_526 (.A(net2403));
 sg13g2_antennanp ANTENNA_527 (.A(net2403));
 sg13g2_antennanp ANTENNA_528 (.A(net2403));
 sg13g2_antennanp ANTENNA_529 (.A(net2403));
 sg13g2_antennanp ANTENNA_530 (.A(net2403));
 sg13g2_antennanp ANTENNA_531 (.A(net2462));
 sg13g2_antennanp ANTENNA_532 (.A(net2462));
 sg13g2_antennanp ANTENNA_533 (.A(net2462));
 sg13g2_antennanp ANTENNA_534 (.A(net2462));
 sg13g2_antennanp ANTENNA_535 (.A(net2462));
 sg13g2_antennanp ANTENNA_536 (.A(net2462));
 sg13g2_antennanp ANTENNA_537 (.A(net2462));
 sg13g2_antennanp ANTENNA_538 (.A(net2462));
 sg13g2_antennanp ANTENNA_539 (.A(net2465));
 sg13g2_antennanp ANTENNA_540 (.A(net2465));
 sg13g2_antennanp ANTENNA_541 (.A(net2465));
 sg13g2_antennanp ANTENNA_542 (.A(net2465));
 sg13g2_antennanp ANTENNA_543 (.A(net2480));
 sg13g2_antennanp ANTENNA_544 (.A(net2480));
 sg13g2_antennanp ANTENNA_545 (.A(net2480));
 sg13g2_antennanp ANTENNA_546 (.A(net2480));
 sg13g2_antennanp ANTENNA_547 (.A(net2480));
 sg13g2_antennanp ANTENNA_548 (.A(net2480));
 sg13g2_antennanp ANTENNA_549 (.A(net2480));
 sg13g2_antennanp ANTENNA_550 (.A(net2480));
 sg13g2_antennanp ANTENNA_551 (.A(net2480));
 sg13g2_antennanp ANTENNA_552 (.A(net2480));
 sg13g2_antennanp ANTENNA_553 (.A(net2480));
 sg13g2_antennanp ANTENNA_554 (.A(net2480));
 sg13g2_antennanp ANTENNA_555 (.A(net2480));
 sg13g2_antennanp ANTENNA_556 (.A(net2480));
 sg13g2_antennanp ANTENNA_557 (.A(net2480));
 sg13g2_antennanp ANTENNA_558 (.A(net2480));
 sg13g2_antennanp ANTENNA_559 (.A(net2480));
 sg13g2_antennanp ANTENNA_560 (.A(net2480));
 sg13g2_antennanp ANTENNA_561 (.A(net2480));
 sg13g2_antennanp ANTENNA_562 (.A(net2480));
 sg13g2_antennanp ANTENNA_563 (.A(net2480));
 sg13g2_antennanp ANTENNA_564 (.A(net2480));
 sg13g2_antennanp ANTENNA_565 (.A(net2501));
 sg13g2_antennanp ANTENNA_566 (.A(net2501));
 sg13g2_antennanp ANTENNA_567 (.A(net2501));
 sg13g2_antennanp ANTENNA_568 (.A(net2501));
 sg13g2_antennanp ANTENNA_569 (.A(net2501));
 sg13g2_antennanp ANTENNA_570 (.A(net2501));
 sg13g2_antennanp ANTENNA_571 (.A(net2501));
 sg13g2_antennanp ANTENNA_572 (.A(net2501));
 sg13g2_antennanp ANTENNA_573 (.A(net2501));
 sg13g2_antennanp ANTENNA_574 (.A(net2501));
 sg13g2_antennanp ANTENNA_575 (.A(net2501));
 sg13g2_antennanp ANTENNA_576 (.A(net2501));
 sg13g2_antennanp ANTENNA_577 (.A(net2501));
 sg13g2_antennanp ANTENNA_578 (.A(net2501));
 sg13g2_antennanp ANTENNA_579 (.A(net2501));
 sg13g2_antennanp ANTENNA_580 (.A(net2501));
 sg13g2_antennanp ANTENNA_581 (.A(net2501));
 sg13g2_antennanp ANTENNA_582 (.A(net2501));
 sg13g2_antennanp ANTENNA_583 (.A(net2501));
 sg13g2_antennanp ANTENNA_584 (.A(net2501));
 sg13g2_antennanp ANTENNA_585 (.A(net2501));
 sg13g2_antennanp ANTENNA_586 (.A(net2501));
 sg13g2_antennanp ANTENNA_587 (.A(net2501));
 sg13g2_antennanp ANTENNA_588 (.A(net2501));
 sg13g2_antennanp ANTENNA_589 (.A(net2501));
 sg13g2_antennanp ANTENNA_590 (.A(net2501));
 sg13g2_antennanp ANTENNA_591 (.A(net2501));
 sg13g2_antennanp ANTENNA_592 (.A(net2501));
 sg13g2_antennanp ANTENNA_593 (.A(net2501));
 sg13g2_antennanp ANTENNA_594 (.A(net2501));
 sg13g2_antennanp ANTENNA_595 (.A(net2501));
 sg13g2_antennanp ANTENNA_596 (.A(net2501));
 sg13g2_antennanp ANTENNA_597 (.A(net2501));
 sg13g2_antennanp ANTENNA_598 (.A(net2501));
 sg13g2_antennanp ANTENNA_599 (.A(net2552));
 sg13g2_antennanp ANTENNA_600 (.A(net2552));
 sg13g2_antennanp ANTENNA_601 (.A(net2552));
 sg13g2_antennanp ANTENNA_602 (.A(net2552));
 sg13g2_antennanp ANTENNA_603 (.A(net2552));
 sg13g2_antennanp ANTENNA_604 (.A(net2552));
 sg13g2_antennanp ANTENNA_605 (.A(net2552));
 sg13g2_antennanp ANTENNA_606 (.A(net2552));
 sg13g2_antennanp ANTENNA_607 (.A(net2552));
 sg13g2_antennanp ANTENNA_608 (.A(net2552));
 sg13g2_antennanp ANTENNA_609 (.A(net2552));
 sg13g2_antennanp ANTENNA_610 (.A(net2552));
 sg13g2_antennanp ANTENNA_611 (.A(net2552));
 sg13g2_antennanp ANTENNA_612 (.A(net2552));
 sg13g2_antennanp ANTENNA_613 (.A(net2552));
 sg13g2_antennanp ANTENNA_614 (.A(net2585));
 sg13g2_antennanp ANTENNA_615 (.A(net2585));
 sg13g2_antennanp ANTENNA_616 (.A(net2585));
 sg13g2_antennanp ANTENNA_617 (.A(net2585));
 sg13g2_antennanp ANTENNA_618 (.A(net2585));
 sg13g2_antennanp ANTENNA_619 (.A(net2585));
 sg13g2_antennanp ANTENNA_620 (.A(net2585));
 sg13g2_antennanp ANTENNA_621 (.A(net2585));
 sg13g2_antennanp ANTENNA_622 (.A(net2585));
 sg13g2_antennanp ANTENNA_623 (.A(net2651));
 sg13g2_antennanp ANTENNA_624 (.A(net2651));
 sg13g2_antennanp ANTENNA_625 (.A(net2651));
 sg13g2_antennanp ANTENNA_626 (.A(net2651));
 sg13g2_antennanp ANTENNA_627 (.A(net2651));
 sg13g2_antennanp ANTENNA_628 (.A(net2651));
 sg13g2_antennanp ANTENNA_629 (.A(net2651));
 sg13g2_antennanp ANTENNA_630 (.A(net2651));
 sg13g2_antennanp ANTENNA_631 (.A(net2651));
 sg13g2_antennanp ANTENNA_632 (.A(net2651));
 sg13g2_antennanp ANTENNA_633 (.A(net2736));
 sg13g2_antennanp ANTENNA_634 (.A(net2736));
 sg13g2_antennanp ANTENNA_635 (.A(net2736));
 sg13g2_antennanp ANTENNA_636 (.A(net2736));
 sg13g2_antennanp ANTENNA_637 (.A(net2736));
 sg13g2_antennanp ANTENNA_638 (.A(net2736));
 sg13g2_antennanp ANTENNA_639 (.A(net2802));
 sg13g2_antennanp ANTENNA_640 (.A(net2802));
 sg13g2_antennanp ANTENNA_641 (.A(net2802));
 sg13g2_antennanp ANTENNA_642 (.A(net2802));
 sg13g2_antennanp ANTENNA_643 (.A(net2802));
 sg13g2_antennanp ANTENNA_644 (.A(net2802));
 sg13g2_antennanp ANTENNA_645 (.A(net2802));
 sg13g2_antennanp ANTENNA_646 (.A(net2802));
 sg13g2_antennanp ANTENNA_647 (.A(net2802));
 sg13g2_antennanp ANTENNA_648 (.A(net2802));
 sg13g2_antennanp ANTENNA_649 (.A(net2802));
 sg13g2_antennanp ANTENNA_650 (.A(net2802));
 sg13g2_antennanp ANTENNA_651 (.A(net2802));
 sg13g2_antennanp ANTENNA_652 (.A(net2802));
 sg13g2_antennanp ANTENNA_653 (.A(net2802));
 sg13g2_antennanp ANTENNA_654 (.A(net2802));
 sg13g2_antennanp ANTENNA_655 (.A(net2802));
 sg13g2_antennanp ANTENNA_656 (.A(net2802));
 sg13g2_antennanp ANTENNA_657 (.A(net2802));
 sg13g2_antennanp ANTENNA_658 (.A(net2802));
 sg13g2_antennanp ANTENNA_659 (.A(net2802));
 sg13g2_antennanp ANTENNA_660 (.A(net2802));
 sg13g2_antennanp ANTENNA_661 (.A(net2802));
 sg13g2_antennanp ANTENNA_662 (.A(net2802));
 sg13g2_antennanp ANTENNA_663 (.A(net2802));
 sg13g2_antennanp ANTENNA_664 (.A(net2802));
 sg13g2_antennanp ANTENNA_665 (.A(net2802));
 sg13g2_antennanp ANTENNA_666 (.A(net2802));
 sg13g2_antennanp ANTENNA_667 (.A(net2802));
 sg13g2_antennanp ANTENNA_668 (.A(net2802));
 sg13g2_antennanp ANTENNA_669 (.A(net2802));
 sg13g2_antennanp ANTENNA_670 (.A(net2802));
 sg13g2_antennanp ANTENNA_671 (.A(net2802));
 sg13g2_antennanp ANTENNA_672 (.A(net2802));
 sg13g2_antennanp ANTENNA_673 (.A(net2802));
 sg13g2_antennanp ANTENNA_674 (.A(net2802));
 sg13g2_antennanp ANTENNA_675 (.A(net2802));
 sg13g2_antennanp ANTENNA_676 (.A(net2802));
 sg13g2_antennanp ANTENNA_677 (.A(net2802));
 sg13g2_antennanp ANTENNA_678 (.A(net2802));
 sg13g2_antennanp ANTENNA_679 (.A(net2802));
 sg13g2_antennanp ANTENNA_680 (.A(net2802));
 sg13g2_antennanp ANTENNA_681 (.A(net2802));
 sg13g2_antennanp ANTENNA_682 (.A(net2802));
 sg13g2_antennanp ANTENNA_683 (.A(net2817));
 sg13g2_antennanp ANTENNA_684 (.A(net2817));
 sg13g2_antennanp ANTENNA_685 (.A(net2817));
 sg13g2_antennanp ANTENNA_686 (.A(net2817));
 sg13g2_antennanp ANTENNA_687 (.A(net2817));
 sg13g2_antennanp ANTENNA_688 (.A(net2817));
 sg13g2_antennanp ANTENNA_689 (.A(net2817));
 sg13g2_antennanp ANTENNA_690 (.A(net2817));
 sg13g2_antennanp ANTENNA_691 (.A(net2817));
 sg13g2_antennanp ANTENNA_692 (.A(net2817));
 sg13g2_antennanp ANTENNA_693 (.A(net2817));
 sg13g2_antennanp ANTENNA_694 (.A(net2817));
 sg13g2_antennanp ANTENNA_695 (.A(net2817));
 sg13g2_antennanp ANTENNA_696 (.A(net2817));
 sg13g2_antennanp ANTENNA_697 (.A(net2817));
 sg13g2_antennanp ANTENNA_698 (.A(net2817));
 sg13g2_antennanp ANTENNA_699 (.A(net2817));
 sg13g2_antennanp ANTENNA_700 (.A(net2817));
 sg13g2_antennanp ANTENNA_701 (.A(net2817));
 sg13g2_antennanp ANTENNA_702 (.A(net2817));
 sg13g2_antennanp ANTENNA_703 (.A(net2817));
 sg13g2_antennanp ANTENNA_704 (.A(net2817));
 sg13g2_antennanp ANTENNA_705 (.A(net2817));
 sg13g2_antennanp ANTENNA_706 (.A(net2817));
 sg13g2_antennanp ANTENNA_707 (.A(net2817));
 sg13g2_antennanp ANTENNA_708 (.A(net2817));
 sg13g2_antennanp ANTENNA_709 (.A(net2817));
 sg13g2_antennanp ANTENNA_710 (.A(net2817));
 sg13g2_antennanp ANTENNA_711 (.A(net2817));
 sg13g2_antennanp ANTENNA_712 (.A(net2817));
 sg13g2_antennanp ANTENNA_713 (.A(net2817));
 sg13g2_antennanp ANTENNA_714 (.A(net2817));
 sg13g2_antennanp ANTENNA_715 (.A(net2850));
 sg13g2_antennanp ANTENNA_716 (.A(net2850));
 sg13g2_antennanp ANTENNA_717 (.A(net2850));
 sg13g2_antennanp ANTENNA_718 (.A(net2850));
 sg13g2_antennanp ANTENNA_719 (.A(net2850));
 sg13g2_antennanp ANTENNA_720 (.A(net2850));
 sg13g2_antennanp ANTENNA_721 (.A(_00472_));
 sg13g2_antennanp ANTENNA_722 (.A(_00472_));
 sg13g2_antennanp ANTENNA_723 (.A(_05176_));
 sg13g2_antennanp ANTENNA_724 (.A(_05176_));
 sg13g2_antennanp ANTENNA_725 (.A(_05176_));
 sg13g2_antennanp ANTENNA_726 (.A(_05176_));
 sg13g2_antennanp ANTENNA_727 (.A(_05176_));
 sg13g2_antennanp ANTENNA_728 (.A(_05176_));
 sg13g2_antennanp ANTENNA_729 (.A(_05176_));
 sg13g2_antennanp ANTENNA_730 (.A(_05176_));
 sg13g2_antennanp ANTENNA_731 (.A(_05176_));
 sg13g2_antennanp ANTENNA_732 (.A(_05176_));
 sg13g2_antennanp ANTENNA_733 (.A(_05176_));
 sg13g2_antennanp ANTENNA_734 (.A(_05176_));
 sg13g2_antennanp ANTENNA_735 (.A(_05176_));
 sg13g2_antennanp ANTENNA_736 (.A(_05176_));
 sg13g2_antennanp ANTENNA_737 (.A(_05176_));
 sg13g2_antennanp ANTENNA_738 (.A(_05176_));
 sg13g2_antennanp ANTENNA_739 (.A(_05176_));
 sg13g2_antennanp ANTENNA_740 (.A(_05858_));
 sg13g2_antennanp ANTENNA_741 (.A(_05858_));
 sg13g2_antennanp ANTENNA_742 (.A(_05858_));
 sg13g2_antennanp ANTENNA_743 (.A(clk));
 sg13g2_antennanp ANTENNA_744 (.A(clk));
 sg13g2_antennanp ANTENNA_745 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_746 (.A(uio_in[7]));
 sg13g2_antennanp ANTENNA_747 (.A(net2199));
 sg13g2_antennanp ANTENNA_748 (.A(net2199));
 sg13g2_antennanp ANTENNA_749 (.A(net2199));
 sg13g2_antennanp ANTENNA_750 (.A(net2199));
 sg13g2_antennanp ANTENNA_751 (.A(net2199));
 sg13g2_antennanp ANTENNA_752 (.A(net2199));
 sg13g2_antennanp ANTENNA_753 (.A(net2199));
 sg13g2_antennanp ANTENNA_754 (.A(net2199));
 sg13g2_antennanp ANTENNA_755 (.A(net2199));
 sg13g2_antennanp ANTENNA_756 (.A(net2199));
 sg13g2_antennanp ANTENNA_757 (.A(net2199));
 sg13g2_antennanp ANTENNA_758 (.A(net2199));
 sg13g2_antennanp ANTENNA_759 (.A(net2199));
 sg13g2_antennanp ANTENNA_760 (.A(net2199));
 sg13g2_antennanp ANTENNA_761 (.A(net2199));
 sg13g2_antennanp ANTENNA_762 (.A(net2199));
 sg13g2_antennanp ANTENNA_763 (.A(net2199));
 sg13g2_antennanp ANTENNA_764 (.A(net2199));
 sg13g2_antennanp ANTENNA_765 (.A(net2266));
 sg13g2_antennanp ANTENNA_766 (.A(net2266));
 sg13g2_antennanp ANTENNA_767 (.A(net2266));
 sg13g2_antennanp ANTENNA_768 (.A(net2266));
 sg13g2_antennanp ANTENNA_769 (.A(net2266));
 sg13g2_antennanp ANTENNA_770 (.A(net2266));
 sg13g2_antennanp ANTENNA_771 (.A(net2266));
 sg13g2_antennanp ANTENNA_772 (.A(net2266));
 sg13g2_antennanp ANTENNA_773 (.A(net2266));
 sg13g2_antennanp ANTENNA_774 (.A(net2266));
 sg13g2_antennanp ANTENNA_775 (.A(net2266));
 sg13g2_antennanp ANTENNA_776 (.A(net2266));
 sg13g2_antennanp ANTENNA_777 (.A(net2284));
 sg13g2_antennanp ANTENNA_778 (.A(net2284));
 sg13g2_antennanp ANTENNA_779 (.A(net2284));
 sg13g2_antennanp ANTENNA_780 (.A(net2284));
 sg13g2_antennanp ANTENNA_781 (.A(net2284));
 sg13g2_antennanp ANTENNA_782 (.A(net2501));
 sg13g2_antennanp ANTENNA_783 (.A(net2501));
 sg13g2_antennanp ANTENNA_784 (.A(net2501));
 sg13g2_antennanp ANTENNA_785 (.A(net2501));
 sg13g2_antennanp ANTENNA_786 (.A(net2501));
 sg13g2_antennanp ANTENNA_787 (.A(net2501));
 sg13g2_antennanp ANTENNA_788 (.A(net2501));
 sg13g2_antennanp ANTENNA_789 (.A(net2501));
 sg13g2_antennanp ANTENNA_790 (.A(net2501));
 sg13g2_antennanp ANTENNA_791 (.A(net2501));
 sg13g2_antennanp ANTENNA_792 (.A(net2501));
 sg13g2_antennanp ANTENNA_793 (.A(net2501));
 sg13g2_antennanp ANTENNA_794 (.A(net2501));
 sg13g2_antennanp ANTENNA_795 (.A(net2501));
 sg13g2_antennanp ANTENNA_796 (.A(net2501));
 sg13g2_antennanp ANTENNA_797 (.A(net2501));
 sg13g2_antennanp ANTENNA_798 (.A(net2501));
 sg13g2_antennanp ANTENNA_799 (.A(net2501));
 sg13g2_antennanp ANTENNA_800 (.A(net2552));
 sg13g2_antennanp ANTENNA_801 (.A(net2552));
 sg13g2_antennanp ANTENNA_802 (.A(net2552));
 sg13g2_antennanp ANTENNA_803 (.A(net2552));
 sg13g2_antennanp ANTENNA_804 (.A(net2552));
 sg13g2_antennanp ANTENNA_805 (.A(net2552));
 sg13g2_antennanp ANTENNA_806 (.A(net2552));
 sg13g2_antennanp ANTENNA_807 (.A(net2552));
 sg13g2_antennanp ANTENNA_808 (.A(net2552));
 sg13g2_antennanp ANTENNA_809 (.A(net2552));
 sg13g2_antennanp ANTENNA_810 (.A(net2552));
 sg13g2_antennanp ANTENNA_811 (.A(net2552));
 sg13g2_antennanp ANTENNA_812 (.A(net2552));
 sg13g2_antennanp ANTENNA_813 (.A(net2552));
 sg13g2_antennanp ANTENNA_814 (.A(net2552));
 sg13g2_antennanp ANTENNA_815 (.A(net2585));
 sg13g2_antennanp ANTENNA_816 (.A(net2585));
 sg13g2_antennanp ANTENNA_817 (.A(net2585));
 sg13g2_antennanp ANTENNA_818 (.A(net2585));
 sg13g2_antennanp ANTENNA_819 (.A(net2585));
 sg13g2_antennanp ANTENNA_820 (.A(net2585));
 sg13g2_antennanp ANTENNA_821 (.A(net2585));
 sg13g2_antennanp ANTENNA_822 (.A(net2585));
 sg13g2_antennanp ANTENNA_823 (.A(net2585));
 sg13g2_antennanp ANTENNA_824 (.A(net2585));
 sg13g2_antennanp ANTENNA_825 (.A(net2850));
 sg13g2_antennanp ANTENNA_826 (.A(net2850));
 sg13g2_antennanp ANTENNA_827 (.A(net2850));
 sg13g2_antennanp ANTENNA_828 (.A(net2850));
 sg13g2_antennanp ANTENNA_829 (.A(net2850));
 sg13g2_antennanp ANTENNA_830 (.A(net2850));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_0_1029 ();
 sg13g2_decap_8 FILLER_0_1036 ();
 sg13g2_decap_8 FILLER_0_1043 ();
 sg13g2_decap_8 FILLER_0_1050 ();
 sg13g2_decap_8 FILLER_0_1057 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_decap_8 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1085 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_8 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1106 ();
 sg13g2_decap_8 FILLER_0_1113 ();
 sg13g2_decap_8 FILLER_0_1120 ();
 sg13g2_decap_8 FILLER_0_1127 ();
 sg13g2_decap_8 FILLER_0_1134 ();
 sg13g2_decap_8 FILLER_0_1141 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_decap_8 FILLER_0_1155 ();
 sg13g2_decap_8 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1169 ();
 sg13g2_decap_8 FILLER_0_1176 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_decap_8 FILLER_0_1456 ();
 sg13g2_decap_8 FILLER_0_1463 ();
 sg13g2_decap_8 FILLER_0_1470 ();
 sg13g2_decap_8 FILLER_0_1477 ();
 sg13g2_decap_8 FILLER_0_1484 ();
 sg13g2_decap_8 FILLER_0_1491 ();
 sg13g2_decap_8 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1540 ();
 sg13g2_decap_8 FILLER_0_1547 ();
 sg13g2_decap_8 FILLER_0_1554 ();
 sg13g2_decap_8 FILLER_0_1561 ();
 sg13g2_decap_8 FILLER_0_1568 ();
 sg13g2_decap_8 FILLER_0_1575 ();
 sg13g2_decap_8 FILLER_0_1582 ();
 sg13g2_decap_8 FILLER_0_1589 ();
 sg13g2_decap_8 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1603 ();
 sg13g2_decap_8 FILLER_0_1610 ();
 sg13g2_decap_8 FILLER_0_1617 ();
 sg13g2_decap_8 FILLER_0_1624 ();
 sg13g2_decap_8 FILLER_0_1631 ();
 sg13g2_decap_8 FILLER_0_1638 ();
 sg13g2_decap_8 FILLER_0_1645 ();
 sg13g2_decap_8 FILLER_0_1652 ();
 sg13g2_decap_8 FILLER_0_1659 ();
 sg13g2_decap_8 FILLER_0_1666 ();
 sg13g2_decap_8 FILLER_0_1673 ();
 sg13g2_decap_8 FILLER_0_1680 ();
 sg13g2_decap_8 FILLER_0_1687 ();
 sg13g2_decap_8 FILLER_0_1694 ();
 sg13g2_decap_8 FILLER_0_1701 ();
 sg13g2_decap_8 FILLER_0_1708 ();
 sg13g2_decap_8 FILLER_0_1715 ();
 sg13g2_decap_8 FILLER_0_1722 ();
 sg13g2_decap_8 FILLER_0_1729 ();
 sg13g2_decap_8 FILLER_0_1736 ();
 sg13g2_decap_8 FILLER_0_1743 ();
 sg13g2_decap_8 FILLER_0_1750 ();
 sg13g2_decap_8 FILLER_0_1757 ();
 sg13g2_decap_4 FILLER_0_1764 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_1_1029 ();
 sg13g2_decap_8 FILLER_1_1036 ();
 sg13g2_decap_8 FILLER_1_1043 ();
 sg13g2_decap_8 FILLER_1_1050 ();
 sg13g2_decap_8 FILLER_1_1057 ();
 sg13g2_decap_8 FILLER_1_1064 ();
 sg13g2_decap_8 FILLER_1_1071 ();
 sg13g2_decap_8 FILLER_1_1078 ();
 sg13g2_decap_8 FILLER_1_1085 ();
 sg13g2_decap_8 FILLER_1_1092 ();
 sg13g2_decap_8 FILLER_1_1099 ();
 sg13g2_decap_8 FILLER_1_1106 ();
 sg13g2_decap_8 FILLER_1_1113 ();
 sg13g2_decap_8 FILLER_1_1120 ();
 sg13g2_decap_8 FILLER_1_1127 ();
 sg13g2_decap_8 FILLER_1_1134 ();
 sg13g2_decap_8 FILLER_1_1141 ();
 sg13g2_decap_8 FILLER_1_1148 ();
 sg13g2_decap_8 FILLER_1_1155 ();
 sg13g2_decap_8 FILLER_1_1162 ();
 sg13g2_decap_8 FILLER_1_1169 ();
 sg13g2_decap_8 FILLER_1_1176 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1190 ();
 sg13g2_decap_8 FILLER_1_1197 ();
 sg13g2_decap_8 FILLER_1_1204 ();
 sg13g2_decap_8 FILLER_1_1211 ();
 sg13g2_decap_8 FILLER_1_1218 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_decap_8 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_decap_8 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1330 ();
 sg13g2_decap_8 FILLER_1_1337 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_decap_8 FILLER_1_1351 ();
 sg13g2_decap_8 FILLER_1_1358 ();
 sg13g2_decap_8 FILLER_1_1365 ();
 sg13g2_decap_8 FILLER_1_1372 ();
 sg13g2_decap_8 FILLER_1_1379 ();
 sg13g2_decap_8 FILLER_1_1386 ();
 sg13g2_decap_8 FILLER_1_1393 ();
 sg13g2_decap_8 FILLER_1_1400 ();
 sg13g2_decap_8 FILLER_1_1407 ();
 sg13g2_decap_8 FILLER_1_1414 ();
 sg13g2_decap_8 FILLER_1_1421 ();
 sg13g2_decap_8 FILLER_1_1428 ();
 sg13g2_decap_8 FILLER_1_1435 ();
 sg13g2_decap_8 FILLER_1_1442 ();
 sg13g2_decap_8 FILLER_1_1449 ();
 sg13g2_decap_8 FILLER_1_1456 ();
 sg13g2_decap_8 FILLER_1_1463 ();
 sg13g2_decap_8 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1477 ();
 sg13g2_decap_8 FILLER_1_1484 ();
 sg13g2_decap_8 FILLER_1_1491 ();
 sg13g2_decap_8 FILLER_1_1498 ();
 sg13g2_decap_8 FILLER_1_1505 ();
 sg13g2_decap_8 FILLER_1_1512 ();
 sg13g2_decap_8 FILLER_1_1519 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1561 ();
 sg13g2_decap_8 FILLER_1_1568 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_8 FILLER_1_1582 ();
 sg13g2_decap_8 FILLER_1_1589 ();
 sg13g2_decap_8 FILLER_1_1596 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_decap_8 FILLER_1_1610 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_8 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1638 ();
 sg13g2_decap_8 FILLER_1_1645 ();
 sg13g2_decap_8 FILLER_1_1652 ();
 sg13g2_decap_8 FILLER_1_1659 ();
 sg13g2_decap_8 FILLER_1_1666 ();
 sg13g2_decap_8 FILLER_1_1673 ();
 sg13g2_decap_8 FILLER_1_1680 ();
 sg13g2_decap_8 FILLER_1_1687 ();
 sg13g2_decap_8 FILLER_1_1694 ();
 sg13g2_decap_8 FILLER_1_1701 ();
 sg13g2_decap_8 FILLER_1_1708 ();
 sg13g2_decap_8 FILLER_1_1715 ();
 sg13g2_decap_8 FILLER_1_1722 ();
 sg13g2_decap_8 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1736 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_decap_8 FILLER_1_1750 ();
 sg13g2_decap_8 FILLER_1_1757 ();
 sg13g2_decap_4 FILLER_1_1764 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1036 ();
 sg13g2_decap_8 FILLER_2_1043 ();
 sg13g2_decap_8 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1057 ();
 sg13g2_decap_8 FILLER_2_1064 ();
 sg13g2_decap_8 FILLER_2_1071 ();
 sg13g2_decap_8 FILLER_2_1078 ();
 sg13g2_decap_8 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1092 ();
 sg13g2_decap_8 FILLER_2_1099 ();
 sg13g2_decap_8 FILLER_2_1106 ();
 sg13g2_decap_8 FILLER_2_1113 ();
 sg13g2_decap_8 FILLER_2_1120 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_8 FILLER_2_1134 ();
 sg13g2_decap_8 FILLER_2_1141 ();
 sg13g2_decap_8 FILLER_2_1148 ();
 sg13g2_decap_8 FILLER_2_1155 ();
 sg13g2_decap_8 FILLER_2_1162 ();
 sg13g2_decap_8 FILLER_2_1169 ();
 sg13g2_decap_8 FILLER_2_1176 ();
 sg13g2_decap_8 FILLER_2_1183 ();
 sg13g2_decap_8 FILLER_2_1190 ();
 sg13g2_decap_8 FILLER_2_1197 ();
 sg13g2_decap_8 FILLER_2_1204 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_decap_8 FILLER_2_1218 ();
 sg13g2_decap_8 FILLER_2_1225 ();
 sg13g2_decap_8 FILLER_2_1232 ();
 sg13g2_decap_8 FILLER_2_1239 ();
 sg13g2_decap_8 FILLER_2_1246 ();
 sg13g2_decap_8 FILLER_2_1253 ();
 sg13g2_decap_8 FILLER_2_1260 ();
 sg13g2_decap_8 FILLER_2_1267 ();
 sg13g2_decap_8 FILLER_2_1274 ();
 sg13g2_decap_8 FILLER_2_1281 ();
 sg13g2_decap_8 FILLER_2_1288 ();
 sg13g2_decap_8 FILLER_2_1295 ();
 sg13g2_decap_8 FILLER_2_1302 ();
 sg13g2_decap_8 FILLER_2_1309 ();
 sg13g2_decap_8 FILLER_2_1316 ();
 sg13g2_decap_8 FILLER_2_1323 ();
 sg13g2_decap_8 FILLER_2_1330 ();
 sg13g2_decap_8 FILLER_2_1337 ();
 sg13g2_decap_8 FILLER_2_1344 ();
 sg13g2_decap_8 FILLER_2_1351 ();
 sg13g2_decap_8 FILLER_2_1358 ();
 sg13g2_decap_8 FILLER_2_1365 ();
 sg13g2_decap_8 FILLER_2_1372 ();
 sg13g2_decap_8 FILLER_2_1379 ();
 sg13g2_decap_8 FILLER_2_1386 ();
 sg13g2_decap_8 FILLER_2_1393 ();
 sg13g2_decap_8 FILLER_2_1400 ();
 sg13g2_decap_8 FILLER_2_1407 ();
 sg13g2_decap_8 FILLER_2_1414 ();
 sg13g2_decap_8 FILLER_2_1421 ();
 sg13g2_decap_8 FILLER_2_1428 ();
 sg13g2_decap_8 FILLER_2_1435 ();
 sg13g2_decap_8 FILLER_2_1442 ();
 sg13g2_decap_8 FILLER_2_1449 ();
 sg13g2_decap_8 FILLER_2_1456 ();
 sg13g2_decap_8 FILLER_2_1463 ();
 sg13g2_decap_8 FILLER_2_1470 ();
 sg13g2_decap_8 FILLER_2_1477 ();
 sg13g2_decap_8 FILLER_2_1484 ();
 sg13g2_decap_8 FILLER_2_1491 ();
 sg13g2_decap_8 FILLER_2_1498 ();
 sg13g2_decap_8 FILLER_2_1505 ();
 sg13g2_decap_8 FILLER_2_1512 ();
 sg13g2_decap_8 FILLER_2_1519 ();
 sg13g2_decap_8 FILLER_2_1526 ();
 sg13g2_decap_8 FILLER_2_1533 ();
 sg13g2_decap_8 FILLER_2_1540 ();
 sg13g2_decap_8 FILLER_2_1547 ();
 sg13g2_decap_8 FILLER_2_1554 ();
 sg13g2_decap_8 FILLER_2_1561 ();
 sg13g2_decap_8 FILLER_2_1568 ();
 sg13g2_decap_8 FILLER_2_1575 ();
 sg13g2_decap_8 FILLER_2_1582 ();
 sg13g2_decap_8 FILLER_2_1589 ();
 sg13g2_decap_8 FILLER_2_1596 ();
 sg13g2_decap_8 FILLER_2_1603 ();
 sg13g2_decap_8 FILLER_2_1610 ();
 sg13g2_decap_8 FILLER_2_1617 ();
 sg13g2_decap_8 FILLER_2_1624 ();
 sg13g2_decap_8 FILLER_2_1631 ();
 sg13g2_decap_8 FILLER_2_1638 ();
 sg13g2_decap_8 FILLER_2_1645 ();
 sg13g2_decap_8 FILLER_2_1652 ();
 sg13g2_decap_8 FILLER_2_1659 ();
 sg13g2_decap_8 FILLER_2_1666 ();
 sg13g2_decap_8 FILLER_2_1673 ();
 sg13g2_decap_8 FILLER_2_1680 ();
 sg13g2_decap_8 FILLER_2_1687 ();
 sg13g2_decap_8 FILLER_2_1694 ();
 sg13g2_decap_8 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1708 ();
 sg13g2_decap_8 FILLER_2_1715 ();
 sg13g2_decap_8 FILLER_2_1722 ();
 sg13g2_decap_8 FILLER_2_1729 ();
 sg13g2_decap_8 FILLER_2_1736 ();
 sg13g2_decap_8 FILLER_2_1743 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_8 FILLER_2_1757 ();
 sg13g2_decap_4 FILLER_2_1764 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_8 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_decap_8 FILLER_3_1029 ();
 sg13g2_decap_8 FILLER_3_1036 ();
 sg13g2_decap_8 FILLER_3_1043 ();
 sg13g2_decap_8 FILLER_3_1050 ();
 sg13g2_decap_8 FILLER_3_1057 ();
 sg13g2_decap_8 FILLER_3_1064 ();
 sg13g2_decap_8 FILLER_3_1071 ();
 sg13g2_decap_8 FILLER_3_1078 ();
 sg13g2_decap_8 FILLER_3_1085 ();
 sg13g2_decap_8 FILLER_3_1092 ();
 sg13g2_decap_8 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1113 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_decap_8 FILLER_3_1134 ();
 sg13g2_decap_8 FILLER_3_1141 ();
 sg13g2_decap_8 FILLER_3_1148 ();
 sg13g2_decap_8 FILLER_3_1155 ();
 sg13g2_decap_8 FILLER_3_1162 ();
 sg13g2_decap_8 FILLER_3_1169 ();
 sg13g2_decap_8 FILLER_3_1176 ();
 sg13g2_decap_8 FILLER_3_1183 ();
 sg13g2_decap_8 FILLER_3_1190 ();
 sg13g2_decap_8 FILLER_3_1197 ();
 sg13g2_decap_8 FILLER_3_1204 ();
 sg13g2_decap_8 FILLER_3_1211 ();
 sg13g2_decap_8 FILLER_3_1218 ();
 sg13g2_decap_8 FILLER_3_1225 ();
 sg13g2_decap_8 FILLER_3_1232 ();
 sg13g2_decap_8 FILLER_3_1239 ();
 sg13g2_decap_8 FILLER_3_1246 ();
 sg13g2_decap_8 FILLER_3_1253 ();
 sg13g2_decap_8 FILLER_3_1260 ();
 sg13g2_decap_8 FILLER_3_1267 ();
 sg13g2_decap_8 FILLER_3_1274 ();
 sg13g2_decap_8 FILLER_3_1281 ();
 sg13g2_decap_8 FILLER_3_1288 ();
 sg13g2_decap_8 FILLER_3_1295 ();
 sg13g2_decap_8 FILLER_3_1302 ();
 sg13g2_decap_8 FILLER_3_1309 ();
 sg13g2_decap_8 FILLER_3_1316 ();
 sg13g2_decap_8 FILLER_3_1323 ();
 sg13g2_decap_8 FILLER_3_1330 ();
 sg13g2_decap_8 FILLER_3_1337 ();
 sg13g2_decap_8 FILLER_3_1344 ();
 sg13g2_decap_8 FILLER_3_1351 ();
 sg13g2_decap_8 FILLER_3_1358 ();
 sg13g2_decap_8 FILLER_3_1365 ();
 sg13g2_decap_8 FILLER_3_1372 ();
 sg13g2_decap_8 FILLER_3_1379 ();
 sg13g2_decap_8 FILLER_3_1386 ();
 sg13g2_decap_8 FILLER_3_1393 ();
 sg13g2_decap_8 FILLER_3_1400 ();
 sg13g2_decap_8 FILLER_3_1407 ();
 sg13g2_decap_8 FILLER_3_1414 ();
 sg13g2_decap_8 FILLER_3_1421 ();
 sg13g2_decap_8 FILLER_3_1428 ();
 sg13g2_decap_8 FILLER_3_1435 ();
 sg13g2_decap_8 FILLER_3_1442 ();
 sg13g2_decap_8 FILLER_3_1449 ();
 sg13g2_decap_8 FILLER_3_1456 ();
 sg13g2_decap_8 FILLER_3_1463 ();
 sg13g2_decap_8 FILLER_3_1470 ();
 sg13g2_decap_8 FILLER_3_1477 ();
 sg13g2_decap_8 FILLER_3_1484 ();
 sg13g2_decap_8 FILLER_3_1491 ();
 sg13g2_decap_8 FILLER_3_1498 ();
 sg13g2_decap_8 FILLER_3_1505 ();
 sg13g2_decap_8 FILLER_3_1512 ();
 sg13g2_decap_8 FILLER_3_1519 ();
 sg13g2_decap_8 FILLER_3_1526 ();
 sg13g2_decap_8 FILLER_3_1533 ();
 sg13g2_decap_8 FILLER_3_1540 ();
 sg13g2_decap_8 FILLER_3_1547 ();
 sg13g2_decap_8 FILLER_3_1554 ();
 sg13g2_decap_8 FILLER_3_1561 ();
 sg13g2_decap_8 FILLER_3_1568 ();
 sg13g2_decap_8 FILLER_3_1575 ();
 sg13g2_decap_8 FILLER_3_1582 ();
 sg13g2_decap_8 FILLER_3_1589 ();
 sg13g2_decap_8 FILLER_3_1596 ();
 sg13g2_decap_8 FILLER_3_1603 ();
 sg13g2_decap_8 FILLER_3_1610 ();
 sg13g2_decap_8 FILLER_3_1617 ();
 sg13g2_decap_8 FILLER_3_1624 ();
 sg13g2_decap_8 FILLER_3_1631 ();
 sg13g2_decap_8 FILLER_3_1638 ();
 sg13g2_decap_8 FILLER_3_1645 ();
 sg13g2_decap_8 FILLER_3_1652 ();
 sg13g2_decap_8 FILLER_3_1659 ();
 sg13g2_decap_8 FILLER_3_1666 ();
 sg13g2_decap_8 FILLER_3_1673 ();
 sg13g2_decap_8 FILLER_3_1680 ();
 sg13g2_decap_8 FILLER_3_1687 ();
 sg13g2_decap_8 FILLER_3_1694 ();
 sg13g2_decap_8 FILLER_3_1701 ();
 sg13g2_decap_8 FILLER_3_1708 ();
 sg13g2_decap_8 FILLER_3_1715 ();
 sg13g2_decap_8 FILLER_3_1722 ();
 sg13g2_decap_8 FILLER_3_1729 ();
 sg13g2_decap_8 FILLER_3_1736 ();
 sg13g2_decap_8 FILLER_3_1743 ();
 sg13g2_decap_8 FILLER_3_1750 ();
 sg13g2_decap_8 FILLER_3_1757 ();
 sg13g2_decap_4 FILLER_3_1764 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_decap_8 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_decap_8 FILLER_4_924 ();
 sg13g2_decap_8 FILLER_4_931 ();
 sg13g2_decap_8 FILLER_4_938 ();
 sg13g2_decap_8 FILLER_4_945 ();
 sg13g2_decap_8 FILLER_4_952 ();
 sg13g2_decap_8 FILLER_4_959 ();
 sg13g2_decap_8 FILLER_4_966 ();
 sg13g2_decap_8 FILLER_4_973 ();
 sg13g2_decap_8 FILLER_4_980 ();
 sg13g2_decap_8 FILLER_4_987 ();
 sg13g2_decap_8 FILLER_4_994 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1015 ();
 sg13g2_decap_8 FILLER_4_1022 ();
 sg13g2_decap_8 FILLER_4_1029 ();
 sg13g2_decap_8 FILLER_4_1036 ();
 sg13g2_decap_8 FILLER_4_1043 ();
 sg13g2_decap_8 FILLER_4_1050 ();
 sg13g2_decap_8 FILLER_4_1057 ();
 sg13g2_decap_8 FILLER_4_1064 ();
 sg13g2_decap_8 FILLER_4_1071 ();
 sg13g2_decap_8 FILLER_4_1078 ();
 sg13g2_decap_8 FILLER_4_1085 ();
 sg13g2_decap_8 FILLER_4_1092 ();
 sg13g2_decap_8 FILLER_4_1099 ();
 sg13g2_decap_8 FILLER_4_1106 ();
 sg13g2_decap_8 FILLER_4_1113 ();
 sg13g2_decap_8 FILLER_4_1120 ();
 sg13g2_decap_8 FILLER_4_1127 ();
 sg13g2_decap_8 FILLER_4_1134 ();
 sg13g2_decap_8 FILLER_4_1141 ();
 sg13g2_decap_8 FILLER_4_1148 ();
 sg13g2_decap_8 FILLER_4_1155 ();
 sg13g2_decap_8 FILLER_4_1162 ();
 sg13g2_decap_8 FILLER_4_1169 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_decap_8 FILLER_4_1183 ();
 sg13g2_decap_8 FILLER_4_1190 ();
 sg13g2_decap_8 FILLER_4_1197 ();
 sg13g2_decap_8 FILLER_4_1204 ();
 sg13g2_decap_8 FILLER_4_1211 ();
 sg13g2_decap_8 FILLER_4_1218 ();
 sg13g2_decap_8 FILLER_4_1225 ();
 sg13g2_decap_8 FILLER_4_1232 ();
 sg13g2_decap_8 FILLER_4_1239 ();
 sg13g2_decap_8 FILLER_4_1246 ();
 sg13g2_decap_8 FILLER_4_1253 ();
 sg13g2_decap_8 FILLER_4_1260 ();
 sg13g2_decap_8 FILLER_4_1267 ();
 sg13g2_decap_8 FILLER_4_1274 ();
 sg13g2_decap_8 FILLER_4_1281 ();
 sg13g2_decap_8 FILLER_4_1288 ();
 sg13g2_decap_8 FILLER_4_1295 ();
 sg13g2_decap_8 FILLER_4_1302 ();
 sg13g2_decap_8 FILLER_4_1309 ();
 sg13g2_decap_8 FILLER_4_1316 ();
 sg13g2_decap_8 FILLER_4_1323 ();
 sg13g2_decap_8 FILLER_4_1330 ();
 sg13g2_decap_8 FILLER_4_1337 ();
 sg13g2_decap_8 FILLER_4_1344 ();
 sg13g2_decap_8 FILLER_4_1351 ();
 sg13g2_decap_8 FILLER_4_1358 ();
 sg13g2_decap_8 FILLER_4_1365 ();
 sg13g2_decap_8 FILLER_4_1372 ();
 sg13g2_decap_8 FILLER_4_1379 ();
 sg13g2_decap_8 FILLER_4_1386 ();
 sg13g2_decap_8 FILLER_4_1393 ();
 sg13g2_decap_8 FILLER_4_1400 ();
 sg13g2_decap_8 FILLER_4_1407 ();
 sg13g2_decap_8 FILLER_4_1414 ();
 sg13g2_decap_8 FILLER_4_1421 ();
 sg13g2_decap_8 FILLER_4_1428 ();
 sg13g2_decap_8 FILLER_4_1435 ();
 sg13g2_decap_8 FILLER_4_1442 ();
 sg13g2_decap_8 FILLER_4_1449 ();
 sg13g2_decap_8 FILLER_4_1456 ();
 sg13g2_decap_8 FILLER_4_1463 ();
 sg13g2_decap_8 FILLER_4_1470 ();
 sg13g2_decap_8 FILLER_4_1477 ();
 sg13g2_decap_8 FILLER_4_1484 ();
 sg13g2_decap_8 FILLER_4_1491 ();
 sg13g2_decap_8 FILLER_4_1498 ();
 sg13g2_decap_8 FILLER_4_1505 ();
 sg13g2_decap_8 FILLER_4_1512 ();
 sg13g2_decap_8 FILLER_4_1519 ();
 sg13g2_decap_8 FILLER_4_1526 ();
 sg13g2_decap_8 FILLER_4_1533 ();
 sg13g2_decap_8 FILLER_4_1540 ();
 sg13g2_decap_8 FILLER_4_1547 ();
 sg13g2_decap_8 FILLER_4_1554 ();
 sg13g2_decap_8 FILLER_4_1561 ();
 sg13g2_decap_8 FILLER_4_1568 ();
 sg13g2_decap_8 FILLER_4_1575 ();
 sg13g2_decap_8 FILLER_4_1582 ();
 sg13g2_decap_8 FILLER_4_1589 ();
 sg13g2_decap_8 FILLER_4_1596 ();
 sg13g2_decap_8 FILLER_4_1603 ();
 sg13g2_decap_8 FILLER_4_1610 ();
 sg13g2_decap_8 FILLER_4_1617 ();
 sg13g2_decap_8 FILLER_4_1624 ();
 sg13g2_decap_8 FILLER_4_1631 ();
 sg13g2_decap_8 FILLER_4_1638 ();
 sg13g2_decap_8 FILLER_4_1645 ();
 sg13g2_decap_8 FILLER_4_1652 ();
 sg13g2_decap_8 FILLER_4_1659 ();
 sg13g2_decap_8 FILLER_4_1666 ();
 sg13g2_decap_8 FILLER_4_1673 ();
 sg13g2_decap_8 FILLER_4_1680 ();
 sg13g2_decap_8 FILLER_4_1687 ();
 sg13g2_decap_8 FILLER_4_1694 ();
 sg13g2_decap_8 FILLER_4_1701 ();
 sg13g2_decap_8 FILLER_4_1708 ();
 sg13g2_decap_8 FILLER_4_1715 ();
 sg13g2_decap_8 FILLER_4_1722 ();
 sg13g2_decap_8 FILLER_4_1729 ();
 sg13g2_decap_8 FILLER_4_1736 ();
 sg13g2_decap_8 FILLER_4_1743 ();
 sg13g2_decap_8 FILLER_4_1750 ();
 sg13g2_decap_8 FILLER_4_1757 ();
 sg13g2_decap_4 FILLER_4_1764 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_decap_8 FILLER_5_875 ();
 sg13g2_decap_8 FILLER_5_882 ();
 sg13g2_decap_8 FILLER_5_889 ();
 sg13g2_decap_8 FILLER_5_896 ();
 sg13g2_decap_8 FILLER_5_903 ();
 sg13g2_decap_8 FILLER_5_910 ();
 sg13g2_decap_8 FILLER_5_917 ();
 sg13g2_decap_8 FILLER_5_924 ();
 sg13g2_decap_8 FILLER_5_931 ();
 sg13g2_decap_8 FILLER_5_938 ();
 sg13g2_decap_8 FILLER_5_945 ();
 sg13g2_decap_8 FILLER_5_952 ();
 sg13g2_decap_8 FILLER_5_959 ();
 sg13g2_decap_8 FILLER_5_966 ();
 sg13g2_decap_8 FILLER_5_973 ();
 sg13g2_decap_8 FILLER_5_980 ();
 sg13g2_decap_8 FILLER_5_987 ();
 sg13g2_decap_8 FILLER_5_994 ();
 sg13g2_decap_8 FILLER_5_1001 ();
 sg13g2_decap_8 FILLER_5_1008 ();
 sg13g2_decap_8 FILLER_5_1015 ();
 sg13g2_decap_8 FILLER_5_1022 ();
 sg13g2_decap_8 FILLER_5_1029 ();
 sg13g2_decap_8 FILLER_5_1036 ();
 sg13g2_decap_8 FILLER_5_1043 ();
 sg13g2_decap_8 FILLER_5_1050 ();
 sg13g2_decap_8 FILLER_5_1057 ();
 sg13g2_decap_8 FILLER_5_1064 ();
 sg13g2_decap_8 FILLER_5_1071 ();
 sg13g2_decap_8 FILLER_5_1078 ();
 sg13g2_decap_8 FILLER_5_1085 ();
 sg13g2_decap_8 FILLER_5_1092 ();
 sg13g2_decap_8 FILLER_5_1099 ();
 sg13g2_decap_8 FILLER_5_1106 ();
 sg13g2_decap_8 FILLER_5_1113 ();
 sg13g2_decap_8 FILLER_5_1120 ();
 sg13g2_decap_8 FILLER_5_1127 ();
 sg13g2_decap_8 FILLER_5_1134 ();
 sg13g2_decap_8 FILLER_5_1141 ();
 sg13g2_decap_8 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1155 ();
 sg13g2_decap_8 FILLER_5_1162 ();
 sg13g2_decap_8 FILLER_5_1169 ();
 sg13g2_decap_8 FILLER_5_1176 ();
 sg13g2_decap_8 FILLER_5_1183 ();
 sg13g2_decap_8 FILLER_5_1190 ();
 sg13g2_decap_8 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1204 ();
 sg13g2_decap_8 FILLER_5_1211 ();
 sg13g2_decap_8 FILLER_5_1218 ();
 sg13g2_decap_8 FILLER_5_1225 ();
 sg13g2_decap_8 FILLER_5_1232 ();
 sg13g2_decap_8 FILLER_5_1239 ();
 sg13g2_decap_8 FILLER_5_1246 ();
 sg13g2_decap_8 FILLER_5_1253 ();
 sg13g2_decap_8 FILLER_5_1260 ();
 sg13g2_decap_8 FILLER_5_1267 ();
 sg13g2_decap_8 FILLER_5_1274 ();
 sg13g2_decap_8 FILLER_5_1281 ();
 sg13g2_decap_8 FILLER_5_1288 ();
 sg13g2_decap_8 FILLER_5_1295 ();
 sg13g2_decap_8 FILLER_5_1302 ();
 sg13g2_decap_8 FILLER_5_1309 ();
 sg13g2_decap_8 FILLER_5_1316 ();
 sg13g2_decap_8 FILLER_5_1323 ();
 sg13g2_decap_8 FILLER_5_1330 ();
 sg13g2_decap_8 FILLER_5_1337 ();
 sg13g2_decap_8 FILLER_5_1344 ();
 sg13g2_decap_8 FILLER_5_1351 ();
 sg13g2_decap_8 FILLER_5_1358 ();
 sg13g2_decap_8 FILLER_5_1365 ();
 sg13g2_decap_8 FILLER_5_1372 ();
 sg13g2_decap_8 FILLER_5_1379 ();
 sg13g2_decap_8 FILLER_5_1386 ();
 sg13g2_decap_8 FILLER_5_1393 ();
 sg13g2_decap_8 FILLER_5_1400 ();
 sg13g2_decap_8 FILLER_5_1407 ();
 sg13g2_decap_8 FILLER_5_1414 ();
 sg13g2_decap_8 FILLER_5_1421 ();
 sg13g2_decap_8 FILLER_5_1428 ();
 sg13g2_decap_8 FILLER_5_1435 ();
 sg13g2_decap_8 FILLER_5_1442 ();
 sg13g2_decap_8 FILLER_5_1449 ();
 sg13g2_decap_8 FILLER_5_1456 ();
 sg13g2_decap_8 FILLER_5_1463 ();
 sg13g2_decap_8 FILLER_5_1470 ();
 sg13g2_decap_8 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1491 ();
 sg13g2_decap_8 FILLER_5_1498 ();
 sg13g2_decap_8 FILLER_5_1505 ();
 sg13g2_decap_8 FILLER_5_1512 ();
 sg13g2_decap_8 FILLER_5_1519 ();
 sg13g2_decap_8 FILLER_5_1526 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_decap_8 FILLER_5_1540 ();
 sg13g2_decap_8 FILLER_5_1547 ();
 sg13g2_decap_8 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1561 ();
 sg13g2_decap_8 FILLER_5_1568 ();
 sg13g2_decap_8 FILLER_5_1575 ();
 sg13g2_decap_8 FILLER_5_1582 ();
 sg13g2_decap_8 FILLER_5_1589 ();
 sg13g2_decap_8 FILLER_5_1596 ();
 sg13g2_decap_8 FILLER_5_1603 ();
 sg13g2_decap_8 FILLER_5_1610 ();
 sg13g2_decap_8 FILLER_5_1617 ();
 sg13g2_decap_8 FILLER_5_1624 ();
 sg13g2_decap_8 FILLER_5_1631 ();
 sg13g2_decap_8 FILLER_5_1638 ();
 sg13g2_decap_8 FILLER_5_1645 ();
 sg13g2_decap_8 FILLER_5_1652 ();
 sg13g2_decap_8 FILLER_5_1659 ();
 sg13g2_decap_8 FILLER_5_1666 ();
 sg13g2_decap_8 FILLER_5_1673 ();
 sg13g2_decap_8 FILLER_5_1680 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_decap_8 FILLER_5_1694 ();
 sg13g2_decap_8 FILLER_5_1701 ();
 sg13g2_decap_8 FILLER_5_1708 ();
 sg13g2_decap_8 FILLER_5_1715 ();
 sg13g2_decap_8 FILLER_5_1722 ();
 sg13g2_decap_8 FILLER_5_1729 ();
 sg13g2_decap_8 FILLER_5_1736 ();
 sg13g2_decap_8 FILLER_5_1743 ();
 sg13g2_decap_8 FILLER_5_1750 ();
 sg13g2_decap_8 FILLER_5_1757 ();
 sg13g2_decap_4 FILLER_5_1764 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_decap_8 FILLER_6_875 ();
 sg13g2_decap_8 FILLER_6_882 ();
 sg13g2_decap_8 FILLER_6_889 ();
 sg13g2_decap_8 FILLER_6_896 ();
 sg13g2_decap_8 FILLER_6_903 ();
 sg13g2_decap_8 FILLER_6_910 ();
 sg13g2_decap_8 FILLER_6_917 ();
 sg13g2_decap_8 FILLER_6_924 ();
 sg13g2_decap_8 FILLER_6_931 ();
 sg13g2_decap_8 FILLER_6_938 ();
 sg13g2_decap_8 FILLER_6_945 ();
 sg13g2_decap_8 FILLER_6_952 ();
 sg13g2_decap_8 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_8 FILLER_6_1015 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_6_1029 ();
 sg13g2_decap_8 FILLER_6_1036 ();
 sg13g2_decap_8 FILLER_6_1043 ();
 sg13g2_decap_8 FILLER_6_1050 ();
 sg13g2_decap_8 FILLER_6_1057 ();
 sg13g2_decap_8 FILLER_6_1064 ();
 sg13g2_decap_8 FILLER_6_1071 ();
 sg13g2_decap_8 FILLER_6_1078 ();
 sg13g2_decap_8 FILLER_6_1085 ();
 sg13g2_decap_8 FILLER_6_1092 ();
 sg13g2_decap_8 FILLER_6_1099 ();
 sg13g2_decap_8 FILLER_6_1106 ();
 sg13g2_decap_8 FILLER_6_1113 ();
 sg13g2_decap_8 FILLER_6_1120 ();
 sg13g2_decap_8 FILLER_6_1127 ();
 sg13g2_decap_8 FILLER_6_1134 ();
 sg13g2_decap_8 FILLER_6_1141 ();
 sg13g2_decap_8 FILLER_6_1148 ();
 sg13g2_decap_8 FILLER_6_1155 ();
 sg13g2_decap_8 FILLER_6_1162 ();
 sg13g2_decap_8 FILLER_6_1169 ();
 sg13g2_decap_8 FILLER_6_1176 ();
 sg13g2_decap_8 FILLER_6_1183 ();
 sg13g2_decap_8 FILLER_6_1190 ();
 sg13g2_decap_8 FILLER_6_1197 ();
 sg13g2_decap_8 FILLER_6_1204 ();
 sg13g2_decap_8 FILLER_6_1211 ();
 sg13g2_decap_8 FILLER_6_1218 ();
 sg13g2_decap_8 FILLER_6_1225 ();
 sg13g2_decap_8 FILLER_6_1232 ();
 sg13g2_decap_8 FILLER_6_1239 ();
 sg13g2_decap_8 FILLER_6_1246 ();
 sg13g2_decap_8 FILLER_6_1253 ();
 sg13g2_decap_8 FILLER_6_1260 ();
 sg13g2_decap_8 FILLER_6_1267 ();
 sg13g2_decap_8 FILLER_6_1274 ();
 sg13g2_decap_8 FILLER_6_1281 ();
 sg13g2_decap_8 FILLER_6_1288 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_decap_8 FILLER_6_1302 ();
 sg13g2_decap_8 FILLER_6_1309 ();
 sg13g2_decap_8 FILLER_6_1316 ();
 sg13g2_decap_8 FILLER_6_1323 ();
 sg13g2_decap_8 FILLER_6_1330 ();
 sg13g2_decap_8 FILLER_6_1337 ();
 sg13g2_decap_8 FILLER_6_1344 ();
 sg13g2_decap_8 FILLER_6_1351 ();
 sg13g2_decap_8 FILLER_6_1358 ();
 sg13g2_decap_8 FILLER_6_1365 ();
 sg13g2_decap_8 FILLER_6_1372 ();
 sg13g2_decap_8 FILLER_6_1379 ();
 sg13g2_decap_8 FILLER_6_1386 ();
 sg13g2_decap_8 FILLER_6_1393 ();
 sg13g2_decap_8 FILLER_6_1400 ();
 sg13g2_decap_8 FILLER_6_1407 ();
 sg13g2_decap_8 FILLER_6_1414 ();
 sg13g2_decap_8 FILLER_6_1421 ();
 sg13g2_decap_8 FILLER_6_1428 ();
 sg13g2_decap_8 FILLER_6_1435 ();
 sg13g2_decap_8 FILLER_6_1442 ();
 sg13g2_decap_8 FILLER_6_1449 ();
 sg13g2_decap_8 FILLER_6_1456 ();
 sg13g2_decap_8 FILLER_6_1463 ();
 sg13g2_decap_8 FILLER_6_1470 ();
 sg13g2_decap_8 FILLER_6_1477 ();
 sg13g2_decap_8 FILLER_6_1484 ();
 sg13g2_decap_8 FILLER_6_1491 ();
 sg13g2_decap_8 FILLER_6_1498 ();
 sg13g2_decap_8 FILLER_6_1505 ();
 sg13g2_decap_8 FILLER_6_1512 ();
 sg13g2_decap_8 FILLER_6_1519 ();
 sg13g2_decap_8 FILLER_6_1526 ();
 sg13g2_decap_8 FILLER_6_1533 ();
 sg13g2_decap_8 FILLER_6_1540 ();
 sg13g2_decap_8 FILLER_6_1547 ();
 sg13g2_decap_8 FILLER_6_1554 ();
 sg13g2_decap_8 FILLER_6_1561 ();
 sg13g2_decap_8 FILLER_6_1568 ();
 sg13g2_decap_8 FILLER_6_1575 ();
 sg13g2_decap_8 FILLER_6_1582 ();
 sg13g2_decap_8 FILLER_6_1589 ();
 sg13g2_decap_8 FILLER_6_1596 ();
 sg13g2_decap_8 FILLER_6_1603 ();
 sg13g2_decap_8 FILLER_6_1610 ();
 sg13g2_decap_8 FILLER_6_1617 ();
 sg13g2_decap_8 FILLER_6_1624 ();
 sg13g2_decap_8 FILLER_6_1631 ();
 sg13g2_decap_8 FILLER_6_1638 ();
 sg13g2_decap_8 FILLER_6_1645 ();
 sg13g2_decap_8 FILLER_6_1652 ();
 sg13g2_decap_8 FILLER_6_1659 ();
 sg13g2_decap_8 FILLER_6_1666 ();
 sg13g2_decap_8 FILLER_6_1673 ();
 sg13g2_decap_8 FILLER_6_1680 ();
 sg13g2_decap_8 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1694 ();
 sg13g2_decap_8 FILLER_6_1701 ();
 sg13g2_decap_8 FILLER_6_1708 ();
 sg13g2_decap_8 FILLER_6_1715 ();
 sg13g2_decap_8 FILLER_6_1722 ();
 sg13g2_decap_8 FILLER_6_1729 ();
 sg13g2_decap_8 FILLER_6_1736 ();
 sg13g2_decap_8 FILLER_6_1743 ();
 sg13g2_decap_8 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1757 ();
 sg13g2_decap_4 FILLER_6_1764 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_7_1029 ();
 sg13g2_decap_8 FILLER_7_1036 ();
 sg13g2_decap_8 FILLER_7_1043 ();
 sg13g2_decap_8 FILLER_7_1050 ();
 sg13g2_decap_8 FILLER_7_1057 ();
 sg13g2_decap_8 FILLER_7_1064 ();
 sg13g2_decap_8 FILLER_7_1071 ();
 sg13g2_decap_8 FILLER_7_1078 ();
 sg13g2_decap_8 FILLER_7_1085 ();
 sg13g2_decap_8 FILLER_7_1092 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_decap_8 FILLER_7_1113 ();
 sg13g2_decap_8 FILLER_7_1120 ();
 sg13g2_decap_8 FILLER_7_1127 ();
 sg13g2_decap_8 FILLER_7_1134 ();
 sg13g2_decap_8 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1155 ();
 sg13g2_decap_8 FILLER_7_1162 ();
 sg13g2_decap_8 FILLER_7_1169 ();
 sg13g2_decap_8 FILLER_7_1176 ();
 sg13g2_decap_8 FILLER_7_1183 ();
 sg13g2_decap_8 FILLER_7_1190 ();
 sg13g2_decap_8 FILLER_7_1197 ();
 sg13g2_decap_8 FILLER_7_1204 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_decap_8 FILLER_7_1218 ();
 sg13g2_decap_8 FILLER_7_1225 ();
 sg13g2_decap_8 FILLER_7_1232 ();
 sg13g2_decap_8 FILLER_7_1239 ();
 sg13g2_decap_8 FILLER_7_1246 ();
 sg13g2_decap_8 FILLER_7_1253 ();
 sg13g2_decap_8 FILLER_7_1260 ();
 sg13g2_decap_8 FILLER_7_1267 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_decap_8 FILLER_7_1323 ();
 sg13g2_decap_8 FILLER_7_1330 ();
 sg13g2_decap_8 FILLER_7_1337 ();
 sg13g2_decap_8 FILLER_7_1344 ();
 sg13g2_decap_8 FILLER_7_1351 ();
 sg13g2_decap_8 FILLER_7_1358 ();
 sg13g2_decap_8 FILLER_7_1365 ();
 sg13g2_decap_8 FILLER_7_1372 ();
 sg13g2_decap_8 FILLER_7_1379 ();
 sg13g2_decap_8 FILLER_7_1386 ();
 sg13g2_decap_8 FILLER_7_1393 ();
 sg13g2_decap_8 FILLER_7_1400 ();
 sg13g2_decap_8 FILLER_7_1407 ();
 sg13g2_decap_8 FILLER_7_1414 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_decap_8 FILLER_7_1428 ();
 sg13g2_decap_8 FILLER_7_1435 ();
 sg13g2_decap_8 FILLER_7_1442 ();
 sg13g2_decap_8 FILLER_7_1449 ();
 sg13g2_decap_8 FILLER_7_1456 ();
 sg13g2_decap_8 FILLER_7_1463 ();
 sg13g2_decap_8 FILLER_7_1470 ();
 sg13g2_decap_8 FILLER_7_1477 ();
 sg13g2_decap_8 FILLER_7_1484 ();
 sg13g2_decap_8 FILLER_7_1491 ();
 sg13g2_decap_8 FILLER_7_1498 ();
 sg13g2_decap_8 FILLER_7_1505 ();
 sg13g2_decap_8 FILLER_7_1512 ();
 sg13g2_decap_8 FILLER_7_1519 ();
 sg13g2_decap_8 FILLER_7_1526 ();
 sg13g2_decap_8 FILLER_7_1533 ();
 sg13g2_decap_8 FILLER_7_1540 ();
 sg13g2_decap_8 FILLER_7_1547 ();
 sg13g2_decap_8 FILLER_7_1554 ();
 sg13g2_decap_8 FILLER_7_1561 ();
 sg13g2_decap_8 FILLER_7_1568 ();
 sg13g2_decap_8 FILLER_7_1575 ();
 sg13g2_decap_8 FILLER_7_1582 ();
 sg13g2_decap_8 FILLER_7_1589 ();
 sg13g2_decap_8 FILLER_7_1596 ();
 sg13g2_decap_8 FILLER_7_1603 ();
 sg13g2_decap_8 FILLER_7_1610 ();
 sg13g2_decap_8 FILLER_7_1617 ();
 sg13g2_decap_8 FILLER_7_1624 ();
 sg13g2_decap_8 FILLER_7_1631 ();
 sg13g2_decap_8 FILLER_7_1638 ();
 sg13g2_decap_8 FILLER_7_1645 ();
 sg13g2_decap_8 FILLER_7_1652 ();
 sg13g2_decap_8 FILLER_7_1659 ();
 sg13g2_decap_8 FILLER_7_1666 ();
 sg13g2_decap_8 FILLER_7_1673 ();
 sg13g2_decap_8 FILLER_7_1680 ();
 sg13g2_decap_8 FILLER_7_1687 ();
 sg13g2_decap_8 FILLER_7_1694 ();
 sg13g2_decap_8 FILLER_7_1701 ();
 sg13g2_decap_8 FILLER_7_1708 ();
 sg13g2_decap_8 FILLER_7_1715 ();
 sg13g2_decap_8 FILLER_7_1722 ();
 sg13g2_decap_8 FILLER_7_1729 ();
 sg13g2_decap_8 FILLER_7_1736 ();
 sg13g2_decap_8 FILLER_7_1743 ();
 sg13g2_decap_8 FILLER_7_1750 ();
 sg13g2_decap_8 FILLER_7_1757 ();
 sg13g2_decap_4 FILLER_7_1764 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_decap_8 FILLER_8_1029 ();
 sg13g2_decap_8 FILLER_8_1036 ();
 sg13g2_decap_8 FILLER_8_1043 ();
 sg13g2_decap_8 FILLER_8_1050 ();
 sg13g2_decap_8 FILLER_8_1057 ();
 sg13g2_decap_8 FILLER_8_1064 ();
 sg13g2_decap_8 FILLER_8_1071 ();
 sg13g2_decap_8 FILLER_8_1078 ();
 sg13g2_decap_8 FILLER_8_1085 ();
 sg13g2_decap_8 FILLER_8_1092 ();
 sg13g2_decap_8 FILLER_8_1099 ();
 sg13g2_decap_8 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1113 ();
 sg13g2_decap_8 FILLER_8_1120 ();
 sg13g2_decap_8 FILLER_8_1127 ();
 sg13g2_decap_8 FILLER_8_1134 ();
 sg13g2_decap_8 FILLER_8_1141 ();
 sg13g2_decap_8 FILLER_8_1148 ();
 sg13g2_decap_8 FILLER_8_1155 ();
 sg13g2_decap_8 FILLER_8_1162 ();
 sg13g2_decap_8 FILLER_8_1169 ();
 sg13g2_decap_8 FILLER_8_1176 ();
 sg13g2_decap_8 FILLER_8_1183 ();
 sg13g2_decap_8 FILLER_8_1190 ();
 sg13g2_decap_8 FILLER_8_1197 ();
 sg13g2_decap_8 FILLER_8_1204 ();
 sg13g2_decap_8 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1218 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_8 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_decap_8 FILLER_8_1253 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_decap_8 FILLER_8_1267 ();
 sg13g2_decap_8 FILLER_8_1274 ();
 sg13g2_decap_8 FILLER_8_1281 ();
 sg13g2_decap_8 FILLER_8_1288 ();
 sg13g2_decap_8 FILLER_8_1295 ();
 sg13g2_decap_8 FILLER_8_1302 ();
 sg13g2_decap_8 FILLER_8_1309 ();
 sg13g2_decap_8 FILLER_8_1316 ();
 sg13g2_decap_8 FILLER_8_1323 ();
 sg13g2_decap_8 FILLER_8_1330 ();
 sg13g2_decap_8 FILLER_8_1337 ();
 sg13g2_decap_8 FILLER_8_1344 ();
 sg13g2_decap_8 FILLER_8_1351 ();
 sg13g2_decap_8 FILLER_8_1358 ();
 sg13g2_decap_8 FILLER_8_1365 ();
 sg13g2_decap_8 FILLER_8_1372 ();
 sg13g2_decap_8 FILLER_8_1379 ();
 sg13g2_decap_8 FILLER_8_1386 ();
 sg13g2_decap_8 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1400 ();
 sg13g2_decap_8 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1414 ();
 sg13g2_decap_8 FILLER_8_1421 ();
 sg13g2_decap_8 FILLER_8_1428 ();
 sg13g2_decap_8 FILLER_8_1435 ();
 sg13g2_decap_8 FILLER_8_1442 ();
 sg13g2_decap_8 FILLER_8_1449 ();
 sg13g2_decap_8 FILLER_8_1456 ();
 sg13g2_decap_8 FILLER_8_1463 ();
 sg13g2_decap_8 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1477 ();
 sg13g2_decap_8 FILLER_8_1484 ();
 sg13g2_decap_8 FILLER_8_1491 ();
 sg13g2_decap_8 FILLER_8_1498 ();
 sg13g2_decap_8 FILLER_8_1505 ();
 sg13g2_decap_8 FILLER_8_1512 ();
 sg13g2_decap_8 FILLER_8_1519 ();
 sg13g2_decap_8 FILLER_8_1526 ();
 sg13g2_decap_8 FILLER_8_1533 ();
 sg13g2_decap_8 FILLER_8_1540 ();
 sg13g2_decap_8 FILLER_8_1547 ();
 sg13g2_decap_8 FILLER_8_1554 ();
 sg13g2_decap_8 FILLER_8_1561 ();
 sg13g2_decap_8 FILLER_8_1568 ();
 sg13g2_decap_8 FILLER_8_1575 ();
 sg13g2_decap_8 FILLER_8_1582 ();
 sg13g2_decap_8 FILLER_8_1589 ();
 sg13g2_decap_8 FILLER_8_1596 ();
 sg13g2_decap_8 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1610 ();
 sg13g2_decap_8 FILLER_8_1617 ();
 sg13g2_decap_8 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1638 ();
 sg13g2_decap_8 FILLER_8_1645 ();
 sg13g2_decap_8 FILLER_8_1652 ();
 sg13g2_decap_8 FILLER_8_1659 ();
 sg13g2_decap_8 FILLER_8_1666 ();
 sg13g2_decap_8 FILLER_8_1673 ();
 sg13g2_decap_8 FILLER_8_1680 ();
 sg13g2_decap_8 FILLER_8_1687 ();
 sg13g2_decap_8 FILLER_8_1694 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_8 FILLER_8_1757 ();
 sg13g2_decap_4 FILLER_8_1764 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_9_1029 ();
 sg13g2_decap_8 FILLER_9_1036 ();
 sg13g2_decap_8 FILLER_9_1043 ();
 sg13g2_decap_8 FILLER_9_1050 ();
 sg13g2_decap_8 FILLER_9_1057 ();
 sg13g2_decap_8 FILLER_9_1064 ();
 sg13g2_decap_8 FILLER_9_1071 ();
 sg13g2_decap_8 FILLER_9_1078 ();
 sg13g2_decap_8 FILLER_9_1085 ();
 sg13g2_decap_8 FILLER_9_1092 ();
 sg13g2_decap_8 FILLER_9_1099 ();
 sg13g2_decap_8 FILLER_9_1106 ();
 sg13g2_decap_8 FILLER_9_1113 ();
 sg13g2_decap_8 FILLER_9_1120 ();
 sg13g2_decap_8 FILLER_9_1127 ();
 sg13g2_decap_8 FILLER_9_1134 ();
 sg13g2_decap_8 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_decap_8 FILLER_9_1155 ();
 sg13g2_decap_8 FILLER_9_1162 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_8 FILLER_9_1183 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_decap_8 FILLER_9_1197 ();
 sg13g2_decap_8 FILLER_9_1204 ();
 sg13g2_decap_8 FILLER_9_1211 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1239 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_decap_8 FILLER_9_1260 ();
 sg13g2_decap_8 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_decap_8 FILLER_9_1323 ();
 sg13g2_decap_8 FILLER_9_1330 ();
 sg13g2_decap_8 FILLER_9_1337 ();
 sg13g2_decap_8 FILLER_9_1344 ();
 sg13g2_decap_8 FILLER_9_1351 ();
 sg13g2_decap_8 FILLER_9_1358 ();
 sg13g2_decap_8 FILLER_9_1365 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_decap_8 FILLER_9_1393 ();
 sg13g2_decap_8 FILLER_9_1400 ();
 sg13g2_decap_8 FILLER_9_1407 ();
 sg13g2_decap_8 FILLER_9_1414 ();
 sg13g2_decap_8 FILLER_9_1421 ();
 sg13g2_decap_8 FILLER_9_1428 ();
 sg13g2_decap_8 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1442 ();
 sg13g2_decap_8 FILLER_9_1449 ();
 sg13g2_decap_8 FILLER_9_1456 ();
 sg13g2_decap_8 FILLER_9_1463 ();
 sg13g2_decap_8 FILLER_9_1470 ();
 sg13g2_decap_8 FILLER_9_1477 ();
 sg13g2_decap_8 FILLER_9_1484 ();
 sg13g2_decap_8 FILLER_9_1491 ();
 sg13g2_decap_8 FILLER_9_1498 ();
 sg13g2_decap_8 FILLER_9_1505 ();
 sg13g2_decap_8 FILLER_9_1512 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1533 ();
 sg13g2_decap_8 FILLER_9_1540 ();
 sg13g2_decap_8 FILLER_9_1547 ();
 sg13g2_decap_8 FILLER_9_1554 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1575 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1603 ();
 sg13g2_decap_8 FILLER_9_1610 ();
 sg13g2_decap_8 FILLER_9_1617 ();
 sg13g2_decap_8 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1631 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_decap_8 FILLER_9_1645 ();
 sg13g2_decap_8 FILLER_9_1652 ();
 sg13g2_decap_8 FILLER_9_1659 ();
 sg13g2_decap_8 FILLER_9_1666 ();
 sg13g2_decap_8 FILLER_9_1673 ();
 sg13g2_decap_8 FILLER_9_1680 ();
 sg13g2_decap_8 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1701 ();
 sg13g2_decap_8 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1715 ();
 sg13g2_decap_8 FILLER_9_1722 ();
 sg13g2_decap_8 FILLER_9_1729 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_decap_8 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_decap_8 FILLER_9_1757 ();
 sg13g2_decap_4 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_decap_8 FILLER_10_875 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_decap_8 FILLER_10_903 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_decap_8 FILLER_10_938 ();
 sg13g2_decap_8 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_8 FILLER_10_1008 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_decap_8 FILLER_10_1022 ();
 sg13g2_decap_8 FILLER_10_1029 ();
 sg13g2_decap_8 FILLER_10_1036 ();
 sg13g2_decap_8 FILLER_10_1043 ();
 sg13g2_decap_8 FILLER_10_1050 ();
 sg13g2_decap_8 FILLER_10_1057 ();
 sg13g2_decap_8 FILLER_10_1064 ();
 sg13g2_decap_8 FILLER_10_1071 ();
 sg13g2_decap_8 FILLER_10_1078 ();
 sg13g2_decap_8 FILLER_10_1085 ();
 sg13g2_decap_8 FILLER_10_1092 ();
 sg13g2_decap_8 FILLER_10_1099 ();
 sg13g2_decap_8 FILLER_10_1106 ();
 sg13g2_decap_8 FILLER_10_1113 ();
 sg13g2_decap_8 FILLER_10_1120 ();
 sg13g2_decap_8 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1134 ();
 sg13g2_decap_8 FILLER_10_1141 ();
 sg13g2_decap_8 FILLER_10_1148 ();
 sg13g2_decap_8 FILLER_10_1155 ();
 sg13g2_decap_8 FILLER_10_1162 ();
 sg13g2_decap_8 FILLER_10_1169 ();
 sg13g2_decap_8 FILLER_10_1176 ();
 sg13g2_decap_8 FILLER_10_1183 ();
 sg13g2_decap_8 FILLER_10_1190 ();
 sg13g2_decap_8 FILLER_10_1197 ();
 sg13g2_decap_8 FILLER_10_1204 ();
 sg13g2_decap_8 FILLER_10_1211 ();
 sg13g2_decap_8 FILLER_10_1218 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1246 ();
 sg13g2_decap_8 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1260 ();
 sg13g2_decap_8 FILLER_10_1267 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_8 FILLER_10_1281 ();
 sg13g2_decap_8 FILLER_10_1288 ();
 sg13g2_decap_8 FILLER_10_1295 ();
 sg13g2_decap_8 FILLER_10_1302 ();
 sg13g2_decap_8 FILLER_10_1309 ();
 sg13g2_decap_8 FILLER_10_1316 ();
 sg13g2_decap_8 FILLER_10_1323 ();
 sg13g2_decap_8 FILLER_10_1330 ();
 sg13g2_decap_8 FILLER_10_1337 ();
 sg13g2_decap_8 FILLER_10_1344 ();
 sg13g2_decap_8 FILLER_10_1351 ();
 sg13g2_decap_8 FILLER_10_1358 ();
 sg13g2_decap_8 FILLER_10_1365 ();
 sg13g2_decap_8 FILLER_10_1372 ();
 sg13g2_decap_8 FILLER_10_1379 ();
 sg13g2_decap_8 FILLER_10_1386 ();
 sg13g2_decap_8 FILLER_10_1393 ();
 sg13g2_decap_8 FILLER_10_1400 ();
 sg13g2_decap_8 FILLER_10_1407 ();
 sg13g2_decap_8 FILLER_10_1414 ();
 sg13g2_decap_8 FILLER_10_1421 ();
 sg13g2_decap_8 FILLER_10_1428 ();
 sg13g2_decap_8 FILLER_10_1435 ();
 sg13g2_decap_8 FILLER_10_1442 ();
 sg13g2_decap_8 FILLER_10_1449 ();
 sg13g2_decap_8 FILLER_10_1456 ();
 sg13g2_decap_8 FILLER_10_1463 ();
 sg13g2_decap_8 FILLER_10_1470 ();
 sg13g2_decap_8 FILLER_10_1477 ();
 sg13g2_decap_8 FILLER_10_1484 ();
 sg13g2_decap_8 FILLER_10_1491 ();
 sg13g2_decap_8 FILLER_10_1498 ();
 sg13g2_decap_8 FILLER_10_1505 ();
 sg13g2_decap_8 FILLER_10_1512 ();
 sg13g2_decap_8 FILLER_10_1519 ();
 sg13g2_decap_8 FILLER_10_1526 ();
 sg13g2_decap_8 FILLER_10_1533 ();
 sg13g2_decap_8 FILLER_10_1540 ();
 sg13g2_decap_8 FILLER_10_1547 ();
 sg13g2_decap_8 FILLER_10_1554 ();
 sg13g2_decap_8 FILLER_10_1561 ();
 sg13g2_decap_8 FILLER_10_1568 ();
 sg13g2_decap_8 FILLER_10_1575 ();
 sg13g2_decap_8 FILLER_10_1582 ();
 sg13g2_decap_8 FILLER_10_1589 ();
 sg13g2_decap_8 FILLER_10_1596 ();
 sg13g2_decap_8 FILLER_10_1603 ();
 sg13g2_decap_8 FILLER_10_1610 ();
 sg13g2_decap_8 FILLER_10_1617 ();
 sg13g2_decap_8 FILLER_10_1624 ();
 sg13g2_decap_8 FILLER_10_1631 ();
 sg13g2_decap_8 FILLER_10_1638 ();
 sg13g2_decap_8 FILLER_10_1645 ();
 sg13g2_decap_8 FILLER_10_1652 ();
 sg13g2_decap_8 FILLER_10_1659 ();
 sg13g2_decap_8 FILLER_10_1666 ();
 sg13g2_decap_8 FILLER_10_1673 ();
 sg13g2_decap_8 FILLER_10_1680 ();
 sg13g2_decap_8 FILLER_10_1687 ();
 sg13g2_decap_8 FILLER_10_1694 ();
 sg13g2_decap_8 FILLER_10_1701 ();
 sg13g2_decap_8 FILLER_10_1708 ();
 sg13g2_decap_8 FILLER_10_1715 ();
 sg13g2_decap_8 FILLER_10_1722 ();
 sg13g2_decap_8 FILLER_10_1729 ();
 sg13g2_decap_8 FILLER_10_1736 ();
 sg13g2_decap_8 FILLER_10_1743 ();
 sg13g2_decap_8 FILLER_10_1750 ();
 sg13g2_decap_8 FILLER_10_1757 ();
 sg13g2_decap_4 FILLER_10_1764 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_8 FILLER_11_1029 ();
 sg13g2_decap_8 FILLER_11_1036 ();
 sg13g2_decap_8 FILLER_11_1043 ();
 sg13g2_decap_8 FILLER_11_1050 ();
 sg13g2_decap_8 FILLER_11_1057 ();
 sg13g2_decap_8 FILLER_11_1064 ();
 sg13g2_decap_8 FILLER_11_1071 ();
 sg13g2_decap_8 FILLER_11_1078 ();
 sg13g2_decap_8 FILLER_11_1085 ();
 sg13g2_decap_8 FILLER_11_1092 ();
 sg13g2_decap_8 FILLER_11_1099 ();
 sg13g2_decap_8 FILLER_11_1106 ();
 sg13g2_decap_8 FILLER_11_1113 ();
 sg13g2_decap_8 FILLER_11_1120 ();
 sg13g2_decap_8 FILLER_11_1127 ();
 sg13g2_decap_8 FILLER_11_1134 ();
 sg13g2_decap_8 FILLER_11_1141 ();
 sg13g2_decap_8 FILLER_11_1148 ();
 sg13g2_decap_8 FILLER_11_1155 ();
 sg13g2_decap_8 FILLER_11_1162 ();
 sg13g2_decap_8 FILLER_11_1169 ();
 sg13g2_decap_8 FILLER_11_1176 ();
 sg13g2_decap_8 FILLER_11_1183 ();
 sg13g2_decap_8 FILLER_11_1190 ();
 sg13g2_decap_8 FILLER_11_1197 ();
 sg13g2_decap_8 FILLER_11_1204 ();
 sg13g2_decap_8 FILLER_11_1211 ();
 sg13g2_decap_8 FILLER_11_1218 ();
 sg13g2_decap_8 FILLER_11_1225 ();
 sg13g2_decap_8 FILLER_11_1232 ();
 sg13g2_decap_8 FILLER_11_1239 ();
 sg13g2_decap_8 FILLER_11_1246 ();
 sg13g2_decap_8 FILLER_11_1253 ();
 sg13g2_decap_8 FILLER_11_1260 ();
 sg13g2_decap_8 FILLER_11_1267 ();
 sg13g2_decap_8 FILLER_11_1274 ();
 sg13g2_decap_8 FILLER_11_1281 ();
 sg13g2_decap_8 FILLER_11_1288 ();
 sg13g2_decap_8 FILLER_11_1295 ();
 sg13g2_decap_8 FILLER_11_1302 ();
 sg13g2_decap_8 FILLER_11_1309 ();
 sg13g2_decap_8 FILLER_11_1316 ();
 sg13g2_decap_8 FILLER_11_1323 ();
 sg13g2_decap_8 FILLER_11_1330 ();
 sg13g2_decap_8 FILLER_11_1337 ();
 sg13g2_decap_8 FILLER_11_1344 ();
 sg13g2_decap_8 FILLER_11_1351 ();
 sg13g2_decap_8 FILLER_11_1358 ();
 sg13g2_decap_8 FILLER_11_1365 ();
 sg13g2_decap_8 FILLER_11_1372 ();
 sg13g2_decap_8 FILLER_11_1379 ();
 sg13g2_decap_8 FILLER_11_1386 ();
 sg13g2_decap_8 FILLER_11_1393 ();
 sg13g2_decap_8 FILLER_11_1400 ();
 sg13g2_decap_8 FILLER_11_1407 ();
 sg13g2_decap_8 FILLER_11_1414 ();
 sg13g2_decap_8 FILLER_11_1421 ();
 sg13g2_decap_8 FILLER_11_1428 ();
 sg13g2_decap_8 FILLER_11_1435 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_8 FILLER_11_1449 ();
 sg13g2_decap_8 FILLER_11_1456 ();
 sg13g2_decap_8 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1470 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_8 FILLER_11_1484 ();
 sg13g2_decap_8 FILLER_11_1491 ();
 sg13g2_decap_8 FILLER_11_1498 ();
 sg13g2_decap_8 FILLER_11_1505 ();
 sg13g2_decap_8 FILLER_11_1512 ();
 sg13g2_decap_8 FILLER_11_1519 ();
 sg13g2_decap_8 FILLER_11_1526 ();
 sg13g2_decap_8 FILLER_11_1533 ();
 sg13g2_decap_8 FILLER_11_1540 ();
 sg13g2_decap_8 FILLER_11_1547 ();
 sg13g2_decap_8 FILLER_11_1554 ();
 sg13g2_decap_8 FILLER_11_1561 ();
 sg13g2_decap_8 FILLER_11_1568 ();
 sg13g2_decap_8 FILLER_11_1575 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_decap_8 FILLER_11_1589 ();
 sg13g2_decap_8 FILLER_11_1596 ();
 sg13g2_decap_8 FILLER_11_1603 ();
 sg13g2_decap_8 FILLER_11_1610 ();
 sg13g2_decap_8 FILLER_11_1617 ();
 sg13g2_decap_8 FILLER_11_1624 ();
 sg13g2_decap_8 FILLER_11_1631 ();
 sg13g2_decap_8 FILLER_11_1638 ();
 sg13g2_decap_8 FILLER_11_1645 ();
 sg13g2_decap_8 FILLER_11_1652 ();
 sg13g2_decap_8 FILLER_11_1659 ();
 sg13g2_decap_8 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1680 ();
 sg13g2_decap_8 FILLER_11_1687 ();
 sg13g2_decap_8 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_decap_8 FILLER_11_1708 ();
 sg13g2_decap_8 FILLER_11_1715 ();
 sg13g2_decap_8 FILLER_11_1722 ();
 sg13g2_decap_8 FILLER_11_1729 ();
 sg13g2_decap_8 FILLER_11_1736 ();
 sg13g2_decap_8 FILLER_11_1743 ();
 sg13g2_decap_8 FILLER_11_1750 ();
 sg13g2_decap_8 FILLER_11_1757 ();
 sg13g2_decap_4 FILLER_11_1764 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_decap_8 FILLER_12_875 ();
 sg13g2_decap_8 FILLER_12_882 ();
 sg13g2_decap_8 FILLER_12_889 ();
 sg13g2_decap_8 FILLER_12_896 ();
 sg13g2_decap_8 FILLER_12_903 ();
 sg13g2_decap_8 FILLER_12_910 ();
 sg13g2_decap_8 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_924 ();
 sg13g2_decap_8 FILLER_12_931 ();
 sg13g2_decap_8 FILLER_12_938 ();
 sg13g2_decap_8 FILLER_12_945 ();
 sg13g2_decap_8 FILLER_12_952 ();
 sg13g2_decap_8 FILLER_12_959 ();
 sg13g2_decap_8 FILLER_12_966 ();
 sg13g2_decap_8 FILLER_12_973 ();
 sg13g2_decap_8 FILLER_12_980 ();
 sg13g2_decap_8 FILLER_12_987 ();
 sg13g2_decap_8 FILLER_12_994 ();
 sg13g2_decap_8 FILLER_12_1001 ();
 sg13g2_decap_8 FILLER_12_1008 ();
 sg13g2_decap_8 FILLER_12_1015 ();
 sg13g2_decap_8 FILLER_12_1022 ();
 sg13g2_decap_8 FILLER_12_1029 ();
 sg13g2_decap_8 FILLER_12_1036 ();
 sg13g2_decap_8 FILLER_12_1043 ();
 sg13g2_decap_8 FILLER_12_1050 ();
 sg13g2_decap_8 FILLER_12_1057 ();
 sg13g2_decap_8 FILLER_12_1064 ();
 sg13g2_decap_8 FILLER_12_1071 ();
 sg13g2_decap_8 FILLER_12_1078 ();
 sg13g2_decap_8 FILLER_12_1085 ();
 sg13g2_decap_8 FILLER_12_1092 ();
 sg13g2_decap_8 FILLER_12_1099 ();
 sg13g2_decap_8 FILLER_12_1106 ();
 sg13g2_decap_8 FILLER_12_1113 ();
 sg13g2_decap_8 FILLER_12_1120 ();
 sg13g2_decap_8 FILLER_12_1127 ();
 sg13g2_decap_8 FILLER_12_1134 ();
 sg13g2_decap_8 FILLER_12_1141 ();
 sg13g2_decap_8 FILLER_12_1148 ();
 sg13g2_decap_8 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1169 ();
 sg13g2_decap_8 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1190 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_decap_8 FILLER_12_1204 ();
 sg13g2_decap_8 FILLER_12_1211 ();
 sg13g2_decap_8 FILLER_12_1218 ();
 sg13g2_decap_8 FILLER_12_1225 ();
 sg13g2_decap_8 FILLER_12_1232 ();
 sg13g2_decap_8 FILLER_12_1239 ();
 sg13g2_decap_8 FILLER_12_1246 ();
 sg13g2_decap_8 FILLER_12_1253 ();
 sg13g2_decap_8 FILLER_12_1260 ();
 sg13g2_decap_8 FILLER_12_1267 ();
 sg13g2_decap_8 FILLER_12_1274 ();
 sg13g2_decap_8 FILLER_12_1281 ();
 sg13g2_decap_8 FILLER_12_1288 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_8 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1316 ();
 sg13g2_decap_8 FILLER_12_1323 ();
 sg13g2_decap_8 FILLER_12_1330 ();
 sg13g2_decap_8 FILLER_12_1337 ();
 sg13g2_decap_8 FILLER_12_1344 ();
 sg13g2_decap_8 FILLER_12_1351 ();
 sg13g2_decap_8 FILLER_12_1358 ();
 sg13g2_decap_8 FILLER_12_1365 ();
 sg13g2_decap_8 FILLER_12_1372 ();
 sg13g2_decap_8 FILLER_12_1379 ();
 sg13g2_decap_8 FILLER_12_1386 ();
 sg13g2_decap_8 FILLER_12_1393 ();
 sg13g2_decap_8 FILLER_12_1400 ();
 sg13g2_decap_8 FILLER_12_1407 ();
 sg13g2_decap_8 FILLER_12_1414 ();
 sg13g2_decap_8 FILLER_12_1421 ();
 sg13g2_decap_8 FILLER_12_1428 ();
 sg13g2_decap_8 FILLER_12_1435 ();
 sg13g2_decap_8 FILLER_12_1442 ();
 sg13g2_decap_8 FILLER_12_1449 ();
 sg13g2_decap_8 FILLER_12_1456 ();
 sg13g2_decap_8 FILLER_12_1463 ();
 sg13g2_decap_8 FILLER_12_1470 ();
 sg13g2_decap_8 FILLER_12_1477 ();
 sg13g2_decap_8 FILLER_12_1484 ();
 sg13g2_decap_8 FILLER_12_1491 ();
 sg13g2_decap_8 FILLER_12_1498 ();
 sg13g2_decap_8 FILLER_12_1505 ();
 sg13g2_decap_8 FILLER_12_1512 ();
 sg13g2_decap_8 FILLER_12_1519 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_8 FILLER_12_1540 ();
 sg13g2_decap_8 FILLER_12_1547 ();
 sg13g2_decap_8 FILLER_12_1554 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_decap_8 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_8 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1617 ();
 sg13g2_decap_8 FILLER_12_1624 ();
 sg13g2_decap_8 FILLER_12_1631 ();
 sg13g2_decap_8 FILLER_12_1638 ();
 sg13g2_decap_8 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1652 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_8 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1673 ();
 sg13g2_decap_8 FILLER_12_1680 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_8 FILLER_12_1701 ();
 sg13g2_decap_8 FILLER_12_1708 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_8 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1750 ();
 sg13g2_decap_8 FILLER_12_1757 ();
 sg13g2_decap_4 FILLER_12_1764 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_decap_8 FILLER_13_875 ();
 sg13g2_decap_8 FILLER_13_882 ();
 sg13g2_decap_8 FILLER_13_889 ();
 sg13g2_decap_8 FILLER_13_896 ();
 sg13g2_decap_8 FILLER_13_903 ();
 sg13g2_decap_8 FILLER_13_910 ();
 sg13g2_decap_8 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_924 ();
 sg13g2_decap_8 FILLER_13_931 ();
 sg13g2_decap_8 FILLER_13_938 ();
 sg13g2_decap_8 FILLER_13_945 ();
 sg13g2_decap_8 FILLER_13_952 ();
 sg13g2_decap_8 FILLER_13_959 ();
 sg13g2_decap_8 FILLER_13_966 ();
 sg13g2_decap_8 FILLER_13_973 ();
 sg13g2_decap_8 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_decap_8 FILLER_13_1015 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_8 FILLER_13_1029 ();
 sg13g2_decap_8 FILLER_13_1036 ();
 sg13g2_decap_8 FILLER_13_1043 ();
 sg13g2_decap_8 FILLER_13_1050 ();
 sg13g2_decap_8 FILLER_13_1057 ();
 sg13g2_decap_8 FILLER_13_1064 ();
 sg13g2_decap_8 FILLER_13_1071 ();
 sg13g2_decap_8 FILLER_13_1078 ();
 sg13g2_decap_8 FILLER_13_1085 ();
 sg13g2_decap_8 FILLER_13_1092 ();
 sg13g2_decap_8 FILLER_13_1099 ();
 sg13g2_decap_8 FILLER_13_1106 ();
 sg13g2_decap_8 FILLER_13_1113 ();
 sg13g2_decap_8 FILLER_13_1120 ();
 sg13g2_decap_8 FILLER_13_1127 ();
 sg13g2_decap_8 FILLER_13_1134 ();
 sg13g2_decap_8 FILLER_13_1141 ();
 sg13g2_decap_8 FILLER_13_1148 ();
 sg13g2_decap_8 FILLER_13_1155 ();
 sg13g2_decap_8 FILLER_13_1162 ();
 sg13g2_decap_8 FILLER_13_1169 ();
 sg13g2_decap_8 FILLER_13_1176 ();
 sg13g2_decap_8 FILLER_13_1183 ();
 sg13g2_decap_8 FILLER_13_1190 ();
 sg13g2_decap_8 FILLER_13_1197 ();
 sg13g2_decap_8 FILLER_13_1204 ();
 sg13g2_decap_8 FILLER_13_1211 ();
 sg13g2_decap_8 FILLER_13_1218 ();
 sg13g2_decap_8 FILLER_13_1225 ();
 sg13g2_decap_8 FILLER_13_1232 ();
 sg13g2_decap_8 FILLER_13_1239 ();
 sg13g2_decap_8 FILLER_13_1246 ();
 sg13g2_decap_8 FILLER_13_1253 ();
 sg13g2_decap_8 FILLER_13_1260 ();
 sg13g2_decap_8 FILLER_13_1267 ();
 sg13g2_decap_8 FILLER_13_1274 ();
 sg13g2_decap_8 FILLER_13_1281 ();
 sg13g2_decap_8 FILLER_13_1288 ();
 sg13g2_decap_8 FILLER_13_1295 ();
 sg13g2_decap_8 FILLER_13_1302 ();
 sg13g2_decap_8 FILLER_13_1309 ();
 sg13g2_decap_8 FILLER_13_1316 ();
 sg13g2_decap_8 FILLER_13_1323 ();
 sg13g2_decap_8 FILLER_13_1330 ();
 sg13g2_decap_8 FILLER_13_1337 ();
 sg13g2_decap_8 FILLER_13_1344 ();
 sg13g2_decap_8 FILLER_13_1351 ();
 sg13g2_decap_8 FILLER_13_1358 ();
 sg13g2_decap_8 FILLER_13_1365 ();
 sg13g2_decap_8 FILLER_13_1372 ();
 sg13g2_decap_8 FILLER_13_1379 ();
 sg13g2_decap_8 FILLER_13_1386 ();
 sg13g2_decap_8 FILLER_13_1393 ();
 sg13g2_decap_8 FILLER_13_1400 ();
 sg13g2_decap_8 FILLER_13_1407 ();
 sg13g2_decap_8 FILLER_13_1414 ();
 sg13g2_decap_8 FILLER_13_1421 ();
 sg13g2_decap_8 FILLER_13_1428 ();
 sg13g2_decap_8 FILLER_13_1435 ();
 sg13g2_decap_8 FILLER_13_1442 ();
 sg13g2_decap_8 FILLER_13_1449 ();
 sg13g2_decap_8 FILLER_13_1456 ();
 sg13g2_decap_8 FILLER_13_1463 ();
 sg13g2_decap_8 FILLER_13_1470 ();
 sg13g2_decap_8 FILLER_13_1477 ();
 sg13g2_decap_8 FILLER_13_1484 ();
 sg13g2_decap_8 FILLER_13_1491 ();
 sg13g2_decap_8 FILLER_13_1498 ();
 sg13g2_decap_8 FILLER_13_1505 ();
 sg13g2_decap_8 FILLER_13_1512 ();
 sg13g2_decap_8 FILLER_13_1519 ();
 sg13g2_decap_8 FILLER_13_1526 ();
 sg13g2_decap_8 FILLER_13_1533 ();
 sg13g2_decap_8 FILLER_13_1540 ();
 sg13g2_decap_8 FILLER_13_1547 ();
 sg13g2_decap_8 FILLER_13_1554 ();
 sg13g2_decap_8 FILLER_13_1561 ();
 sg13g2_decap_8 FILLER_13_1568 ();
 sg13g2_decap_8 FILLER_13_1575 ();
 sg13g2_decap_8 FILLER_13_1582 ();
 sg13g2_decap_8 FILLER_13_1589 ();
 sg13g2_decap_8 FILLER_13_1596 ();
 sg13g2_decap_8 FILLER_13_1603 ();
 sg13g2_decap_8 FILLER_13_1610 ();
 sg13g2_decap_8 FILLER_13_1617 ();
 sg13g2_decap_8 FILLER_13_1624 ();
 sg13g2_decap_8 FILLER_13_1631 ();
 sg13g2_decap_8 FILLER_13_1638 ();
 sg13g2_decap_8 FILLER_13_1645 ();
 sg13g2_decap_8 FILLER_13_1652 ();
 sg13g2_decap_8 FILLER_13_1659 ();
 sg13g2_decap_8 FILLER_13_1666 ();
 sg13g2_decap_8 FILLER_13_1673 ();
 sg13g2_decap_8 FILLER_13_1680 ();
 sg13g2_decap_8 FILLER_13_1687 ();
 sg13g2_decap_8 FILLER_13_1694 ();
 sg13g2_decap_8 FILLER_13_1701 ();
 sg13g2_decap_8 FILLER_13_1708 ();
 sg13g2_decap_8 FILLER_13_1715 ();
 sg13g2_decap_8 FILLER_13_1722 ();
 sg13g2_decap_8 FILLER_13_1729 ();
 sg13g2_decap_8 FILLER_13_1736 ();
 sg13g2_decap_8 FILLER_13_1743 ();
 sg13g2_decap_8 FILLER_13_1750 ();
 sg13g2_decap_8 FILLER_13_1757 ();
 sg13g2_decap_4 FILLER_13_1764 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_14_868 ();
 sg13g2_decap_8 FILLER_14_875 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_8 FILLER_14_889 ();
 sg13g2_decap_8 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_8 FILLER_14_910 ();
 sg13g2_decap_8 FILLER_14_917 ();
 sg13g2_decap_8 FILLER_14_924 ();
 sg13g2_decap_8 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_decap_8 FILLER_14_945 ();
 sg13g2_decap_8 FILLER_14_952 ();
 sg13g2_decap_8 FILLER_14_959 ();
 sg13g2_decap_8 FILLER_14_966 ();
 sg13g2_decap_8 FILLER_14_973 ();
 sg13g2_decap_8 FILLER_14_980 ();
 sg13g2_decap_8 FILLER_14_987 ();
 sg13g2_decap_8 FILLER_14_994 ();
 sg13g2_decap_8 FILLER_14_1001 ();
 sg13g2_decap_8 FILLER_14_1008 ();
 sg13g2_decap_8 FILLER_14_1015 ();
 sg13g2_decap_8 FILLER_14_1022 ();
 sg13g2_decap_8 FILLER_14_1029 ();
 sg13g2_decap_8 FILLER_14_1036 ();
 sg13g2_decap_8 FILLER_14_1043 ();
 sg13g2_decap_8 FILLER_14_1050 ();
 sg13g2_decap_8 FILLER_14_1057 ();
 sg13g2_decap_8 FILLER_14_1064 ();
 sg13g2_decap_8 FILLER_14_1071 ();
 sg13g2_decap_8 FILLER_14_1078 ();
 sg13g2_decap_8 FILLER_14_1085 ();
 sg13g2_decap_8 FILLER_14_1092 ();
 sg13g2_decap_8 FILLER_14_1099 ();
 sg13g2_decap_8 FILLER_14_1106 ();
 sg13g2_decap_8 FILLER_14_1113 ();
 sg13g2_decap_8 FILLER_14_1120 ();
 sg13g2_decap_8 FILLER_14_1127 ();
 sg13g2_decap_8 FILLER_14_1134 ();
 sg13g2_decap_8 FILLER_14_1141 ();
 sg13g2_decap_8 FILLER_14_1148 ();
 sg13g2_decap_8 FILLER_14_1155 ();
 sg13g2_decap_8 FILLER_14_1162 ();
 sg13g2_decap_8 FILLER_14_1169 ();
 sg13g2_decap_8 FILLER_14_1176 ();
 sg13g2_decap_8 FILLER_14_1183 ();
 sg13g2_decap_8 FILLER_14_1190 ();
 sg13g2_decap_8 FILLER_14_1197 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_8 FILLER_14_1211 ();
 sg13g2_decap_8 FILLER_14_1218 ();
 sg13g2_decap_8 FILLER_14_1225 ();
 sg13g2_decap_8 FILLER_14_1232 ();
 sg13g2_decap_8 FILLER_14_1239 ();
 sg13g2_decap_8 FILLER_14_1246 ();
 sg13g2_decap_8 FILLER_14_1253 ();
 sg13g2_decap_8 FILLER_14_1260 ();
 sg13g2_decap_8 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_decap_8 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_decap_8 FILLER_14_1323 ();
 sg13g2_decap_8 FILLER_14_1330 ();
 sg13g2_decap_8 FILLER_14_1337 ();
 sg13g2_decap_8 FILLER_14_1344 ();
 sg13g2_decap_8 FILLER_14_1351 ();
 sg13g2_decap_8 FILLER_14_1358 ();
 sg13g2_decap_8 FILLER_14_1365 ();
 sg13g2_decap_8 FILLER_14_1372 ();
 sg13g2_decap_8 FILLER_14_1379 ();
 sg13g2_decap_8 FILLER_14_1386 ();
 sg13g2_decap_8 FILLER_14_1393 ();
 sg13g2_decap_8 FILLER_14_1400 ();
 sg13g2_decap_8 FILLER_14_1407 ();
 sg13g2_decap_8 FILLER_14_1414 ();
 sg13g2_decap_8 FILLER_14_1421 ();
 sg13g2_decap_8 FILLER_14_1428 ();
 sg13g2_decap_8 FILLER_14_1435 ();
 sg13g2_decap_8 FILLER_14_1442 ();
 sg13g2_decap_8 FILLER_14_1449 ();
 sg13g2_decap_8 FILLER_14_1456 ();
 sg13g2_decap_8 FILLER_14_1463 ();
 sg13g2_decap_8 FILLER_14_1470 ();
 sg13g2_decap_8 FILLER_14_1477 ();
 sg13g2_decap_8 FILLER_14_1484 ();
 sg13g2_decap_8 FILLER_14_1491 ();
 sg13g2_decap_8 FILLER_14_1498 ();
 sg13g2_decap_8 FILLER_14_1505 ();
 sg13g2_decap_8 FILLER_14_1512 ();
 sg13g2_decap_8 FILLER_14_1519 ();
 sg13g2_decap_8 FILLER_14_1526 ();
 sg13g2_decap_8 FILLER_14_1533 ();
 sg13g2_decap_8 FILLER_14_1540 ();
 sg13g2_decap_8 FILLER_14_1547 ();
 sg13g2_decap_8 FILLER_14_1554 ();
 sg13g2_decap_8 FILLER_14_1561 ();
 sg13g2_decap_8 FILLER_14_1568 ();
 sg13g2_decap_8 FILLER_14_1575 ();
 sg13g2_decap_8 FILLER_14_1582 ();
 sg13g2_decap_8 FILLER_14_1589 ();
 sg13g2_decap_8 FILLER_14_1596 ();
 sg13g2_decap_8 FILLER_14_1603 ();
 sg13g2_decap_8 FILLER_14_1610 ();
 sg13g2_decap_8 FILLER_14_1617 ();
 sg13g2_decap_8 FILLER_14_1624 ();
 sg13g2_decap_8 FILLER_14_1631 ();
 sg13g2_decap_8 FILLER_14_1638 ();
 sg13g2_decap_8 FILLER_14_1645 ();
 sg13g2_decap_8 FILLER_14_1652 ();
 sg13g2_decap_8 FILLER_14_1659 ();
 sg13g2_decap_8 FILLER_14_1666 ();
 sg13g2_decap_8 FILLER_14_1673 ();
 sg13g2_decap_8 FILLER_14_1680 ();
 sg13g2_decap_8 FILLER_14_1687 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_decap_8 FILLER_14_1701 ();
 sg13g2_decap_8 FILLER_14_1708 ();
 sg13g2_decap_8 FILLER_14_1715 ();
 sg13g2_decap_8 FILLER_14_1722 ();
 sg13g2_decap_8 FILLER_14_1729 ();
 sg13g2_decap_8 FILLER_14_1736 ();
 sg13g2_decap_8 FILLER_14_1743 ();
 sg13g2_decap_8 FILLER_14_1750 ();
 sg13g2_decap_8 FILLER_14_1757 ();
 sg13g2_decap_4 FILLER_14_1764 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_875 ();
 sg13g2_decap_8 FILLER_15_882 ();
 sg13g2_decap_8 FILLER_15_889 ();
 sg13g2_decap_8 FILLER_15_896 ();
 sg13g2_decap_8 FILLER_15_903 ();
 sg13g2_decap_8 FILLER_15_910 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_decap_8 FILLER_15_924 ();
 sg13g2_decap_8 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_938 ();
 sg13g2_decap_8 FILLER_15_945 ();
 sg13g2_decap_8 FILLER_15_952 ();
 sg13g2_decap_8 FILLER_15_959 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_decap_8 FILLER_15_973 ();
 sg13g2_decap_8 FILLER_15_980 ();
 sg13g2_decap_8 FILLER_15_987 ();
 sg13g2_decap_8 FILLER_15_994 ();
 sg13g2_decap_8 FILLER_15_1001 ();
 sg13g2_decap_8 FILLER_15_1008 ();
 sg13g2_decap_8 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1022 ();
 sg13g2_decap_8 FILLER_15_1029 ();
 sg13g2_decap_8 FILLER_15_1036 ();
 sg13g2_decap_8 FILLER_15_1043 ();
 sg13g2_decap_8 FILLER_15_1050 ();
 sg13g2_decap_8 FILLER_15_1057 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_decap_8 FILLER_15_1071 ();
 sg13g2_decap_8 FILLER_15_1078 ();
 sg13g2_decap_8 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1092 ();
 sg13g2_decap_8 FILLER_15_1099 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_decap_8 FILLER_15_1141 ();
 sg13g2_decap_8 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1155 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1197 ();
 sg13g2_decap_8 FILLER_15_1204 ();
 sg13g2_decap_8 FILLER_15_1211 ();
 sg13g2_decap_8 FILLER_15_1218 ();
 sg13g2_decap_8 FILLER_15_1225 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_decap_8 FILLER_15_1239 ();
 sg13g2_decap_8 FILLER_15_1246 ();
 sg13g2_decap_8 FILLER_15_1253 ();
 sg13g2_decap_8 FILLER_15_1260 ();
 sg13g2_decap_8 FILLER_15_1267 ();
 sg13g2_decap_8 FILLER_15_1274 ();
 sg13g2_decap_8 FILLER_15_1281 ();
 sg13g2_decap_8 FILLER_15_1288 ();
 sg13g2_decap_8 FILLER_15_1295 ();
 sg13g2_decap_8 FILLER_15_1302 ();
 sg13g2_decap_8 FILLER_15_1309 ();
 sg13g2_decap_8 FILLER_15_1316 ();
 sg13g2_decap_8 FILLER_15_1323 ();
 sg13g2_decap_8 FILLER_15_1330 ();
 sg13g2_decap_8 FILLER_15_1337 ();
 sg13g2_decap_8 FILLER_15_1344 ();
 sg13g2_decap_8 FILLER_15_1351 ();
 sg13g2_decap_8 FILLER_15_1358 ();
 sg13g2_decap_8 FILLER_15_1365 ();
 sg13g2_decap_8 FILLER_15_1372 ();
 sg13g2_decap_8 FILLER_15_1379 ();
 sg13g2_decap_8 FILLER_15_1386 ();
 sg13g2_decap_8 FILLER_15_1393 ();
 sg13g2_decap_8 FILLER_15_1400 ();
 sg13g2_decap_8 FILLER_15_1407 ();
 sg13g2_decap_8 FILLER_15_1414 ();
 sg13g2_decap_8 FILLER_15_1421 ();
 sg13g2_decap_8 FILLER_15_1428 ();
 sg13g2_decap_8 FILLER_15_1435 ();
 sg13g2_decap_8 FILLER_15_1442 ();
 sg13g2_decap_8 FILLER_15_1449 ();
 sg13g2_decap_8 FILLER_15_1456 ();
 sg13g2_decap_8 FILLER_15_1463 ();
 sg13g2_decap_8 FILLER_15_1470 ();
 sg13g2_decap_8 FILLER_15_1477 ();
 sg13g2_decap_8 FILLER_15_1484 ();
 sg13g2_decap_8 FILLER_15_1491 ();
 sg13g2_decap_8 FILLER_15_1498 ();
 sg13g2_decap_8 FILLER_15_1505 ();
 sg13g2_decap_8 FILLER_15_1512 ();
 sg13g2_decap_8 FILLER_15_1519 ();
 sg13g2_decap_8 FILLER_15_1526 ();
 sg13g2_decap_8 FILLER_15_1533 ();
 sg13g2_decap_8 FILLER_15_1540 ();
 sg13g2_decap_8 FILLER_15_1547 ();
 sg13g2_decap_8 FILLER_15_1554 ();
 sg13g2_decap_8 FILLER_15_1561 ();
 sg13g2_decap_8 FILLER_15_1568 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_decap_8 FILLER_15_1582 ();
 sg13g2_decap_8 FILLER_15_1589 ();
 sg13g2_decap_8 FILLER_15_1596 ();
 sg13g2_decap_8 FILLER_15_1603 ();
 sg13g2_decap_8 FILLER_15_1610 ();
 sg13g2_decap_8 FILLER_15_1617 ();
 sg13g2_decap_8 FILLER_15_1624 ();
 sg13g2_decap_8 FILLER_15_1631 ();
 sg13g2_decap_8 FILLER_15_1638 ();
 sg13g2_decap_8 FILLER_15_1645 ();
 sg13g2_decap_8 FILLER_15_1652 ();
 sg13g2_decap_8 FILLER_15_1659 ();
 sg13g2_decap_8 FILLER_15_1666 ();
 sg13g2_decap_8 FILLER_15_1673 ();
 sg13g2_decap_8 FILLER_15_1680 ();
 sg13g2_decap_8 FILLER_15_1687 ();
 sg13g2_decap_8 FILLER_15_1694 ();
 sg13g2_decap_8 FILLER_15_1701 ();
 sg13g2_decap_8 FILLER_15_1708 ();
 sg13g2_decap_8 FILLER_15_1715 ();
 sg13g2_decap_8 FILLER_15_1722 ();
 sg13g2_decap_8 FILLER_15_1729 ();
 sg13g2_decap_8 FILLER_15_1736 ();
 sg13g2_decap_8 FILLER_15_1743 ();
 sg13g2_decap_8 FILLER_15_1750 ();
 sg13g2_decap_8 FILLER_15_1757 ();
 sg13g2_decap_4 FILLER_15_1764 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_882 ();
 sg13g2_decap_8 FILLER_16_889 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_decap_8 FILLER_16_1029 ();
 sg13g2_decap_8 FILLER_16_1036 ();
 sg13g2_decap_8 FILLER_16_1043 ();
 sg13g2_decap_8 FILLER_16_1050 ();
 sg13g2_decap_8 FILLER_16_1057 ();
 sg13g2_decap_8 FILLER_16_1064 ();
 sg13g2_decap_8 FILLER_16_1071 ();
 sg13g2_decap_8 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1085 ();
 sg13g2_decap_8 FILLER_16_1092 ();
 sg13g2_decap_8 FILLER_16_1099 ();
 sg13g2_decap_8 FILLER_16_1106 ();
 sg13g2_decap_8 FILLER_16_1113 ();
 sg13g2_decap_8 FILLER_16_1120 ();
 sg13g2_decap_8 FILLER_16_1127 ();
 sg13g2_decap_8 FILLER_16_1134 ();
 sg13g2_decap_8 FILLER_16_1141 ();
 sg13g2_decap_8 FILLER_16_1148 ();
 sg13g2_decap_8 FILLER_16_1155 ();
 sg13g2_decap_8 FILLER_16_1162 ();
 sg13g2_decap_8 FILLER_16_1169 ();
 sg13g2_decap_8 FILLER_16_1176 ();
 sg13g2_decap_8 FILLER_16_1183 ();
 sg13g2_decap_8 FILLER_16_1190 ();
 sg13g2_decap_8 FILLER_16_1197 ();
 sg13g2_decap_8 FILLER_16_1204 ();
 sg13g2_decap_8 FILLER_16_1211 ();
 sg13g2_decap_8 FILLER_16_1218 ();
 sg13g2_decap_8 FILLER_16_1225 ();
 sg13g2_decap_8 FILLER_16_1232 ();
 sg13g2_decap_8 FILLER_16_1239 ();
 sg13g2_decap_8 FILLER_16_1246 ();
 sg13g2_decap_8 FILLER_16_1253 ();
 sg13g2_decap_8 FILLER_16_1260 ();
 sg13g2_decap_8 FILLER_16_1267 ();
 sg13g2_decap_8 FILLER_16_1274 ();
 sg13g2_decap_8 FILLER_16_1281 ();
 sg13g2_decap_8 FILLER_16_1288 ();
 sg13g2_decap_8 FILLER_16_1295 ();
 sg13g2_decap_8 FILLER_16_1302 ();
 sg13g2_decap_8 FILLER_16_1309 ();
 sg13g2_decap_8 FILLER_16_1316 ();
 sg13g2_decap_8 FILLER_16_1323 ();
 sg13g2_decap_8 FILLER_16_1330 ();
 sg13g2_decap_8 FILLER_16_1337 ();
 sg13g2_decap_8 FILLER_16_1344 ();
 sg13g2_decap_8 FILLER_16_1351 ();
 sg13g2_decap_8 FILLER_16_1358 ();
 sg13g2_decap_8 FILLER_16_1365 ();
 sg13g2_decap_8 FILLER_16_1372 ();
 sg13g2_decap_8 FILLER_16_1379 ();
 sg13g2_decap_8 FILLER_16_1386 ();
 sg13g2_decap_8 FILLER_16_1393 ();
 sg13g2_decap_8 FILLER_16_1400 ();
 sg13g2_decap_8 FILLER_16_1407 ();
 sg13g2_decap_8 FILLER_16_1414 ();
 sg13g2_decap_8 FILLER_16_1421 ();
 sg13g2_decap_8 FILLER_16_1428 ();
 sg13g2_decap_8 FILLER_16_1435 ();
 sg13g2_decap_8 FILLER_16_1442 ();
 sg13g2_decap_8 FILLER_16_1449 ();
 sg13g2_decap_8 FILLER_16_1456 ();
 sg13g2_decap_8 FILLER_16_1463 ();
 sg13g2_decap_8 FILLER_16_1470 ();
 sg13g2_decap_8 FILLER_16_1477 ();
 sg13g2_decap_8 FILLER_16_1484 ();
 sg13g2_decap_8 FILLER_16_1491 ();
 sg13g2_decap_8 FILLER_16_1498 ();
 sg13g2_decap_8 FILLER_16_1505 ();
 sg13g2_decap_8 FILLER_16_1512 ();
 sg13g2_decap_8 FILLER_16_1519 ();
 sg13g2_decap_8 FILLER_16_1526 ();
 sg13g2_decap_8 FILLER_16_1533 ();
 sg13g2_decap_8 FILLER_16_1540 ();
 sg13g2_decap_8 FILLER_16_1547 ();
 sg13g2_decap_8 FILLER_16_1554 ();
 sg13g2_decap_8 FILLER_16_1561 ();
 sg13g2_decap_8 FILLER_16_1568 ();
 sg13g2_decap_8 FILLER_16_1575 ();
 sg13g2_decap_8 FILLER_16_1582 ();
 sg13g2_decap_8 FILLER_16_1589 ();
 sg13g2_decap_8 FILLER_16_1596 ();
 sg13g2_decap_8 FILLER_16_1603 ();
 sg13g2_decap_8 FILLER_16_1610 ();
 sg13g2_decap_8 FILLER_16_1617 ();
 sg13g2_decap_8 FILLER_16_1624 ();
 sg13g2_decap_8 FILLER_16_1631 ();
 sg13g2_decap_8 FILLER_16_1638 ();
 sg13g2_decap_8 FILLER_16_1645 ();
 sg13g2_decap_8 FILLER_16_1652 ();
 sg13g2_decap_8 FILLER_16_1659 ();
 sg13g2_decap_8 FILLER_16_1666 ();
 sg13g2_decap_8 FILLER_16_1673 ();
 sg13g2_decap_8 FILLER_16_1680 ();
 sg13g2_decap_8 FILLER_16_1687 ();
 sg13g2_decap_8 FILLER_16_1694 ();
 sg13g2_decap_8 FILLER_16_1701 ();
 sg13g2_decap_8 FILLER_16_1708 ();
 sg13g2_decap_8 FILLER_16_1715 ();
 sg13g2_decap_8 FILLER_16_1722 ();
 sg13g2_decap_8 FILLER_16_1729 ();
 sg13g2_decap_8 FILLER_16_1736 ();
 sg13g2_decap_8 FILLER_16_1743 ();
 sg13g2_decap_8 FILLER_16_1750 ();
 sg13g2_decap_8 FILLER_16_1757 ();
 sg13g2_decap_4 FILLER_16_1764 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_decap_8 FILLER_17_1036 ();
 sg13g2_decap_8 FILLER_17_1043 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_decap_8 FILLER_17_1057 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_decap_8 FILLER_17_1071 ();
 sg13g2_decap_8 FILLER_17_1078 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_8 FILLER_17_1099 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_decap_8 FILLER_17_1323 ();
 sg13g2_decap_8 FILLER_17_1330 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_decap_8 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1358 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_decap_8 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1421 ();
 sg13g2_decap_8 FILLER_17_1428 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1442 ();
 sg13g2_decap_8 FILLER_17_1449 ();
 sg13g2_decap_8 FILLER_17_1456 ();
 sg13g2_decap_8 FILLER_17_1463 ();
 sg13g2_decap_8 FILLER_17_1470 ();
 sg13g2_decap_8 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1484 ();
 sg13g2_decap_8 FILLER_17_1491 ();
 sg13g2_decap_8 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1505 ();
 sg13g2_decap_8 FILLER_17_1512 ();
 sg13g2_decap_8 FILLER_17_1519 ();
 sg13g2_decap_8 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1540 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_decap_8 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_17_1631 ();
 sg13g2_decap_8 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1645 ();
 sg13g2_decap_8 FILLER_17_1652 ();
 sg13g2_decap_8 FILLER_17_1659 ();
 sg13g2_decap_8 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1673 ();
 sg13g2_decap_8 FILLER_17_1680 ();
 sg13g2_decap_8 FILLER_17_1687 ();
 sg13g2_decap_8 FILLER_17_1694 ();
 sg13g2_decap_8 FILLER_17_1701 ();
 sg13g2_decap_8 FILLER_17_1708 ();
 sg13g2_decap_8 FILLER_17_1715 ();
 sg13g2_decap_8 FILLER_17_1722 ();
 sg13g2_decap_8 FILLER_17_1729 ();
 sg13g2_decap_8 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1743 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_decap_4 FILLER_17_1764 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_decap_8 FILLER_18_875 ();
 sg13g2_decap_8 FILLER_18_882 ();
 sg13g2_decap_8 FILLER_18_889 ();
 sg13g2_decap_8 FILLER_18_896 ();
 sg13g2_decap_8 FILLER_18_903 ();
 sg13g2_decap_8 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_917 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_decap_8 FILLER_18_938 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_decap_8 FILLER_18_952 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_decap_8 FILLER_18_1029 ();
 sg13g2_decap_8 FILLER_18_1036 ();
 sg13g2_decap_8 FILLER_18_1043 ();
 sg13g2_decap_8 FILLER_18_1050 ();
 sg13g2_decap_8 FILLER_18_1057 ();
 sg13g2_decap_8 FILLER_18_1064 ();
 sg13g2_decap_8 FILLER_18_1071 ();
 sg13g2_decap_8 FILLER_18_1078 ();
 sg13g2_decap_8 FILLER_18_1085 ();
 sg13g2_decap_8 FILLER_18_1092 ();
 sg13g2_decap_8 FILLER_18_1099 ();
 sg13g2_decap_8 FILLER_18_1106 ();
 sg13g2_decap_8 FILLER_18_1113 ();
 sg13g2_decap_8 FILLER_18_1120 ();
 sg13g2_decap_8 FILLER_18_1127 ();
 sg13g2_decap_8 FILLER_18_1134 ();
 sg13g2_decap_8 FILLER_18_1141 ();
 sg13g2_decap_8 FILLER_18_1148 ();
 sg13g2_decap_8 FILLER_18_1155 ();
 sg13g2_decap_8 FILLER_18_1162 ();
 sg13g2_decap_8 FILLER_18_1169 ();
 sg13g2_decap_8 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_decap_8 FILLER_18_1190 ();
 sg13g2_decap_8 FILLER_18_1197 ();
 sg13g2_decap_8 FILLER_18_1204 ();
 sg13g2_decap_8 FILLER_18_1211 ();
 sg13g2_decap_8 FILLER_18_1218 ();
 sg13g2_decap_8 FILLER_18_1225 ();
 sg13g2_decap_8 FILLER_18_1232 ();
 sg13g2_decap_8 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_8 FILLER_18_1274 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_decap_8 FILLER_18_1323 ();
 sg13g2_decap_8 FILLER_18_1330 ();
 sg13g2_decap_8 FILLER_18_1337 ();
 sg13g2_decap_8 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1351 ();
 sg13g2_decap_8 FILLER_18_1358 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1386 ();
 sg13g2_decap_8 FILLER_18_1393 ();
 sg13g2_decap_8 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1407 ();
 sg13g2_decap_8 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1421 ();
 sg13g2_decap_8 FILLER_18_1428 ();
 sg13g2_decap_8 FILLER_18_1435 ();
 sg13g2_decap_8 FILLER_18_1442 ();
 sg13g2_decap_8 FILLER_18_1449 ();
 sg13g2_decap_8 FILLER_18_1456 ();
 sg13g2_decap_8 FILLER_18_1463 ();
 sg13g2_decap_8 FILLER_18_1470 ();
 sg13g2_decap_8 FILLER_18_1477 ();
 sg13g2_decap_8 FILLER_18_1484 ();
 sg13g2_decap_8 FILLER_18_1491 ();
 sg13g2_decap_8 FILLER_18_1498 ();
 sg13g2_decap_8 FILLER_18_1505 ();
 sg13g2_decap_8 FILLER_18_1512 ();
 sg13g2_decap_8 FILLER_18_1519 ();
 sg13g2_decap_8 FILLER_18_1526 ();
 sg13g2_decap_8 FILLER_18_1533 ();
 sg13g2_decap_8 FILLER_18_1540 ();
 sg13g2_decap_8 FILLER_18_1547 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_decap_8 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1589 ();
 sg13g2_decap_8 FILLER_18_1596 ();
 sg13g2_decap_8 FILLER_18_1603 ();
 sg13g2_decap_8 FILLER_18_1610 ();
 sg13g2_decap_8 FILLER_18_1617 ();
 sg13g2_decap_8 FILLER_18_1624 ();
 sg13g2_decap_8 FILLER_18_1631 ();
 sg13g2_decap_8 FILLER_18_1638 ();
 sg13g2_decap_8 FILLER_18_1645 ();
 sg13g2_decap_8 FILLER_18_1652 ();
 sg13g2_decap_8 FILLER_18_1659 ();
 sg13g2_decap_8 FILLER_18_1666 ();
 sg13g2_decap_8 FILLER_18_1673 ();
 sg13g2_decap_8 FILLER_18_1680 ();
 sg13g2_decap_8 FILLER_18_1687 ();
 sg13g2_decap_8 FILLER_18_1694 ();
 sg13g2_decap_8 FILLER_18_1701 ();
 sg13g2_decap_8 FILLER_18_1708 ();
 sg13g2_decap_8 FILLER_18_1715 ();
 sg13g2_decap_8 FILLER_18_1722 ();
 sg13g2_decap_8 FILLER_18_1729 ();
 sg13g2_decap_8 FILLER_18_1736 ();
 sg13g2_decap_8 FILLER_18_1743 ();
 sg13g2_decap_8 FILLER_18_1750 ();
 sg13g2_decap_8 FILLER_18_1757 ();
 sg13g2_decap_4 FILLER_18_1764 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_decap_8 FILLER_19_875 ();
 sg13g2_decap_8 FILLER_19_882 ();
 sg13g2_decap_8 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_8 FILLER_19_903 ();
 sg13g2_decap_8 FILLER_19_910 ();
 sg13g2_decap_8 FILLER_19_917 ();
 sg13g2_decap_8 FILLER_19_924 ();
 sg13g2_decap_8 FILLER_19_931 ();
 sg13g2_decap_8 FILLER_19_938 ();
 sg13g2_decap_8 FILLER_19_945 ();
 sg13g2_decap_8 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_973 ();
 sg13g2_decap_8 FILLER_19_980 ();
 sg13g2_decap_8 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_decap_8 FILLER_19_1029 ();
 sg13g2_decap_8 FILLER_19_1036 ();
 sg13g2_decap_8 FILLER_19_1043 ();
 sg13g2_decap_8 FILLER_19_1050 ();
 sg13g2_decap_8 FILLER_19_1057 ();
 sg13g2_decap_8 FILLER_19_1064 ();
 sg13g2_decap_8 FILLER_19_1071 ();
 sg13g2_decap_8 FILLER_19_1078 ();
 sg13g2_decap_8 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1092 ();
 sg13g2_decap_8 FILLER_19_1099 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1113 ();
 sg13g2_decap_8 FILLER_19_1120 ();
 sg13g2_decap_8 FILLER_19_1127 ();
 sg13g2_decap_8 FILLER_19_1134 ();
 sg13g2_decap_8 FILLER_19_1141 ();
 sg13g2_decap_8 FILLER_19_1148 ();
 sg13g2_decap_8 FILLER_19_1155 ();
 sg13g2_decap_8 FILLER_19_1162 ();
 sg13g2_decap_8 FILLER_19_1169 ();
 sg13g2_decap_8 FILLER_19_1176 ();
 sg13g2_decap_8 FILLER_19_1183 ();
 sg13g2_decap_8 FILLER_19_1190 ();
 sg13g2_decap_8 FILLER_19_1197 ();
 sg13g2_decap_8 FILLER_19_1204 ();
 sg13g2_decap_8 FILLER_19_1211 ();
 sg13g2_decap_8 FILLER_19_1218 ();
 sg13g2_decap_8 FILLER_19_1225 ();
 sg13g2_decap_8 FILLER_19_1232 ();
 sg13g2_decap_8 FILLER_19_1239 ();
 sg13g2_decap_8 FILLER_19_1246 ();
 sg13g2_decap_8 FILLER_19_1253 ();
 sg13g2_decap_8 FILLER_19_1260 ();
 sg13g2_decap_8 FILLER_19_1267 ();
 sg13g2_decap_8 FILLER_19_1274 ();
 sg13g2_decap_8 FILLER_19_1281 ();
 sg13g2_decap_8 FILLER_19_1288 ();
 sg13g2_decap_8 FILLER_19_1295 ();
 sg13g2_decap_8 FILLER_19_1302 ();
 sg13g2_decap_8 FILLER_19_1309 ();
 sg13g2_decap_8 FILLER_19_1316 ();
 sg13g2_decap_8 FILLER_19_1323 ();
 sg13g2_decap_8 FILLER_19_1330 ();
 sg13g2_decap_8 FILLER_19_1337 ();
 sg13g2_decap_8 FILLER_19_1344 ();
 sg13g2_decap_8 FILLER_19_1351 ();
 sg13g2_decap_8 FILLER_19_1358 ();
 sg13g2_decap_8 FILLER_19_1365 ();
 sg13g2_decap_8 FILLER_19_1372 ();
 sg13g2_decap_8 FILLER_19_1379 ();
 sg13g2_decap_8 FILLER_19_1386 ();
 sg13g2_decap_8 FILLER_19_1393 ();
 sg13g2_decap_8 FILLER_19_1400 ();
 sg13g2_decap_8 FILLER_19_1407 ();
 sg13g2_decap_8 FILLER_19_1414 ();
 sg13g2_decap_8 FILLER_19_1421 ();
 sg13g2_decap_8 FILLER_19_1428 ();
 sg13g2_decap_8 FILLER_19_1435 ();
 sg13g2_decap_8 FILLER_19_1442 ();
 sg13g2_decap_8 FILLER_19_1449 ();
 sg13g2_decap_8 FILLER_19_1456 ();
 sg13g2_decap_8 FILLER_19_1463 ();
 sg13g2_decap_8 FILLER_19_1470 ();
 sg13g2_decap_8 FILLER_19_1477 ();
 sg13g2_decap_8 FILLER_19_1484 ();
 sg13g2_decap_8 FILLER_19_1491 ();
 sg13g2_decap_8 FILLER_19_1498 ();
 sg13g2_decap_8 FILLER_19_1505 ();
 sg13g2_decap_8 FILLER_19_1512 ();
 sg13g2_decap_8 FILLER_19_1519 ();
 sg13g2_decap_8 FILLER_19_1526 ();
 sg13g2_decap_8 FILLER_19_1533 ();
 sg13g2_decap_8 FILLER_19_1540 ();
 sg13g2_decap_8 FILLER_19_1547 ();
 sg13g2_decap_8 FILLER_19_1554 ();
 sg13g2_decap_8 FILLER_19_1561 ();
 sg13g2_decap_8 FILLER_19_1568 ();
 sg13g2_decap_8 FILLER_19_1575 ();
 sg13g2_decap_8 FILLER_19_1582 ();
 sg13g2_decap_8 FILLER_19_1589 ();
 sg13g2_decap_8 FILLER_19_1596 ();
 sg13g2_decap_8 FILLER_19_1603 ();
 sg13g2_decap_8 FILLER_19_1610 ();
 sg13g2_decap_8 FILLER_19_1617 ();
 sg13g2_decap_8 FILLER_19_1624 ();
 sg13g2_decap_8 FILLER_19_1631 ();
 sg13g2_decap_8 FILLER_19_1638 ();
 sg13g2_decap_8 FILLER_19_1645 ();
 sg13g2_decap_8 FILLER_19_1652 ();
 sg13g2_decap_8 FILLER_19_1659 ();
 sg13g2_decap_8 FILLER_19_1666 ();
 sg13g2_decap_8 FILLER_19_1673 ();
 sg13g2_decap_8 FILLER_19_1680 ();
 sg13g2_decap_8 FILLER_19_1687 ();
 sg13g2_decap_8 FILLER_19_1694 ();
 sg13g2_decap_8 FILLER_19_1701 ();
 sg13g2_decap_8 FILLER_19_1708 ();
 sg13g2_decap_8 FILLER_19_1715 ();
 sg13g2_decap_8 FILLER_19_1722 ();
 sg13g2_decap_8 FILLER_19_1729 ();
 sg13g2_decap_8 FILLER_19_1736 ();
 sg13g2_decap_8 FILLER_19_1743 ();
 sg13g2_decap_8 FILLER_19_1750 ();
 sg13g2_decap_8 FILLER_19_1757 ();
 sg13g2_decap_4 FILLER_19_1764 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_868 ();
 sg13g2_decap_8 FILLER_20_875 ();
 sg13g2_decap_8 FILLER_20_882 ();
 sg13g2_decap_8 FILLER_20_889 ();
 sg13g2_decap_8 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_903 ();
 sg13g2_decap_8 FILLER_20_910 ();
 sg13g2_decap_8 FILLER_20_917 ();
 sg13g2_decap_8 FILLER_20_924 ();
 sg13g2_decap_8 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_938 ();
 sg13g2_decap_8 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_952 ();
 sg13g2_decap_8 FILLER_20_959 ();
 sg13g2_decap_8 FILLER_20_966 ();
 sg13g2_decap_8 FILLER_20_973 ();
 sg13g2_decap_8 FILLER_20_980 ();
 sg13g2_decap_8 FILLER_20_987 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_decap_8 FILLER_20_1001 ();
 sg13g2_decap_8 FILLER_20_1008 ();
 sg13g2_decap_8 FILLER_20_1015 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_20_1029 ();
 sg13g2_decap_8 FILLER_20_1036 ();
 sg13g2_decap_8 FILLER_20_1043 ();
 sg13g2_decap_8 FILLER_20_1050 ();
 sg13g2_decap_8 FILLER_20_1057 ();
 sg13g2_decap_8 FILLER_20_1064 ();
 sg13g2_decap_8 FILLER_20_1071 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_8 FILLER_20_1099 ();
 sg13g2_decap_8 FILLER_20_1106 ();
 sg13g2_decap_8 FILLER_20_1113 ();
 sg13g2_decap_8 FILLER_20_1120 ();
 sg13g2_decap_8 FILLER_20_1127 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_decap_8 FILLER_20_1141 ();
 sg13g2_decap_8 FILLER_20_1148 ();
 sg13g2_decap_8 FILLER_20_1155 ();
 sg13g2_decap_8 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1169 ();
 sg13g2_decap_8 FILLER_20_1176 ();
 sg13g2_decap_8 FILLER_20_1183 ();
 sg13g2_decap_8 FILLER_20_1190 ();
 sg13g2_decap_8 FILLER_20_1197 ();
 sg13g2_decap_8 FILLER_20_1204 ();
 sg13g2_decap_8 FILLER_20_1211 ();
 sg13g2_decap_8 FILLER_20_1218 ();
 sg13g2_decap_8 FILLER_20_1225 ();
 sg13g2_decap_8 FILLER_20_1232 ();
 sg13g2_decap_8 FILLER_20_1239 ();
 sg13g2_decap_8 FILLER_20_1246 ();
 sg13g2_decap_8 FILLER_20_1253 ();
 sg13g2_decap_8 FILLER_20_1260 ();
 sg13g2_decap_8 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1274 ();
 sg13g2_decap_8 FILLER_20_1281 ();
 sg13g2_decap_8 FILLER_20_1288 ();
 sg13g2_decap_8 FILLER_20_1295 ();
 sg13g2_decap_8 FILLER_20_1302 ();
 sg13g2_decap_8 FILLER_20_1309 ();
 sg13g2_decap_8 FILLER_20_1316 ();
 sg13g2_decap_8 FILLER_20_1323 ();
 sg13g2_decap_8 FILLER_20_1330 ();
 sg13g2_decap_8 FILLER_20_1337 ();
 sg13g2_decap_8 FILLER_20_1344 ();
 sg13g2_decap_8 FILLER_20_1351 ();
 sg13g2_decap_8 FILLER_20_1358 ();
 sg13g2_decap_8 FILLER_20_1365 ();
 sg13g2_decap_8 FILLER_20_1372 ();
 sg13g2_decap_8 FILLER_20_1379 ();
 sg13g2_decap_8 FILLER_20_1386 ();
 sg13g2_decap_8 FILLER_20_1393 ();
 sg13g2_decap_8 FILLER_20_1400 ();
 sg13g2_decap_8 FILLER_20_1407 ();
 sg13g2_decap_8 FILLER_20_1414 ();
 sg13g2_decap_8 FILLER_20_1421 ();
 sg13g2_decap_8 FILLER_20_1428 ();
 sg13g2_decap_8 FILLER_20_1435 ();
 sg13g2_decap_8 FILLER_20_1442 ();
 sg13g2_decap_8 FILLER_20_1449 ();
 sg13g2_decap_8 FILLER_20_1456 ();
 sg13g2_decap_8 FILLER_20_1463 ();
 sg13g2_decap_8 FILLER_20_1470 ();
 sg13g2_decap_8 FILLER_20_1477 ();
 sg13g2_decap_8 FILLER_20_1484 ();
 sg13g2_decap_8 FILLER_20_1491 ();
 sg13g2_decap_8 FILLER_20_1498 ();
 sg13g2_decap_8 FILLER_20_1505 ();
 sg13g2_decap_8 FILLER_20_1512 ();
 sg13g2_decap_8 FILLER_20_1519 ();
 sg13g2_decap_8 FILLER_20_1526 ();
 sg13g2_decap_8 FILLER_20_1533 ();
 sg13g2_decap_8 FILLER_20_1540 ();
 sg13g2_decap_8 FILLER_20_1547 ();
 sg13g2_decap_8 FILLER_20_1554 ();
 sg13g2_decap_8 FILLER_20_1561 ();
 sg13g2_decap_8 FILLER_20_1568 ();
 sg13g2_decap_8 FILLER_20_1575 ();
 sg13g2_decap_8 FILLER_20_1582 ();
 sg13g2_decap_8 FILLER_20_1589 ();
 sg13g2_decap_8 FILLER_20_1596 ();
 sg13g2_decap_8 FILLER_20_1603 ();
 sg13g2_decap_8 FILLER_20_1610 ();
 sg13g2_decap_8 FILLER_20_1617 ();
 sg13g2_decap_8 FILLER_20_1624 ();
 sg13g2_decap_8 FILLER_20_1631 ();
 sg13g2_decap_8 FILLER_20_1638 ();
 sg13g2_decap_8 FILLER_20_1645 ();
 sg13g2_decap_8 FILLER_20_1652 ();
 sg13g2_decap_8 FILLER_20_1659 ();
 sg13g2_decap_8 FILLER_20_1666 ();
 sg13g2_decap_8 FILLER_20_1673 ();
 sg13g2_decap_8 FILLER_20_1680 ();
 sg13g2_decap_8 FILLER_20_1687 ();
 sg13g2_decap_8 FILLER_20_1694 ();
 sg13g2_decap_8 FILLER_20_1701 ();
 sg13g2_decap_8 FILLER_20_1708 ();
 sg13g2_decap_8 FILLER_20_1715 ();
 sg13g2_decap_8 FILLER_20_1722 ();
 sg13g2_decap_8 FILLER_20_1729 ();
 sg13g2_decap_8 FILLER_20_1736 ();
 sg13g2_decap_8 FILLER_20_1743 ();
 sg13g2_decap_8 FILLER_20_1750 ();
 sg13g2_decap_8 FILLER_20_1757 ();
 sg13g2_decap_4 FILLER_20_1764 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_917 ();
 sg13g2_decap_8 FILLER_21_924 ();
 sg13g2_decap_8 FILLER_21_931 ();
 sg13g2_decap_8 FILLER_21_938 ();
 sg13g2_decap_8 FILLER_21_945 ();
 sg13g2_decap_8 FILLER_21_952 ();
 sg13g2_decap_8 FILLER_21_959 ();
 sg13g2_decap_8 FILLER_21_966 ();
 sg13g2_decap_8 FILLER_21_973 ();
 sg13g2_decap_8 FILLER_21_980 ();
 sg13g2_decap_8 FILLER_21_987 ();
 sg13g2_decap_8 FILLER_21_994 ();
 sg13g2_decap_8 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_8 FILLER_21_1029 ();
 sg13g2_decap_8 FILLER_21_1036 ();
 sg13g2_decap_8 FILLER_21_1043 ();
 sg13g2_decap_8 FILLER_21_1050 ();
 sg13g2_decap_8 FILLER_21_1057 ();
 sg13g2_decap_8 FILLER_21_1064 ();
 sg13g2_decap_8 FILLER_21_1071 ();
 sg13g2_decap_8 FILLER_21_1078 ();
 sg13g2_decap_8 FILLER_21_1085 ();
 sg13g2_decap_8 FILLER_21_1092 ();
 sg13g2_decap_8 FILLER_21_1099 ();
 sg13g2_decap_8 FILLER_21_1106 ();
 sg13g2_decap_8 FILLER_21_1113 ();
 sg13g2_decap_8 FILLER_21_1120 ();
 sg13g2_decap_8 FILLER_21_1127 ();
 sg13g2_decap_8 FILLER_21_1134 ();
 sg13g2_decap_8 FILLER_21_1141 ();
 sg13g2_decap_8 FILLER_21_1148 ();
 sg13g2_decap_8 FILLER_21_1155 ();
 sg13g2_decap_8 FILLER_21_1162 ();
 sg13g2_decap_8 FILLER_21_1169 ();
 sg13g2_decap_8 FILLER_21_1176 ();
 sg13g2_decap_8 FILLER_21_1183 ();
 sg13g2_decap_8 FILLER_21_1190 ();
 sg13g2_decap_8 FILLER_21_1197 ();
 sg13g2_decap_8 FILLER_21_1204 ();
 sg13g2_decap_8 FILLER_21_1211 ();
 sg13g2_decap_8 FILLER_21_1218 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1239 ();
 sg13g2_decap_8 FILLER_21_1246 ();
 sg13g2_decap_8 FILLER_21_1253 ();
 sg13g2_decap_8 FILLER_21_1260 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1274 ();
 sg13g2_decap_8 FILLER_21_1281 ();
 sg13g2_decap_8 FILLER_21_1288 ();
 sg13g2_decap_8 FILLER_21_1295 ();
 sg13g2_decap_8 FILLER_21_1302 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_decap_8 FILLER_21_1316 ();
 sg13g2_decap_8 FILLER_21_1323 ();
 sg13g2_decap_8 FILLER_21_1330 ();
 sg13g2_decap_8 FILLER_21_1337 ();
 sg13g2_decap_8 FILLER_21_1344 ();
 sg13g2_decap_8 FILLER_21_1351 ();
 sg13g2_decap_8 FILLER_21_1358 ();
 sg13g2_decap_8 FILLER_21_1365 ();
 sg13g2_decap_8 FILLER_21_1372 ();
 sg13g2_decap_8 FILLER_21_1379 ();
 sg13g2_decap_8 FILLER_21_1386 ();
 sg13g2_decap_8 FILLER_21_1393 ();
 sg13g2_decap_8 FILLER_21_1400 ();
 sg13g2_decap_8 FILLER_21_1407 ();
 sg13g2_decap_8 FILLER_21_1414 ();
 sg13g2_decap_8 FILLER_21_1421 ();
 sg13g2_decap_8 FILLER_21_1428 ();
 sg13g2_decap_8 FILLER_21_1435 ();
 sg13g2_decap_8 FILLER_21_1442 ();
 sg13g2_decap_8 FILLER_21_1449 ();
 sg13g2_decap_8 FILLER_21_1456 ();
 sg13g2_decap_8 FILLER_21_1463 ();
 sg13g2_decap_8 FILLER_21_1470 ();
 sg13g2_decap_8 FILLER_21_1477 ();
 sg13g2_decap_8 FILLER_21_1484 ();
 sg13g2_decap_8 FILLER_21_1491 ();
 sg13g2_decap_8 FILLER_21_1498 ();
 sg13g2_decap_8 FILLER_21_1505 ();
 sg13g2_decap_8 FILLER_21_1512 ();
 sg13g2_decap_8 FILLER_21_1519 ();
 sg13g2_decap_8 FILLER_21_1526 ();
 sg13g2_decap_8 FILLER_21_1533 ();
 sg13g2_decap_8 FILLER_21_1540 ();
 sg13g2_decap_8 FILLER_21_1547 ();
 sg13g2_decap_8 FILLER_21_1554 ();
 sg13g2_decap_8 FILLER_21_1561 ();
 sg13g2_decap_8 FILLER_21_1568 ();
 sg13g2_decap_8 FILLER_21_1575 ();
 sg13g2_decap_8 FILLER_21_1582 ();
 sg13g2_decap_8 FILLER_21_1589 ();
 sg13g2_decap_8 FILLER_21_1596 ();
 sg13g2_decap_8 FILLER_21_1603 ();
 sg13g2_decap_8 FILLER_21_1610 ();
 sg13g2_decap_8 FILLER_21_1617 ();
 sg13g2_decap_8 FILLER_21_1624 ();
 sg13g2_decap_8 FILLER_21_1631 ();
 sg13g2_decap_8 FILLER_21_1638 ();
 sg13g2_decap_8 FILLER_21_1645 ();
 sg13g2_decap_8 FILLER_21_1652 ();
 sg13g2_decap_8 FILLER_21_1659 ();
 sg13g2_decap_8 FILLER_21_1666 ();
 sg13g2_decap_8 FILLER_21_1673 ();
 sg13g2_decap_8 FILLER_21_1680 ();
 sg13g2_decap_8 FILLER_21_1687 ();
 sg13g2_decap_8 FILLER_21_1694 ();
 sg13g2_decap_8 FILLER_21_1701 ();
 sg13g2_decap_8 FILLER_21_1708 ();
 sg13g2_decap_8 FILLER_21_1715 ();
 sg13g2_decap_8 FILLER_21_1722 ();
 sg13g2_decap_8 FILLER_21_1729 ();
 sg13g2_decap_8 FILLER_21_1736 ();
 sg13g2_decap_8 FILLER_21_1743 ();
 sg13g2_decap_8 FILLER_21_1750 ();
 sg13g2_decap_8 FILLER_21_1757 ();
 sg13g2_decap_4 FILLER_21_1764 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_decap_8 FILLER_22_875 ();
 sg13g2_decap_8 FILLER_22_882 ();
 sg13g2_decap_8 FILLER_22_889 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_decap_8 FILLER_22_903 ();
 sg13g2_decap_8 FILLER_22_910 ();
 sg13g2_decap_8 FILLER_22_917 ();
 sg13g2_decap_8 FILLER_22_924 ();
 sg13g2_decap_8 FILLER_22_931 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_8 FILLER_22_959 ();
 sg13g2_decap_8 FILLER_22_966 ();
 sg13g2_decap_8 FILLER_22_973 ();
 sg13g2_decap_8 FILLER_22_980 ();
 sg13g2_decap_8 FILLER_22_987 ();
 sg13g2_decap_8 FILLER_22_994 ();
 sg13g2_decap_8 FILLER_22_1001 ();
 sg13g2_decap_8 FILLER_22_1008 ();
 sg13g2_decap_8 FILLER_22_1015 ();
 sg13g2_decap_8 FILLER_22_1022 ();
 sg13g2_decap_8 FILLER_22_1029 ();
 sg13g2_decap_8 FILLER_22_1036 ();
 sg13g2_decap_8 FILLER_22_1043 ();
 sg13g2_decap_8 FILLER_22_1050 ();
 sg13g2_decap_8 FILLER_22_1057 ();
 sg13g2_decap_8 FILLER_22_1064 ();
 sg13g2_decap_8 FILLER_22_1071 ();
 sg13g2_decap_8 FILLER_22_1078 ();
 sg13g2_decap_8 FILLER_22_1085 ();
 sg13g2_decap_8 FILLER_22_1092 ();
 sg13g2_decap_8 FILLER_22_1099 ();
 sg13g2_decap_8 FILLER_22_1106 ();
 sg13g2_decap_8 FILLER_22_1113 ();
 sg13g2_decap_8 FILLER_22_1120 ();
 sg13g2_decap_8 FILLER_22_1127 ();
 sg13g2_decap_8 FILLER_22_1134 ();
 sg13g2_decap_8 FILLER_22_1141 ();
 sg13g2_decap_8 FILLER_22_1148 ();
 sg13g2_decap_8 FILLER_22_1155 ();
 sg13g2_decap_8 FILLER_22_1162 ();
 sg13g2_decap_8 FILLER_22_1169 ();
 sg13g2_decap_8 FILLER_22_1176 ();
 sg13g2_decap_8 FILLER_22_1183 ();
 sg13g2_decap_8 FILLER_22_1190 ();
 sg13g2_decap_8 FILLER_22_1197 ();
 sg13g2_decap_8 FILLER_22_1204 ();
 sg13g2_decap_8 FILLER_22_1211 ();
 sg13g2_decap_8 FILLER_22_1218 ();
 sg13g2_decap_8 FILLER_22_1225 ();
 sg13g2_decap_8 FILLER_22_1232 ();
 sg13g2_decap_8 FILLER_22_1239 ();
 sg13g2_decap_8 FILLER_22_1246 ();
 sg13g2_decap_8 FILLER_22_1253 ();
 sg13g2_decap_8 FILLER_22_1260 ();
 sg13g2_decap_8 FILLER_22_1267 ();
 sg13g2_decap_8 FILLER_22_1274 ();
 sg13g2_decap_8 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1288 ();
 sg13g2_decap_8 FILLER_22_1295 ();
 sg13g2_decap_8 FILLER_22_1302 ();
 sg13g2_decap_8 FILLER_22_1309 ();
 sg13g2_decap_8 FILLER_22_1316 ();
 sg13g2_decap_8 FILLER_22_1323 ();
 sg13g2_decap_8 FILLER_22_1330 ();
 sg13g2_decap_8 FILLER_22_1337 ();
 sg13g2_decap_8 FILLER_22_1344 ();
 sg13g2_decap_8 FILLER_22_1351 ();
 sg13g2_decap_8 FILLER_22_1358 ();
 sg13g2_decap_8 FILLER_22_1365 ();
 sg13g2_decap_8 FILLER_22_1372 ();
 sg13g2_decap_8 FILLER_22_1379 ();
 sg13g2_decap_8 FILLER_22_1386 ();
 sg13g2_decap_8 FILLER_22_1393 ();
 sg13g2_decap_8 FILLER_22_1400 ();
 sg13g2_decap_8 FILLER_22_1407 ();
 sg13g2_decap_8 FILLER_22_1414 ();
 sg13g2_decap_8 FILLER_22_1421 ();
 sg13g2_decap_8 FILLER_22_1428 ();
 sg13g2_decap_8 FILLER_22_1435 ();
 sg13g2_decap_8 FILLER_22_1442 ();
 sg13g2_decap_8 FILLER_22_1449 ();
 sg13g2_decap_8 FILLER_22_1456 ();
 sg13g2_decap_8 FILLER_22_1463 ();
 sg13g2_decap_8 FILLER_22_1470 ();
 sg13g2_decap_8 FILLER_22_1477 ();
 sg13g2_decap_8 FILLER_22_1484 ();
 sg13g2_decap_8 FILLER_22_1491 ();
 sg13g2_decap_8 FILLER_22_1498 ();
 sg13g2_decap_8 FILLER_22_1505 ();
 sg13g2_decap_8 FILLER_22_1512 ();
 sg13g2_decap_8 FILLER_22_1519 ();
 sg13g2_decap_8 FILLER_22_1526 ();
 sg13g2_decap_8 FILLER_22_1533 ();
 sg13g2_decap_8 FILLER_22_1540 ();
 sg13g2_decap_8 FILLER_22_1547 ();
 sg13g2_decap_8 FILLER_22_1554 ();
 sg13g2_decap_8 FILLER_22_1561 ();
 sg13g2_decap_8 FILLER_22_1568 ();
 sg13g2_decap_8 FILLER_22_1575 ();
 sg13g2_decap_8 FILLER_22_1582 ();
 sg13g2_decap_8 FILLER_22_1589 ();
 sg13g2_decap_8 FILLER_22_1596 ();
 sg13g2_decap_8 FILLER_22_1603 ();
 sg13g2_decap_8 FILLER_22_1610 ();
 sg13g2_decap_8 FILLER_22_1617 ();
 sg13g2_decap_8 FILLER_22_1624 ();
 sg13g2_decap_8 FILLER_22_1631 ();
 sg13g2_decap_8 FILLER_22_1638 ();
 sg13g2_decap_8 FILLER_22_1645 ();
 sg13g2_decap_8 FILLER_22_1652 ();
 sg13g2_decap_8 FILLER_22_1659 ();
 sg13g2_decap_8 FILLER_22_1666 ();
 sg13g2_decap_8 FILLER_22_1673 ();
 sg13g2_decap_8 FILLER_22_1680 ();
 sg13g2_decap_8 FILLER_22_1687 ();
 sg13g2_decap_8 FILLER_22_1694 ();
 sg13g2_decap_8 FILLER_22_1701 ();
 sg13g2_decap_8 FILLER_22_1708 ();
 sg13g2_decap_8 FILLER_22_1715 ();
 sg13g2_decap_8 FILLER_22_1722 ();
 sg13g2_decap_8 FILLER_22_1729 ();
 sg13g2_decap_8 FILLER_22_1736 ();
 sg13g2_decap_8 FILLER_22_1743 ();
 sg13g2_decap_8 FILLER_22_1750 ();
 sg13g2_decap_8 FILLER_22_1757 ();
 sg13g2_decap_4 FILLER_22_1764 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_decap_8 FILLER_23_882 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_decap_8 FILLER_23_903 ();
 sg13g2_decap_8 FILLER_23_910 ();
 sg13g2_decap_8 FILLER_23_917 ();
 sg13g2_decap_8 FILLER_23_924 ();
 sg13g2_decap_8 FILLER_23_931 ();
 sg13g2_decap_8 FILLER_23_938 ();
 sg13g2_decap_8 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_952 ();
 sg13g2_decap_8 FILLER_23_959 ();
 sg13g2_decap_8 FILLER_23_966 ();
 sg13g2_decap_8 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_decap_8 FILLER_23_987 ();
 sg13g2_decap_8 FILLER_23_994 ();
 sg13g2_decap_8 FILLER_23_1001 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1015 ();
 sg13g2_decap_8 FILLER_23_1022 ();
 sg13g2_decap_8 FILLER_23_1029 ();
 sg13g2_decap_8 FILLER_23_1036 ();
 sg13g2_decap_8 FILLER_23_1043 ();
 sg13g2_decap_8 FILLER_23_1050 ();
 sg13g2_decap_8 FILLER_23_1057 ();
 sg13g2_decap_8 FILLER_23_1064 ();
 sg13g2_decap_8 FILLER_23_1071 ();
 sg13g2_decap_8 FILLER_23_1078 ();
 sg13g2_decap_8 FILLER_23_1085 ();
 sg13g2_decap_8 FILLER_23_1092 ();
 sg13g2_decap_8 FILLER_23_1099 ();
 sg13g2_decap_8 FILLER_23_1106 ();
 sg13g2_decap_8 FILLER_23_1113 ();
 sg13g2_decap_8 FILLER_23_1120 ();
 sg13g2_decap_8 FILLER_23_1127 ();
 sg13g2_decap_8 FILLER_23_1134 ();
 sg13g2_decap_8 FILLER_23_1141 ();
 sg13g2_decap_8 FILLER_23_1148 ();
 sg13g2_decap_8 FILLER_23_1155 ();
 sg13g2_decap_8 FILLER_23_1162 ();
 sg13g2_decap_8 FILLER_23_1169 ();
 sg13g2_decap_8 FILLER_23_1176 ();
 sg13g2_decap_8 FILLER_23_1183 ();
 sg13g2_decap_8 FILLER_23_1190 ();
 sg13g2_decap_8 FILLER_23_1197 ();
 sg13g2_decap_8 FILLER_23_1204 ();
 sg13g2_decap_8 FILLER_23_1211 ();
 sg13g2_decap_8 FILLER_23_1218 ();
 sg13g2_decap_8 FILLER_23_1225 ();
 sg13g2_decap_8 FILLER_23_1232 ();
 sg13g2_decap_8 FILLER_23_1239 ();
 sg13g2_decap_8 FILLER_23_1246 ();
 sg13g2_decap_8 FILLER_23_1253 ();
 sg13g2_decap_8 FILLER_23_1260 ();
 sg13g2_decap_8 FILLER_23_1267 ();
 sg13g2_decap_8 FILLER_23_1274 ();
 sg13g2_decap_8 FILLER_23_1281 ();
 sg13g2_decap_8 FILLER_23_1288 ();
 sg13g2_decap_8 FILLER_23_1295 ();
 sg13g2_decap_8 FILLER_23_1302 ();
 sg13g2_decap_8 FILLER_23_1309 ();
 sg13g2_decap_8 FILLER_23_1316 ();
 sg13g2_decap_8 FILLER_23_1323 ();
 sg13g2_decap_8 FILLER_23_1330 ();
 sg13g2_decap_8 FILLER_23_1337 ();
 sg13g2_decap_8 FILLER_23_1344 ();
 sg13g2_decap_8 FILLER_23_1351 ();
 sg13g2_decap_8 FILLER_23_1358 ();
 sg13g2_decap_8 FILLER_23_1365 ();
 sg13g2_decap_8 FILLER_23_1372 ();
 sg13g2_decap_8 FILLER_23_1379 ();
 sg13g2_decap_8 FILLER_23_1386 ();
 sg13g2_decap_8 FILLER_23_1393 ();
 sg13g2_decap_8 FILLER_23_1400 ();
 sg13g2_decap_8 FILLER_23_1407 ();
 sg13g2_decap_8 FILLER_23_1414 ();
 sg13g2_decap_8 FILLER_23_1421 ();
 sg13g2_decap_8 FILLER_23_1428 ();
 sg13g2_decap_8 FILLER_23_1435 ();
 sg13g2_decap_8 FILLER_23_1442 ();
 sg13g2_decap_8 FILLER_23_1449 ();
 sg13g2_decap_8 FILLER_23_1456 ();
 sg13g2_decap_8 FILLER_23_1463 ();
 sg13g2_decap_8 FILLER_23_1470 ();
 sg13g2_decap_8 FILLER_23_1477 ();
 sg13g2_decap_8 FILLER_23_1484 ();
 sg13g2_decap_8 FILLER_23_1491 ();
 sg13g2_decap_8 FILLER_23_1498 ();
 sg13g2_decap_8 FILLER_23_1505 ();
 sg13g2_decap_8 FILLER_23_1512 ();
 sg13g2_decap_8 FILLER_23_1519 ();
 sg13g2_decap_8 FILLER_23_1526 ();
 sg13g2_decap_8 FILLER_23_1533 ();
 sg13g2_decap_8 FILLER_23_1540 ();
 sg13g2_decap_8 FILLER_23_1547 ();
 sg13g2_decap_8 FILLER_23_1554 ();
 sg13g2_decap_8 FILLER_23_1561 ();
 sg13g2_decap_8 FILLER_23_1568 ();
 sg13g2_decap_8 FILLER_23_1575 ();
 sg13g2_decap_8 FILLER_23_1582 ();
 sg13g2_decap_8 FILLER_23_1589 ();
 sg13g2_decap_8 FILLER_23_1596 ();
 sg13g2_decap_8 FILLER_23_1603 ();
 sg13g2_decap_8 FILLER_23_1610 ();
 sg13g2_decap_8 FILLER_23_1617 ();
 sg13g2_decap_8 FILLER_23_1624 ();
 sg13g2_decap_8 FILLER_23_1631 ();
 sg13g2_decap_8 FILLER_23_1638 ();
 sg13g2_decap_8 FILLER_23_1645 ();
 sg13g2_decap_8 FILLER_23_1652 ();
 sg13g2_decap_8 FILLER_23_1659 ();
 sg13g2_decap_8 FILLER_23_1666 ();
 sg13g2_decap_8 FILLER_23_1673 ();
 sg13g2_decap_8 FILLER_23_1680 ();
 sg13g2_decap_8 FILLER_23_1687 ();
 sg13g2_decap_8 FILLER_23_1694 ();
 sg13g2_decap_8 FILLER_23_1701 ();
 sg13g2_decap_8 FILLER_23_1708 ();
 sg13g2_decap_8 FILLER_23_1715 ();
 sg13g2_decap_8 FILLER_23_1722 ();
 sg13g2_decap_8 FILLER_23_1729 ();
 sg13g2_decap_8 FILLER_23_1736 ();
 sg13g2_decap_8 FILLER_23_1743 ();
 sg13g2_decap_8 FILLER_23_1750 ();
 sg13g2_decap_8 FILLER_23_1757 ();
 sg13g2_decap_4 FILLER_23_1764 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_decap_8 FILLER_24_875 ();
 sg13g2_decap_8 FILLER_24_882 ();
 sg13g2_decap_8 FILLER_24_889 ();
 sg13g2_decap_8 FILLER_24_896 ();
 sg13g2_decap_8 FILLER_24_903 ();
 sg13g2_decap_8 FILLER_24_910 ();
 sg13g2_decap_8 FILLER_24_917 ();
 sg13g2_decap_8 FILLER_24_924 ();
 sg13g2_decap_8 FILLER_24_931 ();
 sg13g2_decap_8 FILLER_24_938 ();
 sg13g2_decap_8 FILLER_24_945 ();
 sg13g2_decap_8 FILLER_24_952 ();
 sg13g2_decap_8 FILLER_24_959 ();
 sg13g2_decap_8 FILLER_24_966 ();
 sg13g2_decap_8 FILLER_24_973 ();
 sg13g2_decap_8 FILLER_24_980 ();
 sg13g2_decap_8 FILLER_24_987 ();
 sg13g2_decap_8 FILLER_24_994 ();
 sg13g2_decap_8 FILLER_24_1001 ();
 sg13g2_decap_8 FILLER_24_1008 ();
 sg13g2_decap_8 FILLER_24_1015 ();
 sg13g2_decap_8 FILLER_24_1022 ();
 sg13g2_decap_8 FILLER_24_1029 ();
 sg13g2_decap_8 FILLER_24_1036 ();
 sg13g2_decap_8 FILLER_24_1043 ();
 sg13g2_decap_8 FILLER_24_1050 ();
 sg13g2_decap_8 FILLER_24_1057 ();
 sg13g2_decap_8 FILLER_24_1064 ();
 sg13g2_decap_8 FILLER_24_1071 ();
 sg13g2_decap_8 FILLER_24_1078 ();
 sg13g2_decap_8 FILLER_24_1085 ();
 sg13g2_decap_8 FILLER_24_1092 ();
 sg13g2_decap_8 FILLER_24_1099 ();
 sg13g2_decap_8 FILLER_24_1106 ();
 sg13g2_decap_8 FILLER_24_1113 ();
 sg13g2_decap_8 FILLER_24_1120 ();
 sg13g2_decap_8 FILLER_24_1127 ();
 sg13g2_decap_8 FILLER_24_1134 ();
 sg13g2_decap_8 FILLER_24_1141 ();
 sg13g2_decap_8 FILLER_24_1148 ();
 sg13g2_decap_8 FILLER_24_1155 ();
 sg13g2_decap_8 FILLER_24_1162 ();
 sg13g2_decap_8 FILLER_24_1169 ();
 sg13g2_decap_8 FILLER_24_1176 ();
 sg13g2_decap_8 FILLER_24_1183 ();
 sg13g2_decap_8 FILLER_24_1190 ();
 sg13g2_decap_8 FILLER_24_1197 ();
 sg13g2_decap_8 FILLER_24_1204 ();
 sg13g2_decap_8 FILLER_24_1211 ();
 sg13g2_decap_8 FILLER_24_1218 ();
 sg13g2_decap_8 FILLER_24_1225 ();
 sg13g2_decap_8 FILLER_24_1232 ();
 sg13g2_decap_8 FILLER_24_1239 ();
 sg13g2_decap_8 FILLER_24_1246 ();
 sg13g2_decap_8 FILLER_24_1253 ();
 sg13g2_decap_8 FILLER_24_1260 ();
 sg13g2_decap_8 FILLER_24_1267 ();
 sg13g2_decap_8 FILLER_24_1274 ();
 sg13g2_decap_8 FILLER_24_1281 ();
 sg13g2_decap_8 FILLER_24_1288 ();
 sg13g2_decap_8 FILLER_24_1295 ();
 sg13g2_decap_8 FILLER_24_1302 ();
 sg13g2_decap_8 FILLER_24_1309 ();
 sg13g2_decap_8 FILLER_24_1316 ();
 sg13g2_decap_8 FILLER_24_1323 ();
 sg13g2_decap_8 FILLER_24_1330 ();
 sg13g2_decap_8 FILLER_24_1337 ();
 sg13g2_decap_8 FILLER_24_1344 ();
 sg13g2_decap_8 FILLER_24_1351 ();
 sg13g2_decap_8 FILLER_24_1358 ();
 sg13g2_decap_8 FILLER_24_1365 ();
 sg13g2_decap_8 FILLER_24_1372 ();
 sg13g2_decap_8 FILLER_24_1379 ();
 sg13g2_decap_8 FILLER_24_1386 ();
 sg13g2_decap_8 FILLER_24_1393 ();
 sg13g2_decap_8 FILLER_24_1400 ();
 sg13g2_decap_8 FILLER_24_1407 ();
 sg13g2_decap_8 FILLER_24_1414 ();
 sg13g2_decap_8 FILLER_24_1421 ();
 sg13g2_decap_8 FILLER_24_1428 ();
 sg13g2_decap_8 FILLER_24_1435 ();
 sg13g2_decap_8 FILLER_24_1442 ();
 sg13g2_decap_8 FILLER_24_1449 ();
 sg13g2_decap_8 FILLER_24_1456 ();
 sg13g2_decap_8 FILLER_24_1463 ();
 sg13g2_decap_8 FILLER_24_1470 ();
 sg13g2_decap_8 FILLER_24_1477 ();
 sg13g2_decap_8 FILLER_24_1484 ();
 sg13g2_decap_8 FILLER_24_1491 ();
 sg13g2_decap_8 FILLER_24_1498 ();
 sg13g2_decap_8 FILLER_24_1505 ();
 sg13g2_decap_8 FILLER_24_1512 ();
 sg13g2_decap_8 FILLER_24_1519 ();
 sg13g2_decap_8 FILLER_24_1526 ();
 sg13g2_decap_8 FILLER_24_1533 ();
 sg13g2_decap_8 FILLER_24_1540 ();
 sg13g2_decap_8 FILLER_24_1547 ();
 sg13g2_decap_8 FILLER_24_1554 ();
 sg13g2_decap_8 FILLER_24_1561 ();
 sg13g2_decap_8 FILLER_24_1568 ();
 sg13g2_decap_8 FILLER_24_1575 ();
 sg13g2_decap_8 FILLER_24_1582 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_decap_8 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_decap_8 FILLER_24_1652 ();
 sg13g2_decap_8 FILLER_24_1659 ();
 sg13g2_decap_8 FILLER_24_1666 ();
 sg13g2_decap_8 FILLER_24_1673 ();
 sg13g2_decap_8 FILLER_24_1680 ();
 sg13g2_decap_8 FILLER_24_1687 ();
 sg13g2_decap_8 FILLER_24_1694 ();
 sg13g2_decap_8 FILLER_24_1701 ();
 sg13g2_decap_8 FILLER_24_1708 ();
 sg13g2_decap_8 FILLER_24_1715 ();
 sg13g2_decap_8 FILLER_24_1722 ();
 sg13g2_decap_8 FILLER_24_1729 ();
 sg13g2_decap_8 FILLER_24_1736 ();
 sg13g2_decap_8 FILLER_24_1743 ();
 sg13g2_decap_8 FILLER_24_1750 ();
 sg13g2_decap_8 FILLER_24_1757 ();
 sg13g2_decap_4 FILLER_24_1764 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_889 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_decap_8 FILLER_25_903 ();
 sg13g2_decap_8 FILLER_25_910 ();
 sg13g2_decap_8 FILLER_25_917 ();
 sg13g2_decap_8 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_931 ();
 sg13g2_decap_8 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_973 ();
 sg13g2_decap_8 FILLER_25_980 ();
 sg13g2_decap_8 FILLER_25_987 ();
 sg13g2_decap_8 FILLER_25_994 ();
 sg13g2_decap_8 FILLER_25_1001 ();
 sg13g2_decap_8 FILLER_25_1008 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1022 ();
 sg13g2_decap_8 FILLER_25_1029 ();
 sg13g2_decap_8 FILLER_25_1036 ();
 sg13g2_decap_8 FILLER_25_1043 ();
 sg13g2_decap_8 FILLER_25_1050 ();
 sg13g2_decap_8 FILLER_25_1057 ();
 sg13g2_decap_8 FILLER_25_1064 ();
 sg13g2_decap_8 FILLER_25_1071 ();
 sg13g2_decap_8 FILLER_25_1078 ();
 sg13g2_decap_8 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1092 ();
 sg13g2_decap_8 FILLER_25_1099 ();
 sg13g2_decap_8 FILLER_25_1106 ();
 sg13g2_decap_8 FILLER_25_1113 ();
 sg13g2_decap_8 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1127 ();
 sg13g2_decap_8 FILLER_25_1134 ();
 sg13g2_decap_8 FILLER_25_1141 ();
 sg13g2_decap_8 FILLER_25_1148 ();
 sg13g2_decap_8 FILLER_25_1155 ();
 sg13g2_decap_8 FILLER_25_1162 ();
 sg13g2_decap_8 FILLER_25_1169 ();
 sg13g2_decap_8 FILLER_25_1176 ();
 sg13g2_decap_8 FILLER_25_1183 ();
 sg13g2_decap_8 FILLER_25_1190 ();
 sg13g2_decap_8 FILLER_25_1197 ();
 sg13g2_decap_8 FILLER_25_1204 ();
 sg13g2_decap_8 FILLER_25_1211 ();
 sg13g2_decap_8 FILLER_25_1218 ();
 sg13g2_decap_8 FILLER_25_1225 ();
 sg13g2_decap_8 FILLER_25_1232 ();
 sg13g2_decap_8 FILLER_25_1239 ();
 sg13g2_decap_8 FILLER_25_1246 ();
 sg13g2_decap_8 FILLER_25_1253 ();
 sg13g2_decap_8 FILLER_25_1260 ();
 sg13g2_decap_8 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1274 ();
 sg13g2_decap_8 FILLER_25_1281 ();
 sg13g2_decap_8 FILLER_25_1288 ();
 sg13g2_decap_8 FILLER_25_1295 ();
 sg13g2_decap_8 FILLER_25_1302 ();
 sg13g2_decap_8 FILLER_25_1309 ();
 sg13g2_decap_8 FILLER_25_1316 ();
 sg13g2_decap_8 FILLER_25_1323 ();
 sg13g2_decap_8 FILLER_25_1330 ();
 sg13g2_decap_8 FILLER_25_1337 ();
 sg13g2_decap_8 FILLER_25_1344 ();
 sg13g2_decap_8 FILLER_25_1351 ();
 sg13g2_decap_8 FILLER_25_1358 ();
 sg13g2_decap_8 FILLER_25_1365 ();
 sg13g2_decap_8 FILLER_25_1372 ();
 sg13g2_decap_8 FILLER_25_1379 ();
 sg13g2_decap_8 FILLER_25_1386 ();
 sg13g2_decap_8 FILLER_25_1393 ();
 sg13g2_decap_8 FILLER_25_1400 ();
 sg13g2_decap_8 FILLER_25_1407 ();
 sg13g2_decap_8 FILLER_25_1414 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_decap_8 FILLER_25_1428 ();
 sg13g2_decap_8 FILLER_25_1435 ();
 sg13g2_decap_8 FILLER_25_1442 ();
 sg13g2_decap_8 FILLER_25_1449 ();
 sg13g2_decap_8 FILLER_25_1456 ();
 sg13g2_decap_8 FILLER_25_1463 ();
 sg13g2_decap_8 FILLER_25_1470 ();
 sg13g2_decap_8 FILLER_25_1477 ();
 sg13g2_decap_8 FILLER_25_1484 ();
 sg13g2_decap_8 FILLER_25_1491 ();
 sg13g2_decap_8 FILLER_25_1498 ();
 sg13g2_decap_8 FILLER_25_1505 ();
 sg13g2_decap_8 FILLER_25_1512 ();
 sg13g2_decap_8 FILLER_25_1519 ();
 sg13g2_decap_8 FILLER_25_1526 ();
 sg13g2_decap_8 FILLER_25_1533 ();
 sg13g2_decap_8 FILLER_25_1540 ();
 sg13g2_decap_8 FILLER_25_1547 ();
 sg13g2_decap_8 FILLER_25_1554 ();
 sg13g2_decap_8 FILLER_25_1561 ();
 sg13g2_decap_8 FILLER_25_1568 ();
 sg13g2_decap_8 FILLER_25_1575 ();
 sg13g2_decap_8 FILLER_25_1582 ();
 sg13g2_decap_8 FILLER_25_1589 ();
 sg13g2_decap_8 FILLER_25_1596 ();
 sg13g2_decap_8 FILLER_25_1603 ();
 sg13g2_decap_8 FILLER_25_1610 ();
 sg13g2_decap_8 FILLER_25_1617 ();
 sg13g2_decap_8 FILLER_25_1624 ();
 sg13g2_decap_8 FILLER_25_1631 ();
 sg13g2_decap_8 FILLER_25_1638 ();
 sg13g2_decap_8 FILLER_25_1645 ();
 sg13g2_decap_8 FILLER_25_1652 ();
 sg13g2_decap_8 FILLER_25_1659 ();
 sg13g2_decap_8 FILLER_25_1666 ();
 sg13g2_decap_8 FILLER_25_1673 ();
 sg13g2_decap_8 FILLER_25_1680 ();
 sg13g2_decap_8 FILLER_25_1687 ();
 sg13g2_decap_8 FILLER_25_1694 ();
 sg13g2_decap_8 FILLER_25_1701 ();
 sg13g2_decap_8 FILLER_25_1708 ();
 sg13g2_decap_8 FILLER_25_1715 ();
 sg13g2_decap_8 FILLER_25_1722 ();
 sg13g2_decap_8 FILLER_25_1729 ();
 sg13g2_decap_8 FILLER_25_1736 ();
 sg13g2_decap_8 FILLER_25_1743 ();
 sg13g2_decap_8 FILLER_25_1750 ();
 sg13g2_decap_8 FILLER_25_1757 ();
 sg13g2_decap_4 FILLER_25_1764 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_decap_8 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_decap_8 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_931 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_26_1029 ();
 sg13g2_decap_8 FILLER_26_1036 ();
 sg13g2_decap_8 FILLER_26_1043 ();
 sg13g2_decap_8 FILLER_26_1050 ();
 sg13g2_decap_8 FILLER_26_1057 ();
 sg13g2_decap_8 FILLER_26_1064 ();
 sg13g2_decap_8 FILLER_26_1071 ();
 sg13g2_decap_8 FILLER_26_1078 ();
 sg13g2_decap_8 FILLER_26_1085 ();
 sg13g2_decap_8 FILLER_26_1092 ();
 sg13g2_decap_8 FILLER_26_1099 ();
 sg13g2_decap_8 FILLER_26_1106 ();
 sg13g2_decap_8 FILLER_26_1113 ();
 sg13g2_decap_8 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1127 ();
 sg13g2_decap_8 FILLER_26_1134 ();
 sg13g2_decap_8 FILLER_26_1141 ();
 sg13g2_decap_8 FILLER_26_1148 ();
 sg13g2_decap_8 FILLER_26_1155 ();
 sg13g2_decap_8 FILLER_26_1162 ();
 sg13g2_decap_8 FILLER_26_1169 ();
 sg13g2_decap_8 FILLER_26_1176 ();
 sg13g2_decap_8 FILLER_26_1183 ();
 sg13g2_decap_8 FILLER_26_1190 ();
 sg13g2_decap_8 FILLER_26_1197 ();
 sg13g2_decap_8 FILLER_26_1204 ();
 sg13g2_decap_8 FILLER_26_1211 ();
 sg13g2_decap_8 FILLER_26_1218 ();
 sg13g2_decap_8 FILLER_26_1225 ();
 sg13g2_decap_8 FILLER_26_1232 ();
 sg13g2_decap_8 FILLER_26_1239 ();
 sg13g2_decap_8 FILLER_26_1246 ();
 sg13g2_decap_8 FILLER_26_1253 ();
 sg13g2_decap_8 FILLER_26_1260 ();
 sg13g2_decap_8 FILLER_26_1267 ();
 sg13g2_decap_8 FILLER_26_1274 ();
 sg13g2_decap_8 FILLER_26_1281 ();
 sg13g2_decap_8 FILLER_26_1288 ();
 sg13g2_decap_8 FILLER_26_1295 ();
 sg13g2_decap_8 FILLER_26_1302 ();
 sg13g2_decap_8 FILLER_26_1309 ();
 sg13g2_decap_8 FILLER_26_1316 ();
 sg13g2_decap_8 FILLER_26_1323 ();
 sg13g2_decap_8 FILLER_26_1330 ();
 sg13g2_decap_8 FILLER_26_1337 ();
 sg13g2_decap_8 FILLER_26_1344 ();
 sg13g2_decap_8 FILLER_26_1351 ();
 sg13g2_decap_8 FILLER_26_1358 ();
 sg13g2_decap_8 FILLER_26_1365 ();
 sg13g2_decap_8 FILLER_26_1372 ();
 sg13g2_decap_8 FILLER_26_1379 ();
 sg13g2_decap_8 FILLER_26_1386 ();
 sg13g2_decap_8 FILLER_26_1393 ();
 sg13g2_decap_8 FILLER_26_1400 ();
 sg13g2_decap_8 FILLER_26_1407 ();
 sg13g2_decap_8 FILLER_26_1414 ();
 sg13g2_decap_8 FILLER_26_1421 ();
 sg13g2_decap_8 FILLER_26_1428 ();
 sg13g2_decap_8 FILLER_26_1435 ();
 sg13g2_decap_8 FILLER_26_1442 ();
 sg13g2_decap_8 FILLER_26_1449 ();
 sg13g2_decap_8 FILLER_26_1456 ();
 sg13g2_decap_8 FILLER_26_1463 ();
 sg13g2_decap_8 FILLER_26_1470 ();
 sg13g2_decap_8 FILLER_26_1477 ();
 sg13g2_decap_8 FILLER_26_1484 ();
 sg13g2_decap_8 FILLER_26_1491 ();
 sg13g2_decap_8 FILLER_26_1498 ();
 sg13g2_decap_8 FILLER_26_1505 ();
 sg13g2_decap_8 FILLER_26_1512 ();
 sg13g2_decap_8 FILLER_26_1519 ();
 sg13g2_decap_8 FILLER_26_1526 ();
 sg13g2_decap_8 FILLER_26_1533 ();
 sg13g2_decap_8 FILLER_26_1540 ();
 sg13g2_decap_8 FILLER_26_1547 ();
 sg13g2_decap_8 FILLER_26_1554 ();
 sg13g2_decap_8 FILLER_26_1561 ();
 sg13g2_decap_8 FILLER_26_1568 ();
 sg13g2_decap_8 FILLER_26_1575 ();
 sg13g2_decap_8 FILLER_26_1582 ();
 sg13g2_decap_8 FILLER_26_1589 ();
 sg13g2_decap_8 FILLER_26_1596 ();
 sg13g2_decap_8 FILLER_26_1603 ();
 sg13g2_decap_8 FILLER_26_1610 ();
 sg13g2_decap_8 FILLER_26_1617 ();
 sg13g2_decap_8 FILLER_26_1624 ();
 sg13g2_decap_8 FILLER_26_1631 ();
 sg13g2_decap_8 FILLER_26_1638 ();
 sg13g2_decap_8 FILLER_26_1645 ();
 sg13g2_decap_8 FILLER_26_1652 ();
 sg13g2_decap_8 FILLER_26_1659 ();
 sg13g2_decap_8 FILLER_26_1666 ();
 sg13g2_decap_8 FILLER_26_1673 ();
 sg13g2_decap_8 FILLER_26_1680 ();
 sg13g2_decap_8 FILLER_26_1687 ();
 sg13g2_decap_8 FILLER_26_1694 ();
 sg13g2_decap_8 FILLER_26_1701 ();
 sg13g2_decap_8 FILLER_26_1708 ();
 sg13g2_decap_8 FILLER_26_1715 ();
 sg13g2_decap_8 FILLER_26_1722 ();
 sg13g2_decap_8 FILLER_26_1729 ();
 sg13g2_decap_8 FILLER_26_1736 ();
 sg13g2_decap_8 FILLER_26_1743 ();
 sg13g2_decap_8 FILLER_26_1750 ();
 sg13g2_decap_8 FILLER_26_1757 ();
 sg13g2_decap_4 FILLER_26_1764 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_decap_8 FILLER_27_1029 ();
 sg13g2_decap_8 FILLER_27_1036 ();
 sg13g2_decap_8 FILLER_27_1043 ();
 sg13g2_decap_8 FILLER_27_1050 ();
 sg13g2_decap_8 FILLER_27_1057 ();
 sg13g2_decap_8 FILLER_27_1064 ();
 sg13g2_decap_8 FILLER_27_1071 ();
 sg13g2_decap_8 FILLER_27_1078 ();
 sg13g2_decap_8 FILLER_27_1085 ();
 sg13g2_decap_8 FILLER_27_1092 ();
 sg13g2_decap_8 FILLER_27_1099 ();
 sg13g2_decap_8 FILLER_27_1106 ();
 sg13g2_decap_8 FILLER_27_1113 ();
 sg13g2_decap_8 FILLER_27_1120 ();
 sg13g2_decap_8 FILLER_27_1127 ();
 sg13g2_decap_8 FILLER_27_1134 ();
 sg13g2_decap_8 FILLER_27_1141 ();
 sg13g2_decap_8 FILLER_27_1148 ();
 sg13g2_decap_8 FILLER_27_1155 ();
 sg13g2_decap_8 FILLER_27_1162 ();
 sg13g2_decap_8 FILLER_27_1169 ();
 sg13g2_decap_8 FILLER_27_1176 ();
 sg13g2_decap_8 FILLER_27_1183 ();
 sg13g2_decap_8 FILLER_27_1190 ();
 sg13g2_decap_8 FILLER_27_1197 ();
 sg13g2_decap_8 FILLER_27_1204 ();
 sg13g2_decap_8 FILLER_27_1211 ();
 sg13g2_decap_8 FILLER_27_1218 ();
 sg13g2_decap_8 FILLER_27_1225 ();
 sg13g2_decap_8 FILLER_27_1232 ();
 sg13g2_decap_8 FILLER_27_1239 ();
 sg13g2_decap_8 FILLER_27_1246 ();
 sg13g2_decap_8 FILLER_27_1253 ();
 sg13g2_decap_8 FILLER_27_1260 ();
 sg13g2_decap_8 FILLER_27_1267 ();
 sg13g2_decap_8 FILLER_27_1274 ();
 sg13g2_decap_8 FILLER_27_1281 ();
 sg13g2_decap_8 FILLER_27_1288 ();
 sg13g2_decap_8 FILLER_27_1295 ();
 sg13g2_decap_8 FILLER_27_1302 ();
 sg13g2_decap_8 FILLER_27_1309 ();
 sg13g2_decap_8 FILLER_27_1316 ();
 sg13g2_decap_8 FILLER_27_1323 ();
 sg13g2_decap_8 FILLER_27_1330 ();
 sg13g2_decap_8 FILLER_27_1337 ();
 sg13g2_decap_8 FILLER_27_1344 ();
 sg13g2_decap_8 FILLER_27_1351 ();
 sg13g2_decap_8 FILLER_27_1358 ();
 sg13g2_decap_8 FILLER_27_1365 ();
 sg13g2_decap_8 FILLER_27_1372 ();
 sg13g2_decap_8 FILLER_27_1379 ();
 sg13g2_decap_8 FILLER_27_1386 ();
 sg13g2_decap_8 FILLER_27_1393 ();
 sg13g2_decap_8 FILLER_27_1400 ();
 sg13g2_decap_8 FILLER_27_1407 ();
 sg13g2_decap_8 FILLER_27_1414 ();
 sg13g2_decap_8 FILLER_27_1421 ();
 sg13g2_decap_8 FILLER_27_1428 ();
 sg13g2_decap_8 FILLER_27_1435 ();
 sg13g2_decap_8 FILLER_27_1442 ();
 sg13g2_decap_8 FILLER_27_1449 ();
 sg13g2_decap_8 FILLER_27_1456 ();
 sg13g2_decap_8 FILLER_27_1463 ();
 sg13g2_decap_8 FILLER_27_1470 ();
 sg13g2_decap_8 FILLER_27_1477 ();
 sg13g2_decap_8 FILLER_27_1484 ();
 sg13g2_decap_8 FILLER_27_1491 ();
 sg13g2_decap_8 FILLER_27_1498 ();
 sg13g2_decap_8 FILLER_27_1505 ();
 sg13g2_decap_8 FILLER_27_1512 ();
 sg13g2_decap_8 FILLER_27_1519 ();
 sg13g2_decap_8 FILLER_27_1526 ();
 sg13g2_decap_8 FILLER_27_1533 ();
 sg13g2_decap_8 FILLER_27_1540 ();
 sg13g2_decap_8 FILLER_27_1547 ();
 sg13g2_decap_8 FILLER_27_1554 ();
 sg13g2_decap_8 FILLER_27_1561 ();
 sg13g2_decap_8 FILLER_27_1568 ();
 sg13g2_decap_8 FILLER_27_1575 ();
 sg13g2_decap_8 FILLER_27_1582 ();
 sg13g2_decap_8 FILLER_27_1589 ();
 sg13g2_decap_8 FILLER_27_1596 ();
 sg13g2_decap_8 FILLER_27_1603 ();
 sg13g2_decap_8 FILLER_27_1610 ();
 sg13g2_decap_8 FILLER_27_1617 ();
 sg13g2_decap_8 FILLER_27_1624 ();
 sg13g2_decap_8 FILLER_27_1631 ();
 sg13g2_decap_8 FILLER_27_1638 ();
 sg13g2_decap_8 FILLER_27_1645 ();
 sg13g2_decap_8 FILLER_27_1652 ();
 sg13g2_decap_8 FILLER_27_1659 ();
 sg13g2_decap_8 FILLER_27_1666 ();
 sg13g2_decap_8 FILLER_27_1673 ();
 sg13g2_decap_8 FILLER_27_1680 ();
 sg13g2_decap_8 FILLER_27_1687 ();
 sg13g2_decap_8 FILLER_27_1694 ();
 sg13g2_decap_8 FILLER_27_1701 ();
 sg13g2_decap_8 FILLER_27_1708 ();
 sg13g2_decap_8 FILLER_27_1715 ();
 sg13g2_decap_8 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_27_1729 ();
 sg13g2_decap_8 FILLER_27_1736 ();
 sg13g2_decap_8 FILLER_27_1743 ();
 sg13g2_decap_8 FILLER_27_1750 ();
 sg13g2_decap_8 FILLER_27_1757 ();
 sg13g2_decap_4 FILLER_27_1764 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_decap_8 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_28_868 ();
 sg13g2_decap_8 FILLER_28_875 ();
 sg13g2_decap_8 FILLER_28_882 ();
 sg13g2_decap_8 FILLER_28_889 ();
 sg13g2_decap_8 FILLER_28_896 ();
 sg13g2_decap_8 FILLER_28_903 ();
 sg13g2_decap_8 FILLER_28_910 ();
 sg13g2_decap_8 FILLER_28_917 ();
 sg13g2_decap_8 FILLER_28_924 ();
 sg13g2_decap_8 FILLER_28_931 ();
 sg13g2_decap_8 FILLER_28_938 ();
 sg13g2_decap_8 FILLER_28_945 ();
 sg13g2_decap_8 FILLER_28_952 ();
 sg13g2_decap_8 FILLER_28_959 ();
 sg13g2_decap_8 FILLER_28_966 ();
 sg13g2_decap_8 FILLER_28_973 ();
 sg13g2_decap_8 FILLER_28_980 ();
 sg13g2_decap_8 FILLER_28_987 ();
 sg13g2_decap_8 FILLER_28_994 ();
 sg13g2_decap_8 FILLER_28_1001 ();
 sg13g2_decap_8 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1015 ();
 sg13g2_decap_8 FILLER_28_1022 ();
 sg13g2_decap_8 FILLER_28_1029 ();
 sg13g2_decap_8 FILLER_28_1036 ();
 sg13g2_decap_8 FILLER_28_1043 ();
 sg13g2_decap_8 FILLER_28_1050 ();
 sg13g2_decap_8 FILLER_28_1057 ();
 sg13g2_decap_8 FILLER_28_1064 ();
 sg13g2_decap_8 FILLER_28_1071 ();
 sg13g2_decap_8 FILLER_28_1078 ();
 sg13g2_decap_8 FILLER_28_1085 ();
 sg13g2_decap_8 FILLER_28_1092 ();
 sg13g2_decap_8 FILLER_28_1099 ();
 sg13g2_decap_8 FILLER_28_1106 ();
 sg13g2_decap_8 FILLER_28_1113 ();
 sg13g2_decap_8 FILLER_28_1120 ();
 sg13g2_decap_8 FILLER_28_1127 ();
 sg13g2_decap_8 FILLER_28_1134 ();
 sg13g2_decap_8 FILLER_28_1141 ();
 sg13g2_decap_8 FILLER_28_1148 ();
 sg13g2_decap_8 FILLER_28_1155 ();
 sg13g2_decap_8 FILLER_28_1162 ();
 sg13g2_decap_8 FILLER_28_1169 ();
 sg13g2_decap_8 FILLER_28_1176 ();
 sg13g2_decap_8 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1190 ();
 sg13g2_decap_8 FILLER_28_1197 ();
 sg13g2_decap_8 FILLER_28_1204 ();
 sg13g2_decap_8 FILLER_28_1211 ();
 sg13g2_decap_8 FILLER_28_1218 ();
 sg13g2_decap_8 FILLER_28_1225 ();
 sg13g2_decap_8 FILLER_28_1232 ();
 sg13g2_decap_8 FILLER_28_1239 ();
 sg13g2_decap_8 FILLER_28_1246 ();
 sg13g2_decap_8 FILLER_28_1253 ();
 sg13g2_decap_8 FILLER_28_1260 ();
 sg13g2_decap_8 FILLER_28_1267 ();
 sg13g2_decap_8 FILLER_28_1274 ();
 sg13g2_decap_8 FILLER_28_1281 ();
 sg13g2_decap_8 FILLER_28_1288 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1302 ();
 sg13g2_decap_8 FILLER_28_1309 ();
 sg13g2_decap_8 FILLER_28_1316 ();
 sg13g2_decap_8 FILLER_28_1323 ();
 sg13g2_decap_8 FILLER_28_1330 ();
 sg13g2_decap_8 FILLER_28_1337 ();
 sg13g2_decap_8 FILLER_28_1344 ();
 sg13g2_decap_8 FILLER_28_1351 ();
 sg13g2_decap_8 FILLER_28_1358 ();
 sg13g2_decap_8 FILLER_28_1365 ();
 sg13g2_decap_8 FILLER_28_1372 ();
 sg13g2_decap_8 FILLER_28_1379 ();
 sg13g2_decap_8 FILLER_28_1386 ();
 sg13g2_decap_8 FILLER_28_1393 ();
 sg13g2_decap_8 FILLER_28_1400 ();
 sg13g2_decap_8 FILLER_28_1407 ();
 sg13g2_decap_8 FILLER_28_1414 ();
 sg13g2_decap_8 FILLER_28_1421 ();
 sg13g2_decap_8 FILLER_28_1428 ();
 sg13g2_decap_8 FILLER_28_1435 ();
 sg13g2_decap_8 FILLER_28_1442 ();
 sg13g2_decap_8 FILLER_28_1449 ();
 sg13g2_decap_8 FILLER_28_1456 ();
 sg13g2_decap_8 FILLER_28_1463 ();
 sg13g2_decap_8 FILLER_28_1470 ();
 sg13g2_decap_8 FILLER_28_1477 ();
 sg13g2_decap_8 FILLER_28_1484 ();
 sg13g2_decap_8 FILLER_28_1491 ();
 sg13g2_decap_8 FILLER_28_1498 ();
 sg13g2_decap_8 FILLER_28_1505 ();
 sg13g2_decap_8 FILLER_28_1512 ();
 sg13g2_decap_8 FILLER_28_1519 ();
 sg13g2_decap_8 FILLER_28_1526 ();
 sg13g2_decap_8 FILLER_28_1533 ();
 sg13g2_decap_8 FILLER_28_1540 ();
 sg13g2_decap_8 FILLER_28_1547 ();
 sg13g2_decap_8 FILLER_28_1554 ();
 sg13g2_decap_8 FILLER_28_1561 ();
 sg13g2_decap_8 FILLER_28_1568 ();
 sg13g2_decap_8 FILLER_28_1575 ();
 sg13g2_decap_8 FILLER_28_1582 ();
 sg13g2_decap_8 FILLER_28_1589 ();
 sg13g2_decap_8 FILLER_28_1596 ();
 sg13g2_decap_8 FILLER_28_1603 ();
 sg13g2_decap_8 FILLER_28_1610 ();
 sg13g2_decap_8 FILLER_28_1617 ();
 sg13g2_decap_8 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_8 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1652 ();
 sg13g2_decap_8 FILLER_28_1659 ();
 sg13g2_decap_8 FILLER_28_1666 ();
 sg13g2_decap_8 FILLER_28_1673 ();
 sg13g2_decap_8 FILLER_28_1680 ();
 sg13g2_decap_8 FILLER_28_1687 ();
 sg13g2_decap_8 FILLER_28_1694 ();
 sg13g2_decap_8 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1708 ();
 sg13g2_decap_8 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1722 ();
 sg13g2_decap_8 FILLER_28_1729 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_8 FILLER_28_1757 ();
 sg13g2_decap_4 FILLER_28_1764 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_decap_8 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_882 ();
 sg13g2_decap_8 FILLER_29_889 ();
 sg13g2_decap_8 FILLER_29_896 ();
 sg13g2_decap_8 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_910 ();
 sg13g2_decap_8 FILLER_29_917 ();
 sg13g2_decap_8 FILLER_29_924 ();
 sg13g2_decap_8 FILLER_29_931 ();
 sg13g2_decap_8 FILLER_29_938 ();
 sg13g2_decap_8 FILLER_29_945 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_decap_8 FILLER_29_959 ();
 sg13g2_decap_8 FILLER_29_966 ();
 sg13g2_decap_8 FILLER_29_973 ();
 sg13g2_decap_8 FILLER_29_980 ();
 sg13g2_decap_8 FILLER_29_987 ();
 sg13g2_decap_8 FILLER_29_994 ();
 sg13g2_decap_8 FILLER_29_1001 ();
 sg13g2_decap_8 FILLER_29_1008 ();
 sg13g2_decap_8 FILLER_29_1015 ();
 sg13g2_decap_8 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_29_1029 ();
 sg13g2_decap_8 FILLER_29_1036 ();
 sg13g2_decap_8 FILLER_29_1043 ();
 sg13g2_decap_8 FILLER_29_1050 ();
 sg13g2_decap_8 FILLER_29_1057 ();
 sg13g2_decap_8 FILLER_29_1064 ();
 sg13g2_decap_8 FILLER_29_1071 ();
 sg13g2_decap_8 FILLER_29_1078 ();
 sg13g2_decap_8 FILLER_29_1085 ();
 sg13g2_decap_8 FILLER_29_1092 ();
 sg13g2_decap_8 FILLER_29_1099 ();
 sg13g2_decap_8 FILLER_29_1106 ();
 sg13g2_decap_8 FILLER_29_1113 ();
 sg13g2_decap_8 FILLER_29_1120 ();
 sg13g2_decap_8 FILLER_29_1127 ();
 sg13g2_decap_8 FILLER_29_1134 ();
 sg13g2_decap_8 FILLER_29_1141 ();
 sg13g2_decap_8 FILLER_29_1148 ();
 sg13g2_decap_8 FILLER_29_1155 ();
 sg13g2_decap_8 FILLER_29_1162 ();
 sg13g2_decap_8 FILLER_29_1169 ();
 sg13g2_decap_8 FILLER_29_1176 ();
 sg13g2_decap_8 FILLER_29_1183 ();
 sg13g2_decap_8 FILLER_29_1190 ();
 sg13g2_decap_8 FILLER_29_1197 ();
 sg13g2_decap_8 FILLER_29_1204 ();
 sg13g2_decap_8 FILLER_29_1211 ();
 sg13g2_decap_8 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1225 ();
 sg13g2_decap_8 FILLER_29_1232 ();
 sg13g2_decap_8 FILLER_29_1239 ();
 sg13g2_decap_8 FILLER_29_1246 ();
 sg13g2_decap_8 FILLER_29_1253 ();
 sg13g2_decap_8 FILLER_29_1260 ();
 sg13g2_decap_8 FILLER_29_1267 ();
 sg13g2_decap_8 FILLER_29_1274 ();
 sg13g2_decap_8 FILLER_29_1281 ();
 sg13g2_decap_8 FILLER_29_1288 ();
 sg13g2_decap_8 FILLER_29_1295 ();
 sg13g2_decap_8 FILLER_29_1302 ();
 sg13g2_decap_8 FILLER_29_1309 ();
 sg13g2_decap_8 FILLER_29_1316 ();
 sg13g2_decap_8 FILLER_29_1323 ();
 sg13g2_decap_8 FILLER_29_1330 ();
 sg13g2_decap_8 FILLER_29_1337 ();
 sg13g2_decap_8 FILLER_29_1344 ();
 sg13g2_decap_8 FILLER_29_1351 ();
 sg13g2_decap_8 FILLER_29_1358 ();
 sg13g2_decap_8 FILLER_29_1365 ();
 sg13g2_decap_8 FILLER_29_1372 ();
 sg13g2_decap_8 FILLER_29_1379 ();
 sg13g2_decap_8 FILLER_29_1386 ();
 sg13g2_decap_8 FILLER_29_1393 ();
 sg13g2_decap_8 FILLER_29_1400 ();
 sg13g2_decap_8 FILLER_29_1407 ();
 sg13g2_decap_8 FILLER_29_1414 ();
 sg13g2_decap_8 FILLER_29_1421 ();
 sg13g2_decap_8 FILLER_29_1428 ();
 sg13g2_decap_8 FILLER_29_1435 ();
 sg13g2_decap_8 FILLER_29_1442 ();
 sg13g2_decap_8 FILLER_29_1449 ();
 sg13g2_decap_8 FILLER_29_1456 ();
 sg13g2_decap_8 FILLER_29_1463 ();
 sg13g2_decap_8 FILLER_29_1470 ();
 sg13g2_decap_8 FILLER_29_1477 ();
 sg13g2_decap_8 FILLER_29_1484 ();
 sg13g2_decap_8 FILLER_29_1491 ();
 sg13g2_decap_8 FILLER_29_1498 ();
 sg13g2_decap_8 FILLER_29_1505 ();
 sg13g2_decap_8 FILLER_29_1512 ();
 sg13g2_decap_8 FILLER_29_1519 ();
 sg13g2_decap_8 FILLER_29_1526 ();
 sg13g2_decap_8 FILLER_29_1533 ();
 sg13g2_decap_8 FILLER_29_1540 ();
 sg13g2_decap_8 FILLER_29_1547 ();
 sg13g2_decap_8 FILLER_29_1554 ();
 sg13g2_decap_8 FILLER_29_1561 ();
 sg13g2_decap_8 FILLER_29_1568 ();
 sg13g2_decap_8 FILLER_29_1575 ();
 sg13g2_decap_8 FILLER_29_1582 ();
 sg13g2_decap_8 FILLER_29_1589 ();
 sg13g2_decap_8 FILLER_29_1596 ();
 sg13g2_decap_8 FILLER_29_1603 ();
 sg13g2_decap_8 FILLER_29_1610 ();
 sg13g2_decap_8 FILLER_29_1617 ();
 sg13g2_decap_8 FILLER_29_1624 ();
 sg13g2_decap_8 FILLER_29_1631 ();
 sg13g2_decap_8 FILLER_29_1638 ();
 sg13g2_decap_8 FILLER_29_1645 ();
 sg13g2_decap_8 FILLER_29_1652 ();
 sg13g2_decap_8 FILLER_29_1659 ();
 sg13g2_decap_8 FILLER_29_1666 ();
 sg13g2_decap_8 FILLER_29_1673 ();
 sg13g2_decap_8 FILLER_29_1680 ();
 sg13g2_decap_8 FILLER_29_1687 ();
 sg13g2_decap_8 FILLER_29_1694 ();
 sg13g2_decap_8 FILLER_29_1701 ();
 sg13g2_decap_8 FILLER_29_1708 ();
 sg13g2_decap_8 FILLER_29_1715 ();
 sg13g2_decap_8 FILLER_29_1722 ();
 sg13g2_decap_8 FILLER_29_1729 ();
 sg13g2_decap_8 FILLER_29_1736 ();
 sg13g2_decap_8 FILLER_29_1743 ();
 sg13g2_decap_8 FILLER_29_1750 ();
 sg13g2_decap_8 FILLER_29_1757 ();
 sg13g2_decap_4 FILLER_29_1764 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_decap_8 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_30_1029 ();
 sg13g2_decap_8 FILLER_30_1036 ();
 sg13g2_decap_8 FILLER_30_1043 ();
 sg13g2_decap_8 FILLER_30_1050 ();
 sg13g2_decap_8 FILLER_30_1057 ();
 sg13g2_decap_8 FILLER_30_1064 ();
 sg13g2_decap_8 FILLER_30_1071 ();
 sg13g2_decap_8 FILLER_30_1078 ();
 sg13g2_decap_8 FILLER_30_1085 ();
 sg13g2_decap_8 FILLER_30_1092 ();
 sg13g2_decap_8 FILLER_30_1099 ();
 sg13g2_decap_8 FILLER_30_1106 ();
 sg13g2_decap_8 FILLER_30_1113 ();
 sg13g2_decap_8 FILLER_30_1120 ();
 sg13g2_decap_8 FILLER_30_1127 ();
 sg13g2_decap_8 FILLER_30_1134 ();
 sg13g2_decap_8 FILLER_30_1141 ();
 sg13g2_decap_8 FILLER_30_1148 ();
 sg13g2_decap_8 FILLER_30_1155 ();
 sg13g2_decap_8 FILLER_30_1162 ();
 sg13g2_decap_8 FILLER_30_1169 ();
 sg13g2_decap_8 FILLER_30_1176 ();
 sg13g2_decap_8 FILLER_30_1183 ();
 sg13g2_decap_8 FILLER_30_1190 ();
 sg13g2_decap_8 FILLER_30_1197 ();
 sg13g2_decap_8 FILLER_30_1204 ();
 sg13g2_decap_8 FILLER_30_1211 ();
 sg13g2_decap_8 FILLER_30_1218 ();
 sg13g2_decap_8 FILLER_30_1225 ();
 sg13g2_decap_8 FILLER_30_1232 ();
 sg13g2_decap_8 FILLER_30_1239 ();
 sg13g2_decap_8 FILLER_30_1246 ();
 sg13g2_decap_8 FILLER_30_1253 ();
 sg13g2_decap_8 FILLER_30_1260 ();
 sg13g2_decap_8 FILLER_30_1267 ();
 sg13g2_decap_8 FILLER_30_1274 ();
 sg13g2_decap_8 FILLER_30_1281 ();
 sg13g2_decap_8 FILLER_30_1288 ();
 sg13g2_decap_8 FILLER_30_1295 ();
 sg13g2_decap_8 FILLER_30_1302 ();
 sg13g2_decap_8 FILLER_30_1309 ();
 sg13g2_decap_8 FILLER_30_1316 ();
 sg13g2_decap_8 FILLER_30_1323 ();
 sg13g2_decap_8 FILLER_30_1330 ();
 sg13g2_decap_8 FILLER_30_1337 ();
 sg13g2_decap_8 FILLER_30_1344 ();
 sg13g2_decap_8 FILLER_30_1351 ();
 sg13g2_decap_8 FILLER_30_1358 ();
 sg13g2_decap_8 FILLER_30_1365 ();
 sg13g2_decap_8 FILLER_30_1372 ();
 sg13g2_decap_8 FILLER_30_1379 ();
 sg13g2_decap_8 FILLER_30_1386 ();
 sg13g2_decap_8 FILLER_30_1393 ();
 sg13g2_decap_8 FILLER_30_1400 ();
 sg13g2_decap_8 FILLER_30_1407 ();
 sg13g2_decap_8 FILLER_30_1414 ();
 sg13g2_decap_8 FILLER_30_1421 ();
 sg13g2_decap_8 FILLER_30_1428 ();
 sg13g2_decap_8 FILLER_30_1435 ();
 sg13g2_decap_8 FILLER_30_1442 ();
 sg13g2_decap_8 FILLER_30_1449 ();
 sg13g2_decap_8 FILLER_30_1456 ();
 sg13g2_decap_8 FILLER_30_1463 ();
 sg13g2_decap_8 FILLER_30_1470 ();
 sg13g2_decap_8 FILLER_30_1477 ();
 sg13g2_decap_8 FILLER_30_1484 ();
 sg13g2_decap_8 FILLER_30_1491 ();
 sg13g2_decap_8 FILLER_30_1498 ();
 sg13g2_decap_8 FILLER_30_1505 ();
 sg13g2_decap_8 FILLER_30_1512 ();
 sg13g2_decap_8 FILLER_30_1519 ();
 sg13g2_decap_8 FILLER_30_1526 ();
 sg13g2_decap_8 FILLER_30_1533 ();
 sg13g2_decap_8 FILLER_30_1540 ();
 sg13g2_decap_8 FILLER_30_1547 ();
 sg13g2_decap_8 FILLER_30_1554 ();
 sg13g2_decap_8 FILLER_30_1561 ();
 sg13g2_decap_8 FILLER_30_1568 ();
 sg13g2_decap_8 FILLER_30_1575 ();
 sg13g2_decap_8 FILLER_30_1582 ();
 sg13g2_decap_8 FILLER_30_1589 ();
 sg13g2_decap_8 FILLER_30_1596 ();
 sg13g2_decap_8 FILLER_30_1603 ();
 sg13g2_decap_8 FILLER_30_1610 ();
 sg13g2_decap_8 FILLER_30_1617 ();
 sg13g2_decap_8 FILLER_30_1624 ();
 sg13g2_decap_8 FILLER_30_1631 ();
 sg13g2_decap_8 FILLER_30_1638 ();
 sg13g2_decap_8 FILLER_30_1645 ();
 sg13g2_decap_8 FILLER_30_1652 ();
 sg13g2_decap_8 FILLER_30_1659 ();
 sg13g2_decap_8 FILLER_30_1666 ();
 sg13g2_decap_8 FILLER_30_1673 ();
 sg13g2_decap_8 FILLER_30_1680 ();
 sg13g2_decap_8 FILLER_30_1687 ();
 sg13g2_decap_8 FILLER_30_1694 ();
 sg13g2_decap_8 FILLER_30_1701 ();
 sg13g2_decap_8 FILLER_30_1708 ();
 sg13g2_decap_8 FILLER_30_1715 ();
 sg13g2_decap_8 FILLER_30_1722 ();
 sg13g2_decap_8 FILLER_30_1729 ();
 sg13g2_decap_8 FILLER_30_1736 ();
 sg13g2_decap_8 FILLER_30_1743 ();
 sg13g2_decap_8 FILLER_30_1750 ();
 sg13g2_decap_8 FILLER_30_1757 ();
 sg13g2_decap_4 FILLER_30_1764 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_31_1029 ();
 sg13g2_decap_8 FILLER_31_1036 ();
 sg13g2_decap_8 FILLER_31_1043 ();
 sg13g2_decap_8 FILLER_31_1050 ();
 sg13g2_decap_8 FILLER_31_1057 ();
 sg13g2_decap_8 FILLER_31_1064 ();
 sg13g2_decap_8 FILLER_31_1071 ();
 sg13g2_decap_8 FILLER_31_1078 ();
 sg13g2_decap_8 FILLER_31_1085 ();
 sg13g2_decap_8 FILLER_31_1092 ();
 sg13g2_decap_8 FILLER_31_1099 ();
 sg13g2_decap_8 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1113 ();
 sg13g2_decap_8 FILLER_31_1120 ();
 sg13g2_decap_8 FILLER_31_1127 ();
 sg13g2_decap_8 FILLER_31_1134 ();
 sg13g2_decap_8 FILLER_31_1141 ();
 sg13g2_decap_8 FILLER_31_1148 ();
 sg13g2_decap_8 FILLER_31_1155 ();
 sg13g2_decap_8 FILLER_31_1162 ();
 sg13g2_decap_8 FILLER_31_1169 ();
 sg13g2_decap_8 FILLER_31_1176 ();
 sg13g2_decap_8 FILLER_31_1183 ();
 sg13g2_decap_8 FILLER_31_1190 ();
 sg13g2_decap_8 FILLER_31_1197 ();
 sg13g2_decap_8 FILLER_31_1204 ();
 sg13g2_decap_8 FILLER_31_1211 ();
 sg13g2_decap_8 FILLER_31_1218 ();
 sg13g2_decap_8 FILLER_31_1225 ();
 sg13g2_decap_8 FILLER_31_1232 ();
 sg13g2_decap_8 FILLER_31_1239 ();
 sg13g2_decap_8 FILLER_31_1246 ();
 sg13g2_decap_8 FILLER_31_1253 ();
 sg13g2_decap_8 FILLER_31_1260 ();
 sg13g2_decap_8 FILLER_31_1267 ();
 sg13g2_decap_8 FILLER_31_1274 ();
 sg13g2_decap_8 FILLER_31_1281 ();
 sg13g2_decap_8 FILLER_31_1288 ();
 sg13g2_decap_8 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1302 ();
 sg13g2_decap_8 FILLER_31_1309 ();
 sg13g2_decap_8 FILLER_31_1316 ();
 sg13g2_decap_8 FILLER_31_1323 ();
 sg13g2_decap_8 FILLER_31_1330 ();
 sg13g2_decap_8 FILLER_31_1337 ();
 sg13g2_decap_8 FILLER_31_1344 ();
 sg13g2_decap_8 FILLER_31_1351 ();
 sg13g2_decap_8 FILLER_31_1358 ();
 sg13g2_decap_8 FILLER_31_1365 ();
 sg13g2_decap_8 FILLER_31_1372 ();
 sg13g2_decap_8 FILLER_31_1379 ();
 sg13g2_decap_8 FILLER_31_1386 ();
 sg13g2_decap_8 FILLER_31_1393 ();
 sg13g2_decap_8 FILLER_31_1400 ();
 sg13g2_decap_8 FILLER_31_1407 ();
 sg13g2_decap_8 FILLER_31_1414 ();
 sg13g2_decap_8 FILLER_31_1421 ();
 sg13g2_decap_8 FILLER_31_1428 ();
 sg13g2_decap_8 FILLER_31_1435 ();
 sg13g2_decap_8 FILLER_31_1442 ();
 sg13g2_decap_8 FILLER_31_1449 ();
 sg13g2_decap_8 FILLER_31_1456 ();
 sg13g2_decap_8 FILLER_31_1463 ();
 sg13g2_decap_8 FILLER_31_1470 ();
 sg13g2_decap_8 FILLER_31_1477 ();
 sg13g2_decap_8 FILLER_31_1484 ();
 sg13g2_decap_8 FILLER_31_1491 ();
 sg13g2_decap_8 FILLER_31_1498 ();
 sg13g2_decap_8 FILLER_31_1505 ();
 sg13g2_decap_8 FILLER_31_1512 ();
 sg13g2_decap_8 FILLER_31_1519 ();
 sg13g2_decap_8 FILLER_31_1526 ();
 sg13g2_decap_8 FILLER_31_1533 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_decap_8 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1568 ();
 sg13g2_decap_8 FILLER_31_1575 ();
 sg13g2_decap_8 FILLER_31_1582 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_decap_8 FILLER_31_1603 ();
 sg13g2_decap_8 FILLER_31_1610 ();
 sg13g2_decap_8 FILLER_31_1617 ();
 sg13g2_decap_8 FILLER_31_1624 ();
 sg13g2_decap_8 FILLER_31_1631 ();
 sg13g2_decap_8 FILLER_31_1638 ();
 sg13g2_decap_8 FILLER_31_1645 ();
 sg13g2_decap_8 FILLER_31_1652 ();
 sg13g2_decap_8 FILLER_31_1659 ();
 sg13g2_decap_8 FILLER_31_1666 ();
 sg13g2_decap_8 FILLER_31_1673 ();
 sg13g2_decap_8 FILLER_31_1680 ();
 sg13g2_decap_8 FILLER_31_1687 ();
 sg13g2_decap_8 FILLER_31_1694 ();
 sg13g2_decap_8 FILLER_31_1701 ();
 sg13g2_decap_8 FILLER_31_1708 ();
 sg13g2_decap_8 FILLER_31_1715 ();
 sg13g2_decap_8 FILLER_31_1722 ();
 sg13g2_decap_8 FILLER_31_1729 ();
 sg13g2_decap_8 FILLER_31_1736 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_4 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_decap_8 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_32_847 ();
 sg13g2_decap_8 FILLER_32_854 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_882 ();
 sg13g2_decap_8 FILLER_32_889 ();
 sg13g2_decap_8 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_903 ();
 sg13g2_decap_8 FILLER_32_910 ();
 sg13g2_decap_8 FILLER_32_917 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_8 FILLER_32_931 ();
 sg13g2_decap_8 FILLER_32_938 ();
 sg13g2_decap_8 FILLER_32_945 ();
 sg13g2_decap_8 FILLER_32_952 ();
 sg13g2_decap_8 FILLER_32_959 ();
 sg13g2_decap_8 FILLER_32_966 ();
 sg13g2_decap_8 FILLER_32_973 ();
 sg13g2_decap_8 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_987 ();
 sg13g2_decap_8 FILLER_32_994 ();
 sg13g2_decap_8 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1008 ();
 sg13g2_decap_8 FILLER_32_1015 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_32_1029 ();
 sg13g2_decap_8 FILLER_32_1036 ();
 sg13g2_decap_8 FILLER_32_1043 ();
 sg13g2_decap_8 FILLER_32_1050 ();
 sg13g2_decap_8 FILLER_32_1057 ();
 sg13g2_decap_8 FILLER_32_1064 ();
 sg13g2_decap_8 FILLER_32_1071 ();
 sg13g2_decap_8 FILLER_32_1078 ();
 sg13g2_decap_8 FILLER_32_1085 ();
 sg13g2_decap_8 FILLER_32_1092 ();
 sg13g2_decap_8 FILLER_32_1099 ();
 sg13g2_decap_8 FILLER_32_1106 ();
 sg13g2_decap_8 FILLER_32_1113 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_8 FILLER_32_1169 ();
 sg13g2_decap_8 FILLER_32_1176 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1204 ();
 sg13g2_decap_8 FILLER_32_1211 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_decap_8 FILLER_32_1246 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_8 FILLER_32_1309 ();
 sg13g2_decap_8 FILLER_32_1316 ();
 sg13g2_decap_8 FILLER_32_1323 ();
 sg13g2_decap_8 FILLER_32_1330 ();
 sg13g2_decap_8 FILLER_32_1337 ();
 sg13g2_decap_8 FILLER_32_1344 ();
 sg13g2_decap_8 FILLER_32_1351 ();
 sg13g2_decap_8 FILLER_32_1358 ();
 sg13g2_decap_8 FILLER_32_1365 ();
 sg13g2_decap_8 FILLER_32_1372 ();
 sg13g2_decap_8 FILLER_32_1379 ();
 sg13g2_decap_8 FILLER_32_1386 ();
 sg13g2_decap_8 FILLER_32_1393 ();
 sg13g2_decap_8 FILLER_32_1400 ();
 sg13g2_decap_8 FILLER_32_1407 ();
 sg13g2_decap_8 FILLER_32_1414 ();
 sg13g2_decap_8 FILLER_32_1421 ();
 sg13g2_decap_8 FILLER_32_1428 ();
 sg13g2_decap_8 FILLER_32_1435 ();
 sg13g2_decap_8 FILLER_32_1442 ();
 sg13g2_decap_8 FILLER_32_1449 ();
 sg13g2_decap_8 FILLER_32_1456 ();
 sg13g2_decap_8 FILLER_32_1463 ();
 sg13g2_decap_8 FILLER_32_1470 ();
 sg13g2_decap_8 FILLER_32_1477 ();
 sg13g2_decap_8 FILLER_32_1484 ();
 sg13g2_decap_8 FILLER_32_1491 ();
 sg13g2_decap_8 FILLER_32_1498 ();
 sg13g2_decap_8 FILLER_32_1505 ();
 sg13g2_decap_8 FILLER_32_1512 ();
 sg13g2_decap_8 FILLER_32_1519 ();
 sg13g2_decap_8 FILLER_32_1526 ();
 sg13g2_decap_8 FILLER_32_1533 ();
 sg13g2_decap_8 FILLER_32_1540 ();
 sg13g2_decap_8 FILLER_32_1547 ();
 sg13g2_decap_8 FILLER_32_1554 ();
 sg13g2_decap_8 FILLER_32_1561 ();
 sg13g2_decap_8 FILLER_32_1568 ();
 sg13g2_decap_8 FILLER_32_1575 ();
 sg13g2_decap_8 FILLER_32_1582 ();
 sg13g2_decap_8 FILLER_32_1589 ();
 sg13g2_decap_8 FILLER_32_1596 ();
 sg13g2_decap_8 FILLER_32_1603 ();
 sg13g2_decap_8 FILLER_32_1610 ();
 sg13g2_decap_8 FILLER_32_1617 ();
 sg13g2_decap_8 FILLER_32_1624 ();
 sg13g2_decap_8 FILLER_32_1631 ();
 sg13g2_decap_8 FILLER_32_1638 ();
 sg13g2_decap_8 FILLER_32_1645 ();
 sg13g2_decap_8 FILLER_32_1652 ();
 sg13g2_decap_8 FILLER_32_1659 ();
 sg13g2_decap_8 FILLER_32_1666 ();
 sg13g2_decap_8 FILLER_32_1673 ();
 sg13g2_decap_8 FILLER_32_1680 ();
 sg13g2_decap_8 FILLER_32_1687 ();
 sg13g2_decap_8 FILLER_32_1694 ();
 sg13g2_decap_8 FILLER_32_1701 ();
 sg13g2_decap_8 FILLER_32_1708 ();
 sg13g2_decap_8 FILLER_32_1715 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_8 FILLER_32_1729 ();
 sg13g2_decap_8 FILLER_32_1736 ();
 sg13g2_decap_8 FILLER_32_1743 ();
 sg13g2_decap_8 FILLER_32_1750 ();
 sg13g2_decap_8 FILLER_32_1757 ();
 sg13g2_decap_4 FILLER_32_1764 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_33_1029 ();
 sg13g2_decap_8 FILLER_33_1036 ();
 sg13g2_decap_8 FILLER_33_1043 ();
 sg13g2_decap_8 FILLER_33_1050 ();
 sg13g2_decap_8 FILLER_33_1057 ();
 sg13g2_decap_8 FILLER_33_1064 ();
 sg13g2_decap_8 FILLER_33_1071 ();
 sg13g2_decap_8 FILLER_33_1078 ();
 sg13g2_decap_8 FILLER_33_1085 ();
 sg13g2_decap_8 FILLER_33_1092 ();
 sg13g2_decap_8 FILLER_33_1099 ();
 sg13g2_decap_8 FILLER_33_1106 ();
 sg13g2_decap_8 FILLER_33_1113 ();
 sg13g2_decap_8 FILLER_33_1120 ();
 sg13g2_decap_8 FILLER_33_1127 ();
 sg13g2_decap_8 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1141 ();
 sg13g2_decap_8 FILLER_33_1148 ();
 sg13g2_decap_8 FILLER_33_1155 ();
 sg13g2_decap_8 FILLER_33_1162 ();
 sg13g2_decap_8 FILLER_33_1169 ();
 sg13g2_decap_8 FILLER_33_1176 ();
 sg13g2_decap_8 FILLER_33_1183 ();
 sg13g2_decap_8 FILLER_33_1190 ();
 sg13g2_decap_8 FILLER_33_1197 ();
 sg13g2_decap_8 FILLER_33_1204 ();
 sg13g2_decap_8 FILLER_33_1211 ();
 sg13g2_decap_8 FILLER_33_1218 ();
 sg13g2_decap_8 FILLER_33_1225 ();
 sg13g2_decap_8 FILLER_33_1232 ();
 sg13g2_decap_8 FILLER_33_1239 ();
 sg13g2_decap_8 FILLER_33_1246 ();
 sg13g2_decap_8 FILLER_33_1253 ();
 sg13g2_decap_8 FILLER_33_1260 ();
 sg13g2_decap_8 FILLER_33_1267 ();
 sg13g2_decap_8 FILLER_33_1274 ();
 sg13g2_decap_8 FILLER_33_1281 ();
 sg13g2_decap_8 FILLER_33_1288 ();
 sg13g2_decap_8 FILLER_33_1295 ();
 sg13g2_decap_8 FILLER_33_1302 ();
 sg13g2_decap_8 FILLER_33_1309 ();
 sg13g2_decap_8 FILLER_33_1316 ();
 sg13g2_decap_8 FILLER_33_1323 ();
 sg13g2_decap_8 FILLER_33_1330 ();
 sg13g2_decap_8 FILLER_33_1337 ();
 sg13g2_decap_8 FILLER_33_1344 ();
 sg13g2_decap_8 FILLER_33_1351 ();
 sg13g2_decap_8 FILLER_33_1358 ();
 sg13g2_decap_8 FILLER_33_1365 ();
 sg13g2_decap_8 FILLER_33_1372 ();
 sg13g2_decap_8 FILLER_33_1379 ();
 sg13g2_decap_8 FILLER_33_1386 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_8 FILLER_33_1400 ();
 sg13g2_decap_8 FILLER_33_1407 ();
 sg13g2_decap_8 FILLER_33_1414 ();
 sg13g2_decap_8 FILLER_33_1421 ();
 sg13g2_decap_8 FILLER_33_1428 ();
 sg13g2_decap_8 FILLER_33_1435 ();
 sg13g2_decap_8 FILLER_33_1442 ();
 sg13g2_decap_8 FILLER_33_1449 ();
 sg13g2_decap_8 FILLER_33_1456 ();
 sg13g2_decap_8 FILLER_33_1463 ();
 sg13g2_decap_8 FILLER_33_1470 ();
 sg13g2_decap_8 FILLER_33_1477 ();
 sg13g2_decap_8 FILLER_33_1484 ();
 sg13g2_decap_8 FILLER_33_1491 ();
 sg13g2_decap_8 FILLER_33_1498 ();
 sg13g2_decap_8 FILLER_33_1505 ();
 sg13g2_decap_8 FILLER_33_1512 ();
 sg13g2_decap_8 FILLER_33_1519 ();
 sg13g2_decap_8 FILLER_33_1526 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_decap_8 FILLER_33_1540 ();
 sg13g2_decap_8 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1554 ();
 sg13g2_decap_8 FILLER_33_1561 ();
 sg13g2_decap_8 FILLER_33_1568 ();
 sg13g2_decap_8 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1582 ();
 sg13g2_decap_8 FILLER_33_1589 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1603 ();
 sg13g2_decap_8 FILLER_33_1610 ();
 sg13g2_decap_8 FILLER_33_1617 ();
 sg13g2_decap_8 FILLER_33_1624 ();
 sg13g2_decap_8 FILLER_33_1631 ();
 sg13g2_decap_8 FILLER_33_1638 ();
 sg13g2_decap_8 FILLER_33_1645 ();
 sg13g2_decap_8 FILLER_33_1652 ();
 sg13g2_decap_8 FILLER_33_1659 ();
 sg13g2_decap_8 FILLER_33_1666 ();
 sg13g2_decap_8 FILLER_33_1673 ();
 sg13g2_decap_8 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1687 ();
 sg13g2_decap_8 FILLER_33_1694 ();
 sg13g2_decap_8 FILLER_33_1701 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_8 FILLER_33_1722 ();
 sg13g2_decap_8 FILLER_33_1729 ();
 sg13g2_decap_8 FILLER_33_1736 ();
 sg13g2_decap_8 FILLER_33_1743 ();
 sg13g2_decap_8 FILLER_33_1750 ();
 sg13g2_decap_8 FILLER_33_1757 ();
 sg13g2_decap_4 FILLER_33_1764 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_34_847 ();
 sg13g2_decap_8 FILLER_34_854 ();
 sg13g2_decap_8 FILLER_34_861 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_decap_8 FILLER_34_896 ();
 sg13g2_decap_8 FILLER_34_903 ();
 sg13g2_decap_8 FILLER_34_910 ();
 sg13g2_decap_8 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_34_1029 ();
 sg13g2_decap_8 FILLER_34_1036 ();
 sg13g2_decap_8 FILLER_34_1043 ();
 sg13g2_decap_8 FILLER_34_1050 ();
 sg13g2_decap_8 FILLER_34_1057 ();
 sg13g2_decap_8 FILLER_34_1064 ();
 sg13g2_decap_8 FILLER_34_1071 ();
 sg13g2_decap_8 FILLER_34_1078 ();
 sg13g2_decap_8 FILLER_34_1085 ();
 sg13g2_decap_8 FILLER_34_1092 ();
 sg13g2_decap_8 FILLER_34_1099 ();
 sg13g2_decap_8 FILLER_34_1106 ();
 sg13g2_decap_8 FILLER_34_1113 ();
 sg13g2_decap_8 FILLER_34_1120 ();
 sg13g2_decap_8 FILLER_34_1127 ();
 sg13g2_decap_8 FILLER_34_1134 ();
 sg13g2_decap_8 FILLER_34_1141 ();
 sg13g2_decap_8 FILLER_34_1148 ();
 sg13g2_decap_8 FILLER_34_1155 ();
 sg13g2_decap_8 FILLER_34_1162 ();
 sg13g2_decap_8 FILLER_34_1169 ();
 sg13g2_decap_8 FILLER_34_1176 ();
 sg13g2_decap_8 FILLER_34_1183 ();
 sg13g2_decap_8 FILLER_34_1190 ();
 sg13g2_decap_8 FILLER_34_1197 ();
 sg13g2_decap_8 FILLER_34_1204 ();
 sg13g2_decap_8 FILLER_34_1211 ();
 sg13g2_decap_8 FILLER_34_1218 ();
 sg13g2_decap_8 FILLER_34_1225 ();
 sg13g2_decap_8 FILLER_34_1232 ();
 sg13g2_decap_8 FILLER_34_1239 ();
 sg13g2_decap_8 FILLER_34_1246 ();
 sg13g2_decap_8 FILLER_34_1253 ();
 sg13g2_decap_8 FILLER_34_1260 ();
 sg13g2_decap_8 FILLER_34_1267 ();
 sg13g2_decap_8 FILLER_34_1274 ();
 sg13g2_decap_8 FILLER_34_1281 ();
 sg13g2_decap_8 FILLER_34_1288 ();
 sg13g2_decap_8 FILLER_34_1295 ();
 sg13g2_decap_8 FILLER_34_1302 ();
 sg13g2_decap_8 FILLER_34_1309 ();
 sg13g2_decap_8 FILLER_34_1316 ();
 sg13g2_decap_8 FILLER_34_1323 ();
 sg13g2_decap_8 FILLER_34_1330 ();
 sg13g2_decap_8 FILLER_34_1337 ();
 sg13g2_decap_8 FILLER_34_1344 ();
 sg13g2_decap_8 FILLER_34_1351 ();
 sg13g2_decap_8 FILLER_34_1358 ();
 sg13g2_decap_8 FILLER_34_1365 ();
 sg13g2_decap_8 FILLER_34_1372 ();
 sg13g2_decap_8 FILLER_34_1379 ();
 sg13g2_decap_8 FILLER_34_1386 ();
 sg13g2_decap_8 FILLER_34_1393 ();
 sg13g2_decap_8 FILLER_34_1400 ();
 sg13g2_decap_8 FILLER_34_1407 ();
 sg13g2_decap_8 FILLER_34_1414 ();
 sg13g2_decap_8 FILLER_34_1421 ();
 sg13g2_decap_8 FILLER_34_1428 ();
 sg13g2_decap_8 FILLER_34_1435 ();
 sg13g2_decap_8 FILLER_34_1442 ();
 sg13g2_decap_8 FILLER_34_1449 ();
 sg13g2_decap_8 FILLER_34_1456 ();
 sg13g2_decap_8 FILLER_34_1463 ();
 sg13g2_decap_8 FILLER_34_1470 ();
 sg13g2_decap_8 FILLER_34_1477 ();
 sg13g2_decap_8 FILLER_34_1484 ();
 sg13g2_decap_8 FILLER_34_1491 ();
 sg13g2_decap_8 FILLER_34_1498 ();
 sg13g2_decap_8 FILLER_34_1505 ();
 sg13g2_decap_8 FILLER_34_1512 ();
 sg13g2_decap_8 FILLER_34_1519 ();
 sg13g2_decap_8 FILLER_34_1526 ();
 sg13g2_decap_8 FILLER_34_1533 ();
 sg13g2_decap_8 FILLER_34_1540 ();
 sg13g2_decap_8 FILLER_34_1547 ();
 sg13g2_decap_8 FILLER_34_1554 ();
 sg13g2_decap_8 FILLER_34_1561 ();
 sg13g2_decap_8 FILLER_34_1568 ();
 sg13g2_decap_8 FILLER_34_1575 ();
 sg13g2_decap_8 FILLER_34_1582 ();
 sg13g2_decap_8 FILLER_34_1589 ();
 sg13g2_decap_8 FILLER_34_1596 ();
 sg13g2_decap_8 FILLER_34_1603 ();
 sg13g2_decap_8 FILLER_34_1610 ();
 sg13g2_decap_8 FILLER_34_1617 ();
 sg13g2_decap_8 FILLER_34_1624 ();
 sg13g2_decap_8 FILLER_34_1631 ();
 sg13g2_decap_8 FILLER_34_1638 ();
 sg13g2_decap_8 FILLER_34_1645 ();
 sg13g2_decap_8 FILLER_34_1652 ();
 sg13g2_decap_8 FILLER_34_1659 ();
 sg13g2_decap_8 FILLER_34_1666 ();
 sg13g2_decap_8 FILLER_34_1673 ();
 sg13g2_decap_8 FILLER_34_1680 ();
 sg13g2_decap_8 FILLER_34_1687 ();
 sg13g2_decap_8 FILLER_34_1694 ();
 sg13g2_decap_8 FILLER_34_1701 ();
 sg13g2_decap_8 FILLER_34_1708 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_8 FILLER_34_1729 ();
 sg13g2_decap_8 FILLER_34_1736 ();
 sg13g2_decap_8 FILLER_34_1743 ();
 sg13g2_decap_8 FILLER_34_1750 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_4 FILLER_34_1764 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_decap_8 FILLER_35_875 ();
 sg13g2_decap_8 FILLER_35_882 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_decap_8 FILLER_35_896 ();
 sg13g2_decap_8 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_910 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_945 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_8 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_973 ();
 sg13g2_decap_8 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_8 FILLER_35_994 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_decap_8 FILLER_35_1043 ();
 sg13g2_decap_8 FILLER_35_1050 ();
 sg13g2_decap_8 FILLER_35_1057 ();
 sg13g2_decap_8 FILLER_35_1064 ();
 sg13g2_decap_8 FILLER_35_1071 ();
 sg13g2_decap_8 FILLER_35_1078 ();
 sg13g2_decap_8 FILLER_35_1085 ();
 sg13g2_decap_8 FILLER_35_1092 ();
 sg13g2_decap_8 FILLER_35_1099 ();
 sg13g2_decap_8 FILLER_35_1106 ();
 sg13g2_decap_8 FILLER_35_1113 ();
 sg13g2_decap_8 FILLER_35_1120 ();
 sg13g2_decap_8 FILLER_35_1127 ();
 sg13g2_decap_8 FILLER_35_1134 ();
 sg13g2_decap_8 FILLER_35_1141 ();
 sg13g2_decap_8 FILLER_35_1148 ();
 sg13g2_decap_8 FILLER_35_1155 ();
 sg13g2_decap_8 FILLER_35_1162 ();
 sg13g2_decap_8 FILLER_35_1169 ();
 sg13g2_decap_8 FILLER_35_1176 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_decap_8 FILLER_35_1190 ();
 sg13g2_decap_8 FILLER_35_1197 ();
 sg13g2_decap_8 FILLER_35_1204 ();
 sg13g2_decap_8 FILLER_35_1211 ();
 sg13g2_decap_8 FILLER_35_1218 ();
 sg13g2_decap_8 FILLER_35_1225 ();
 sg13g2_decap_8 FILLER_35_1232 ();
 sg13g2_decap_8 FILLER_35_1239 ();
 sg13g2_decap_8 FILLER_35_1246 ();
 sg13g2_decap_8 FILLER_35_1253 ();
 sg13g2_decap_8 FILLER_35_1260 ();
 sg13g2_decap_8 FILLER_35_1267 ();
 sg13g2_decap_8 FILLER_35_1274 ();
 sg13g2_decap_8 FILLER_35_1281 ();
 sg13g2_decap_8 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_decap_8 FILLER_35_1309 ();
 sg13g2_decap_8 FILLER_35_1316 ();
 sg13g2_decap_8 FILLER_35_1323 ();
 sg13g2_decap_8 FILLER_35_1330 ();
 sg13g2_decap_8 FILLER_35_1337 ();
 sg13g2_decap_8 FILLER_35_1344 ();
 sg13g2_decap_8 FILLER_35_1351 ();
 sg13g2_decap_8 FILLER_35_1358 ();
 sg13g2_decap_8 FILLER_35_1365 ();
 sg13g2_decap_8 FILLER_35_1372 ();
 sg13g2_decap_8 FILLER_35_1379 ();
 sg13g2_decap_8 FILLER_35_1386 ();
 sg13g2_decap_8 FILLER_35_1393 ();
 sg13g2_decap_8 FILLER_35_1400 ();
 sg13g2_decap_8 FILLER_35_1407 ();
 sg13g2_decap_8 FILLER_35_1414 ();
 sg13g2_decap_8 FILLER_35_1421 ();
 sg13g2_decap_8 FILLER_35_1428 ();
 sg13g2_decap_8 FILLER_35_1435 ();
 sg13g2_decap_8 FILLER_35_1442 ();
 sg13g2_decap_8 FILLER_35_1449 ();
 sg13g2_decap_8 FILLER_35_1456 ();
 sg13g2_decap_8 FILLER_35_1463 ();
 sg13g2_decap_8 FILLER_35_1470 ();
 sg13g2_decap_8 FILLER_35_1477 ();
 sg13g2_decap_8 FILLER_35_1484 ();
 sg13g2_decap_8 FILLER_35_1491 ();
 sg13g2_decap_8 FILLER_35_1498 ();
 sg13g2_decap_8 FILLER_35_1505 ();
 sg13g2_decap_8 FILLER_35_1512 ();
 sg13g2_decap_8 FILLER_35_1519 ();
 sg13g2_decap_8 FILLER_35_1526 ();
 sg13g2_decap_8 FILLER_35_1533 ();
 sg13g2_decap_8 FILLER_35_1540 ();
 sg13g2_decap_8 FILLER_35_1547 ();
 sg13g2_decap_8 FILLER_35_1554 ();
 sg13g2_decap_8 FILLER_35_1561 ();
 sg13g2_decap_8 FILLER_35_1568 ();
 sg13g2_decap_8 FILLER_35_1575 ();
 sg13g2_decap_8 FILLER_35_1582 ();
 sg13g2_decap_8 FILLER_35_1589 ();
 sg13g2_decap_8 FILLER_35_1596 ();
 sg13g2_decap_8 FILLER_35_1603 ();
 sg13g2_decap_8 FILLER_35_1610 ();
 sg13g2_decap_8 FILLER_35_1617 ();
 sg13g2_decap_8 FILLER_35_1624 ();
 sg13g2_decap_8 FILLER_35_1631 ();
 sg13g2_decap_8 FILLER_35_1638 ();
 sg13g2_decap_8 FILLER_35_1645 ();
 sg13g2_decap_8 FILLER_35_1652 ();
 sg13g2_decap_8 FILLER_35_1659 ();
 sg13g2_decap_8 FILLER_35_1666 ();
 sg13g2_decap_8 FILLER_35_1673 ();
 sg13g2_decap_8 FILLER_35_1680 ();
 sg13g2_decap_8 FILLER_35_1687 ();
 sg13g2_decap_8 FILLER_35_1694 ();
 sg13g2_decap_8 FILLER_35_1701 ();
 sg13g2_decap_8 FILLER_35_1708 ();
 sg13g2_decap_8 FILLER_35_1715 ();
 sg13g2_decap_8 FILLER_35_1722 ();
 sg13g2_decap_8 FILLER_35_1729 ();
 sg13g2_decap_8 FILLER_35_1736 ();
 sg13g2_decap_8 FILLER_35_1743 ();
 sg13g2_decap_8 FILLER_35_1750 ();
 sg13g2_decap_8 FILLER_35_1757 ();
 sg13g2_decap_4 FILLER_35_1764 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_36_868 ();
 sg13g2_decap_8 FILLER_36_875 ();
 sg13g2_decap_8 FILLER_36_882 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_decap_8 FILLER_36_896 ();
 sg13g2_decap_8 FILLER_36_903 ();
 sg13g2_decap_8 FILLER_36_910 ();
 sg13g2_decap_8 FILLER_36_917 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_decap_8 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_36_1029 ();
 sg13g2_decap_8 FILLER_36_1036 ();
 sg13g2_decap_8 FILLER_36_1043 ();
 sg13g2_decap_8 FILLER_36_1050 ();
 sg13g2_decap_8 FILLER_36_1057 ();
 sg13g2_decap_8 FILLER_36_1064 ();
 sg13g2_decap_8 FILLER_36_1071 ();
 sg13g2_decap_8 FILLER_36_1078 ();
 sg13g2_decap_8 FILLER_36_1085 ();
 sg13g2_decap_8 FILLER_36_1092 ();
 sg13g2_decap_8 FILLER_36_1099 ();
 sg13g2_decap_8 FILLER_36_1106 ();
 sg13g2_decap_8 FILLER_36_1113 ();
 sg13g2_decap_8 FILLER_36_1120 ();
 sg13g2_decap_8 FILLER_36_1127 ();
 sg13g2_decap_8 FILLER_36_1134 ();
 sg13g2_decap_8 FILLER_36_1141 ();
 sg13g2_decap_8 FILLER_36_1148 ();
 sg13g2_decap_8 FILLER_36_1155 ();
 sg13g2_decap_8 FILLER_36_1162 ();
 sg13g2_decap_8 FILLER_36_1169 ();
 sg13g2_decap_8 FILLER_36_1176 ();
 sg13g2_decap_8 FILLER_36_1183 ();
 sg13g2_decap_8 FILLER_36_1190 ();
 sg13g2_decap_8 FILLER_36_1197 ();
 sg13g2_decap_8 FILLER_36_1204 ();
 sg13g2_decap_8 FILLER_36_1211 ();
 sg13g2_decap_8 FILLER_36_1218 ();
 sg13g2_decap_8 FILLER_36_1225 ();
 sg13g2_decap_8 FILLER_36_1232 ();
 sg13g2_decap_8 FILLER_36_1239 ();
 sg13g2_decap_8 FILLER_36_1246 ();
 sg13g2_decap_8 FILLER_36_1253 ();
 sg13g2_decap_8 FILLER_36_1260 ();
 sg13g2_decap_8 FILLER_36_1267 ();
 sg13g2_decap_8 FILLER_36_1274 ();
 sg13g2_decap_8 FILLER_36_1281 ();
 sg13g2_decap_8 FILLER_36_1288 ();
 sg13g2_decap_8 FILLER_36_1295 ();
 sg13g2_decap_8 FILLER_36_1302 ();
 sg13g2_decap_8 FILLER_36_1309 ();
 sg13g2_decap_8 FILLER_36_1316 ();
 sg13g2_decap_8 FILLER_36_1323 ();
 sg13g2_decap_8 FILLER_36_1330 ();
 sg13g2_decap_8 FILLER_36_1337 ();
 sg13g2_decap_8 FILLER_36_1344 ();
 sg13g2_decap_8 FILLER_36_1351 ();
 sg13g2_decap_8 FILLER_36_1358 ();
 sg13g2_decap_8 FILLER_36_1365 ();
 sg13g2_decap_8 FILLER_36_1372 ();
 sg13g2_decap_8 FILLER_36_1379 ();
 sg13g2_decap_8 FILLER_36_1386 ();
 sg13g2_decap_8 FILLER_36_1393 ();
 sg13g2_decap_8 FILLER_36_1400 ();
 sg13g2_decap_8 FILLER_36_1407 ();
 sg13g2_decap_8 FILLER_36_1414 ();
 sg13g2_decap_8 FILLER_36_1421 ();
 sg13g2_decap_8 FILLER_36_1428 ();
 sg13g2_decap_8 FILLER_36_1435 ();
 sg13g2_decap_8 FILLER_36_1442 ();
 sg13g2_decap_8 FILLER_36_1449 ();
 sg13g2_decap_8 FILLER_36_1456 ();
 sg13g2_decap_8 FILLER_36_1463 ();
 sg13g2_decap_8 FILLER_36_1470 ();
 sg13g2_decap_8 FILLER_36_1477 ();
 sg13g2_decap_8 FILLER_36_1484 ();
 sg13g2_decap_8 FILLER_36_1491 ();
 sg13g2_decap_8 FILLER_36_1498 ();
 sg13g2_decap_8 FILLER_36_1505 ();
 sg13g2_decap_8 FILLER_36_1512 ();
 sg13g2_decap_8 FILLER_36_1519 ();
 sg13g2_decap_8 FILLER_36_1526 ();
 sg13g2_decap_8 FILLER_36_1533 ();
 sg13g2_decap_8 FILLER_36_1540 ();
 sg13g2_decap_8 FILLER_36_1547 ();
 sg13g2_decap_8 FILLER_36_1554 ();
 sg13g2_decap_8 FILLER_36_1561 ();
 sg13g2_decap_8 FILLER_36_1568 ();
 sg13g2_decap_8 FILLER_36_1575 ();
 sg13g2_decap_8 FILLER_36_1582 ();
 sg13g2_decap_8 FILLER_36_1589 ();
 sg13g2_decap_8 FILLER_36_1596 ();
 sg13g2_decap_8 FILLER_36_1603 ();
 sg13g2_decap_8 FILLER_36_1610 ();
 sg13g2_decap_8 FILLER_36_1617 ();
 sg13g2_decap_8 FILLER_36_1624 ();
 sg13g2_decap_8 FILLER_36_1631 ();
 sg13g2_decap_8 FILLER_36_1638 ();
 sg13g2_decap_8 FILLER_36_1645 ();
 sg13g2_decap_8 FILLER_36_1652 ();
 sg13g2_decap_8 FILLER_36_1659 ();
 sg13g2_decap_8 FILLER_36_1666 ();
 sg13g2_decap_8 FILLER_36_1673 ();
 sg13g2_decap_8 FILLER_36_1680 ();
 sg13g2_decap_8 FILLER_36_1687 ();
 sg13g2_decap_8 FILLER_36_1694 ();
 sg13g2_decap_8 FILLER_36_1701 ();
 sg13g2_decap_8 FILLER_36_1708 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_decap_8 FILLER_36_1722 ();
 sg13g2_decap_8 FILLER_36_1729 ();
 sg13g2_decap_8 FILLER_36_1736 ();
 sg13g2_decap_8 FILLER_36_1743 ();
 sg13g2_decap_8 FILLER_36_1750 ();
 sg13g2_decap_8 FILLER_36_1757 ();
 sg13g2_decap_4 FILLER_36_1764 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_37_1029 ();
 sg13g2_decap_8 FILLER_37_1036 ();
 sg13g2_decap_8 FILLER_37_1043 ();
 sg13g2_decap_8 FILLER_37_1050 ();
 sg13g2_decap_8 FILLER_37_1057 ();
 sg13g2_decap_8 FILLER_37_1064 ();
 sg13g2_decap_8 FILLER_37_1071 ();
 sg13g2_decap_8 FILLER_37_1078 ();
 sg13g2_decap_8 FILLER_37_1085 ();
 sg13g2_decap_8 FILLER_37_1092 ();
 sg13g2_decap_8 FILLER_37_1099 ();
 sg13g2_decap_8 FILLER_37_1106 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_decap_8 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_decap_8 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1155 ();
 sg13g2_decap_8 FILLER_37_1162 ();
 sg13g2_decap_8 FILLER_37_1169 ();
 sg13g2_decap_8 FILLER_37_1176 ();
 sg13g2_decap_8 FILLER_37_1183 ();
 sg13g2_decap_8 FILLER_37_1190 ();
 sg13g2_decap_8 FILLER_37_1197 ();
 sg13g2_decap_8 FILLER_37_1204 ();
 sg13g2_decap_8 FILLER_37_1211 ();
 sg13g2_decap_8 FILLER_37_1218 ();
 sg13g2_decap_8 FILLER_37_1225 ();
 sg13g2_decap_8 FILLER_37_1232 ();
 sg13g2_decap_8 FILLER_37_1239 ();
 sg13g2_decap_8 FILLER_37_1246 ();
 sg13g2_decap_8 FILLER_37_1253 ();
 sg13g2_decap_8 FILLER_37_1260 ();
 sg13g2_decap_8 FILLER_37_1267 ();
 sg13g2_decap_8 FILLER_37_1274 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_decap_8 FILLER_37_1288 ();
 sg13g2_decap_8 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1302 ();
 sg13g2_decap_8 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_decap_8 FILLER_37_1323 ();
 sg13g2_decap_8 FILLER_37_1330 ();
 sg13g2_decap_8 FILLER_37_1337 ();
 sg13g2_decap_8 FILLER_37_1344 ();
 sg13g2_decap_8 FILLER_37_1351 ();
 sg13g2_decap_8 FILLER_37_1358 ();
 sg13g2_decap_8 FILLER_37_1365 ();
 sg13g2_decap_8 FILLER_37_1372 ();
 sg13g2_decap_8 FILLER_37_1379 ();
 sg13g2_decap_8 FILLER_37_1386 ();
 sg13g2_decap_8 FILLER_37_1393 ();
 sg13g2_decap_8 FILLER_37_1400 ();
 sg13g2_decap_8 FILLER_37_1407 ();
 sg13g2_decap_8 FILLER_37_1414 ();
 sg13g2_decap_8 FILLER_37_1421 ();
 sg13g2_decap_8 FILLER_37_1428 ();
 sg13g2_decap_8 FILLER_37_1435 ();
 sg13g2_decap_8 FILLER_37_1442 ();
 sg13g2_decap_8 FILLER_37_1449 ();
 sg13g2_decap_8 FILLER_37_1456 ();
 sg13g2_decap_8 FILLER_37_1463 ();
 sg13g2_decap_8 FILLER_37_1470 ();
 sg13g2_decap_8 FILLER_37_1477 ();
 sg13g2_decap_8 FILLER_37_1484 ();
 sg13g2_decap_8 FILLER_37_1491 ();
 sg13g2_decap_8 FILLER_37_1498 ();
 sg13g2_decap_8 FILLER_37_1505 ();
 sg13g2_decap_8 FILLER_37_1512 ();
 sg13g2_decap_8 FILLER_37_1519 ();
 sg13g2_decap_8 FILLER_37_1526 ();
 sg13g2_decap_8 FILLER_37_1533 ();
 sg13g2_decap_8 FILLER_37_1540 ();
 sg13g2_decap_8 FILLER_37_1547 ();
 sg13g2_decap_8 FILLER_37_1554 ();
 sg13g2_decap_8 FILLER_37_1561 ();
 sg13g2_decap_8 FILLER_37_1568 ();
 sg13g2_decap_8 FILLER_37_1575 ();
 sg13g2_decap_8 FILLER_37_1582 ();
 sg13g2_decap_8 FILLER_37_1589 ();
 sg13g2_decap_8 FILLER_37_1596 ();
 sg13g2_decap_8 FILLER_37_1603 ();
 sg13g2_decap_8 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1617 ();
 sg13g2_decap_8 FILLER_37_1624 ();
 sg13g2_decap_8 FILLER_37_1631 ();
 sg13g2_decap_8 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1645 ();
 sg13g2_decap_8 FILLER_37_1652 ();
 sg13g2_decap_8 FILLER_37_1659 ();
 sg13g2_decap_8 FILLER_37_1666 ();
 sg13g2_decap_8 FILLER_37_1673 ();
 sg13g2_decap_8 FILLER_37_1680 ();
 sg13g2_decap_8 FILLER_37_1687 ();
 sg13g2_decap_8 FILLER_37_1694 ();
 sg13g2_decap_8 FILLER_37_1701 ();
 sg13g2_decap_8 FILLER_37_1708 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_decap_8 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1743 ();
 sg13g2_decap_8 FILLER_37_1750 ();
 sg13g2_decap_8 FILLER_37_1757 ();
 sg13g2_decap_4 FILLER_37_1764 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_38_1029 ();
 sg13g2_decap_8 FILLER_38_1036 ();
 sg13g2_decap_8 FILLER_38_1043 ();
 sg13g2_decap_8 FILLER_38_1050 ();
 sg13g2_decap_8 FILLER_38_1057 ();
 sg13g2_decap_8 FILLER_38_1064 ();
 sg13g2_decap_8 FILLER_38_1071 ();
 sg13g2_decap_8 FILLER_38_1078 ();
 sg13g2_decap_8 FILLER_38_1085 ();
 sg13g2_decap_8 FILLER_38_1092 ();
 sg13g2_decap_8 FILLER_38_1099 ();
 sg13g2_decap_8 FILLER_38_1106 ();
 sg13g2_decap_8 FILLER_38_1113 ();
 sg13g2_decap_8 FILLER_38_1120 ();
 sg13g2_decap_8 FILLER_38_1127 ();
 sg13g2_decap_8 FILLER_38_1134 ();
 sg13g2_decap_8 FILLER_38_1141 ();
 sg13g2_decap_8 FILLER_38_1148 ();
 sg13g2_decap_8 FILLER_38_1155 ();
 sg13g2_decap_8 FILLER_38_1162 ();
 sg13g2_decap_8 FILLER_38_1169 ();
 sg13g2_decap_8 FILLER_38_1176 ();
 sg13g2_decap_8 FILLER_38_1183 ();
 sg13g2_decap_8 FILLER_38_1190 ();
 sg13g2_decap_8 FILLER_38_1197 ();
 sg13g2_decap_8 FILLER_38_1204 ();
 sg13g2_decap_8 FILLER_38_1211 ();
 sg13g2_decap_8 FILLER_38_1218 ();
 sg13g2_decap_8 FILLER_38_1225 ();
 sg13g2_decap_8 FILLER_38_1232 ();
 sg13g2_decap_8 FILLER_38_1239 ();
 sg13g2_decap_8 FILLER_38_1246 ();
 sg13g2_decap_8 FILLER_38_1253 ();
 sg13g2_decap_8 FILLER_38_1260 ();
 sg13g2_decap_8 FILLER_38_1267 ();
 sg13g2_decap_8 FILLER_38_1274 ();
 sg13g2_decap_8 FILLER_38_1281 ();
 sg13g2_decap_8 FILLER_38_1288 ();
 sg13g2_decap_8 FILLER_38_1295 ();
 sg13g2_decap_8 FILLER_38_1302 ();
 sg13g2_decap_8 FILLER_38_1309 ();
 sg13g2_decap_8 FILLER_38_1316 ();
 sg13g2_decap_8 FILLER_38_1323 ();
 sg13g2_decap_8 FILLER_38_1330 ();
 sg13g2_decap_8 FILLER_38_1337 ();
 sg13g2_decap_8 FILLER_38_1344 ();
 sg13g2_decap_8 FILLER_38_1351 ();
 sg13g2_decap_8 FILLER_38_1358 ();
 sg13g2_decap_8 FILLER_38_1365 ();
 sg13g2_decap_8 FILLER_38_1372 ();
 sg13g2_decap_8 FILLER_38_1379 ();
 sg13g2_decap_8 FILLER_38_1386 ();
 sg13g2_decap_8 FILLER_38_1393 ();
 sg13g2_decap_8 FILLER_38_1400 ();
 sg13g2_decap_8 FILLER_38_1407 ();
 sg13g2_decap_8 FILLER_38_1414 ();
 sg13g2_decap_8 FILLER_38_1421 ();
 sg13g2_decap_8 FILLER_38_1428 ();
 sg13g2_decap_8 FILLER_38_1435 ();
 sg13g2_decap_8 FILLER_38_1442 ();
 sg13g2_decap_8 FILLER_38_1449 ();
 sg13g2_decap_8 FILLER_38_1456 ();
 sg13g2_decap_8 FILLER_38_1463 ();
 sg13g2_decap_8 FILLER_38_1470 ();
 sg13g2_decap_8 FILLER_38_1477 ();
 sg13g2_decap_8 FILLER_38_1484 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_decap_8 FILLER_38_1498 ();
 sg13g2_decap_8 FILLER_38_1505 ();
 sg13g2_decap_8 FILLER_38_1512 ();
 sg13g2_decap_8 FILLER_38_1519 ();
 sg13g2_decap_8 FILLER_38_1526 ();
 sg13g2_decap_8 FILLER_38_1533 ();
 sg13g2_decap_8 FILLER_38_1540 ();
 sg13g2_decap_8 FILLER_38_1547 ();
 sg13g2_decap_8 FILLER_38_1554 ();
 sg13g2_decap_8 FILLER_38_1561 ();
 sg13g2_decap_8 FILLER_38_1568 ();
 sg13g2_decap_8 FILLER_38_1575 ();
 sg13g2_decap_8 FILLER_38_1582 ();
 sg13g2_decap_8 FILLER_38_1589 ();
 sg13g2_decap_8 FILLER_38_1596 ();
 sg13g2_decap_8 FILLER_38_1603 ();
 sg13g2_decap_8 FILLER_38_1610 ();
 sg13g2_decap_8 FILLER_38_1617 ();
 sg13g2_decap_8 FILLER_38_1624 ();
 sg13g2_decap_8 FILLER_38_1631 ();
 sg13g2_decap_8 FILLER_38_1638 ();
 sg13g2_decap_8 FILLER_38_1645 ();
 sg13g2_decap_8 FILLER_38_1652 ();
 sg13g2_decap_8 FILLER_38_1659 ();
 sg13g2_decap_8 FILLER_38_1666 ();
 sg13g2_decap_8 FILLER_38_1673 ();
 sg13g2_decap_8 FILLER_38_1680 ();
 sg13g2_decap_8 FILLER_38_1687 ();
 sg13g2_decap_8 FILLER_38_1694 ();
 sg13g2_decap_8 FILLER_38_1701 ();
 sg13g2_decap_8 FILLER_38_1708 ();
 sg13g2_decap_8 FILLER_38_1715 ();
 sg13g2_decap_8 FILLER_38_1722 ();
 sg13g2_decap_8 FILLER_38_1729 ();
 sg13g2_decap_8 FILLER_38_1736 ();
 sg13g2_decap_8 FILLER_38_1743 ();
 sg13g2_decap_8 FILLER_38_1750 ();
 sg13g2_decap_8 FILLER_38_1757 ();
 sg13g2_decap_4 FILLER_38_1764 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_4 FILLER_39_826 ();
 sg13g2_fill_1 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_39_931 ();
 sg13g2_decap_8 FILLER_39_938 ();
 sg13g2_decap_8 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_966 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_decap_8 FILLER_39_980 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_8 FILLER_39_1029 ();
 sg13g2_decap_8 FILLER_39_1036 ();
 sg13g2_decap_8 FILLER_39_1043 ();
 sg13g2_decap_8 FILLER_39_1050 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_decap_8 FILLER_39_1064 ();
 sg13g2_decap_8 FILLER_39_1071 ();
 sg13g2_decap_8 FILLER_39_1078 ();
 sg13g2_decap_8 FILLER_39_1085 ();
 sg13g2_decap_8 FILLER_39_1092 ();
 sg13g2_decap_8 FILLER_39_1099 ();
 sg13g2_decap_8 FILLER_39_1106 ();
 sg13g2_decap_8 FILLER_39_1113 ();
 sg13g2_decap_8 FILLER_39_1120 ();
 sg13g2_decap_8 FILLER_39_1127 ();
 sg13g2_decap_8 FILLER_39_1134 ();
 sg13g2_decap_8 FILLER_39_1141 ();
 sg13g2_decap_8 FILLER_39_1148 ();
 sg13g2_decap_8 FILLER_39_1155 ();
 sg13g2_decap_8 FILLER_39_1162 ();
 sg13g2_decap_8 FILLER_39_1169 ();
 sg13g2_decap_8 FILLER_39_1176 ();
 sg13g2_decap_8 FILLER_39_1183 ();
 sg13g2_decap_8 FILLER_39_1190 ();
 sg13g2_decap_8 FILLER_39_1197 ();
 sg13g2_decap_8 FILLER_39_1204 ();
 sg13g2_decap_8 FILLER_39_1211 ();
 sg13g2_decap_8 FILLER_39_1218 ();
 sg13g2_decap_8 FILLER_39_1225 ();
 sg13g2_decap_8 FILLER_39_1232 ();
 sg13g2_decap_8 FILLER_39_1239 ();
 sg13g2_decap_8 FILLER_39_1246 ();
 sg13g2_decap_8 FILLER_39_1253 ();
 sg13g2_decap_8 FILLER_39_1260 ();
 sg13g2_decap_8 FILLER_39_1267 ();
 sg13g2_decap_8 FILLER_39_1274 ();
 sg13g2_decap_8 FILLER_39_1281 ();
 sg13g2_decap_8 FILLER_39_1288 ();
 sg13g2_decap_8 FILLER_39_1295 ();
 sg13g2_decap_8 FILLER_39_1302 ();
 sg13g2_decap_8 FILLER_39_1309 ();
 sg13g2_decap_8 FILLER_39_1316 ();
 sg13g2_decap_8 FILLER_39_1323 ();
 sg13g2_decap_8 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1337 ();
 sg13g2_decap_8 FILLER_39_1344 ();
 sg13g2_decap_8 FILLER_39_1351 ();
 sg13g2_decap_8 FILLER_39_1358 ();
 sg13g2_decap_8 FILLER_39_1365 ();
 sg13g2_decap_8 FILLER_39_1372 ();
 sg13g2_decap_8 FILLER_39_1379 ();
 sg13g2_decap_8 FILLER_39_1386 ();
 sg13g2_decap_8 FILLER_39_1393 ();
 sg13g2_decap_8 FILLER_39_1400 ();
 sg13g2_decap_8 FILLER_39_1407 ();
 sg13g2_decap_8 FILLER_39_1414 ();
 sg13g2_decap_8 FILLER_39_1421 ();
 sg13g2_decap_8 FILLER_39_1428 ();
 sg13g2_decap_8 FILLER_39_1435 ();
 sg13g2_decap_8 FILLER_39_1442 ();
 sg13g2_decap_8 FILLER_39_1449 ();
 sg13g2_decap_8 FILLER_39_1456 ();
 sg13g2_decap_8 FILLER_39_1463 ();
 sg13g2_decap_8 FILLER_39_1470 ();
 sg13g2_decap_8 FILLER_39_1477 ();
 sg13g2_decap_8 FILLER_39_1484 ();
 sg13g2_decap_8 FILLER_39_1491 ();
 sg13g2_decap_8 FILLER_39_1498 ();
 sg13g2_decap_8 FILLER_39_1505 ();
 sg13g2_decap_8 FILLER_39_1512 ();
 sg13g2_decap_8 FILLER_39_1519 ();
 sg13g2_decap_8 FILLER_39_1526 ();
 sg13g2_decap_8 FILLER_39_1533 ();
 sg13g2_decap_8 FILLER_39_1540 ();
 sg13g2_decap_8 FILLER_39_1547 ();
 sg13g2_decap_8 FILLER_39_1554 ();
 sg13g2_decap_8 FILLER_39_1561 ();
 sg13g2_decap_8 FILLER_39_1568 ();
 sg13g2_decap_8 FILLER_39_1575 ();
 sg13g2_decap_8 FILLER_39_1582 ();
 sg13g2_decap_8 FILLER_39_1589 ();
 sg13g2_decap_8 FILLER_39_1596 ();
 sg13g2_decap_8 FILLER_39_1603 ();
 sg13g2_decap_8 FILLER_39_1610 ();
 sg13g2_decap_8 FILLER_39_1617 ();
 sg13g2_decap_8 FILLER_39_1624 ();
 sg13g2_decap_8 FILLER_39_1631 ();
 sg13g2_decap_8 FILLER_39_1638 ();
 sg13g2_decap_8 FILLER_39_1645 ();
 sg13g2_decap_8 FILLER_39_1652 ();
 sg13g2_decap_8 FILLER_39_1659 ();
 sg13g2_decap_8 FILLER_39_1666 ();
 sg13g2_decap_8 FILLER_39_1673 ();
 sg13g2_decap_8 FILLER_39_1680 ();
 sg13g2_decap_8 FILLER_39_1687 ();
 sg13g2_decap_8 FILLER_39_1694 ();
 sg13g2_decap_8 FILLER_39_1701 ();
 sg13g2_decap_8 FILLER_39_1708 ();
 sg13g2_decap_8 FILLER_39_1715 ();
 sg13g2_decap_8 FILLER_39_1722 ();
 sg13g2_decap_8 FILLER_39_1729 ();
 sg13g2_decap_8 FILLER_39_1736 ();
 sg13g2_decap_8 FILLER_39_1743 ();
 sg13g2_decap_8 FILLER_39_1750 ();
 sg13g2_decap_8 FILLER_39_1757 ();
 sg13g2_decap_4 FILLER_39_1764 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_4 FILLER_40_812 ();
 sg13g2_fill_1 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_848 ();
 sg13g2_fill_2 FILLER_40_855 ();
 sg13g2_fill_1 FILLER_40_857 ();
 sg13g2_fill_2 FILLER_40_863 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_decap_8 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_40_884 ();
 sg13g2_decap_8 FILLER_40_891 ();
 sg13g2_fill_2 FILLER_40_898 ();
 sg13g2_fill_1 FILLER_40_900 ();
 sg13g2_fill_2 FILLER_40_904 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_8 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_8 FILLER_40_956 ();
 sg13g2_decap_8 FILLER_40_963 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_984 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_8 FILLER_40_998 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_decap_8 FILLER_40_1026 ();
 sg13g2_decap_8 FILLER_40_1033 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_decap_8 FILLER_40_1054 ();
 sg13g2_decap_8 FILLER_40_1061 ();
 sg13g2_decap_8 FILLER_40_1068 ();
 sg13g2_decap_8 FILLER_40_1075 ();
 sg13g2_decap_8 FILLER_40_1082 ();
 sg13g2_decap_8 FILLER_40_1089 ();
 sg13g2_decap_8 FILLER_40_1096 ();
 sg13g2_decap_8 FILLER_40_1103 ();
 sg13g2_decap_8 FILLER_40_1110 ();
 sg13g2_decap_8 FILLER_40_1117 ();
 sg13g2_decap_8 FILLER_40_1124 ();
 sg13g2_decap_8 FILLER_40_1131 ();
 sg13g2_decap_8 FILLER_40_1138 ();
 sg13g2_decap_8 FILLER_40_1145 ();
 sg13g2_decap_8 FILLER_40_1152 ();
 sg13g2_decap_8 FILLER_40_1159 ();
 sg13g2_decap_8 FILLER_40_1166 ();
 sg13g2_decap_8 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1180 ();
 sg13g2_decap_8 FILLER_40_1187 ();
 sg13g2_decap_8 FILLER_40_1194 ();
 sg13g2_decap_8 FILLER_40_1201 ();
 sg13g2_decap_8 FILLER_40_1208 ();
 sg13g2_decap_8 FILLER_40_1215 ();
 sg13g2_decap_8 FILLER_40_1222 ();
 sg13g2_decap_8 FILLER_40_1229 ();
 sg13g2_decap_8 FILLER_40_1236 ();
 sg13g2_decap_8 FILLER_40_1243 ();
 sg13g2_decap_8 FILLER_40_1250 ();
 sg13g2_decap_8 FILLER_40_1257 ();
 sg13g2_decap_8 FILLER_40_1264 ();
 sg13g2_decap_8 FILLER_40_1271 ();
 sg13g2_decap_8 FILLER_40_1278 ();
 sg13g2_decap_8 FILLER_40_1285 ();
 sg13g2_decap_8 FILLER_40_1292 ();
 sg13g2_decap_8 FILLER_40_1299 ();
 sg13g2_decap_8 FILLER_40_1306 ();
 sg13g2_decap_8 FILLER_40_1313 ();
 sg13g2_decap_8 FILLER_40_1320 ();
 sg13g2_decap_8 FILLER_40_1327 ();
 sg13g2_decap_8 FILLER_40_1334 ();
 sg13g2_decap_8 FILLER_40_1341 ();
 sg13g2_decap_8 FILLER_40_1348 ();
 sg13g2_decap_8 FILLER_40_1355 ();
 sg13g2_decap_8 FILLER_40_1362 ();
 sg13g2_decap_8 FILLER_40_1369 ();
 sg13g2_decap_8 FILLER_40_1376 ();
 sg13g2_decap_8 FILLER_40_1383 ();
 sg13g2_decap_8 FILLER_40_1390 ();
 sg13g2_decap_8 FILLER_40_1397 ();
 sg13g2_decap_8 FILLER_40_1404 ();
 sg13g2_decap_8 FILLER_40_1411 ();
 sg13g2_decap_8 FILLER_40_1418 ();
 sg13g2_decap_8 FILLER_40_1425 ();
 sg13g2_decap_8 FILLER_40_1432 ();
 sg13g2_decap_8 FILLER_40_1439 ();
 sg13g2_decap_8 FILLER_40_1446 ();
 sg13g2_decap_8 FILLER_40_1453 ();
 sg13g2_decap_8 FILLER_40_1460 ();
 sg13g2_decap_8 FILLER_40_1467 ();
 sg13g2_decap_8 FILLER_40_1474 ();
 sg13g2_decap_8 FILLER_40_1481 ();
 sg13g2_decap_8 FILLER_40_1488 ();
 sg13g2_decap_8 FILLER_40_1495 ();
 sg13g2_decap_8 FILLER_40_1502 ();
 sg13g2_decap_8 FILLER_40_1509 ();
 sg13g2_decap_8 FILLER_40_1516 ();
 sg13g2_decap_8 FILLER_40_1523 ();
 sg13g2_decap_8 FILLER_40_1530 ();
 sg13g2_decap_8 FILLER_40_1537 ();
 sg13g2_decap_8 FILLER_40_1544 ();
 sg13g2_decap_8 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1558 ();
 sg13g2_decap_8 FILLER_40_1565 ();
 sg13g2_decap_8 FILLER_40_1572 ();
 sg13g2_decap_8 FILLER_40_1579 ();
 sg13g2_decap_8 FILLER_40_1586 ();
 sg13g2_decap_8 FILLER_40_1593 ();
 sg13g2_decap_8 FILLER_40_1600 ();
 sg13g2_decap_8 FILLER_40_1607 ();
 sg13g2_decap_8 FILLER_40_1614 ();
 sg13g2_decap_8 FILLER_40_1621 ();
 sg13g2_decap_8 FILLER_40_1628 ();
 sg13g2_decap_8 FILLER_40_1635 ();
 sg13g2_decap_8 FILLER_40_1642 ();
 sg13g2_decap_8 FILLER_40_1649 ();
 sg13g2_decap_8 FILLER_40_1656 ();
 sg13g2_decap_8 FILLER_40_1663 ();
 sg13g2_decap_8 FILLER_40_1670 ();
 sg13g2_decap_8 FILLER_40_1677 ();
 sg13g2_decap_8 FILLER_40_1684 ();
 sg13g2_decap_8 FILLER_40_1691 ();
 sg13g2_decap_8 FILLER_40_1698 ();
 sg13g2_decap_8 FILLER_40_1705 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_4 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_792 ();
 sg13g2_decap_8 FILLER_41_799 ();
 sg13g2_fill_2 FILLER_41_818 ();
 sg13g2_fill_1 FILLER_41_851 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_fill_1 FILLER_41_862 ();
 sg13g2_decap_8 FILLER_41_876 ();
 sg13g2_decap_4 FILLER_41_883 ();
 sg13g2_fill_1 FILLER_41_887 ();
 sg13g2_fill_2 FILLER_41_895 ();
 sg13g2_fill_1 FILLER_41_897 ();
 sg13g2_fill_2 FILLER_41_903 ();
 sg13g2_fill_1 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_914 ();
 sg13g2_decap_8 FILLER_41_921 ();
 sg13g2_fill_1 FILLER_41_928 ();
 sg13g2_fill_2 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_fill_1 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_991 ();
 sg13g2_decap_8 FILLER_41_998 ();
 sg13g2_decap_8 FILLER_41_1005 ();
 sg13g2_decap_8 FILLER_41_1012 ();
 sg13g2_decap_8 FILLER_41_1019 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_8 FILLER_41_1033 ();
 sg13g2_decap_8 FILLER_41_1040 ();
 sg13g2_decap_8 FILLER_41_1047 ();
 sg13g2_decap_8 FILLER_41_1054 ();
 sg13g2_decap_8 FILLER_41_1061 ();
 sg13g2_decap_8 FILLER_41_1068 ();
 sg13g2_decap_8 FILLER_41_1075 ();
 sg13g2_decap_8 FILLER_41_1082 ();
 sg13g2_decap_8 FILLER_41_1089 ();
 sg13g2_decap_8 FILLER_41_1096 ();
 sg13g2_decap_8 FILLER_41_1103 ();
 sg13g2_decap_8 FILLER_41_1110 ();
 sg13g2_decap_8 FILLER_41_1117 ();
 sg13g2_decap_8 FILLER_41_1124 ();
 sg13g2_decap_8 FILLER_41_1131 ();
 sg13g2_decap_8 FILLER_41_1138 ();
 sg13g2_decap_8 FILLER_41_1145 ();
 sg13g2_decap_8 FILLER_41_1152 ();
 sg13g2_decap_8 FILLER_41_1159 ();
 sg13g2_decap_8 FILLER_41_1166 ();
 sg13g2_decap_8 FILLER_41_1173 ();
 sg13g2_decap_8 FILLER_41_1180 ();
 sg13g2_decap_8 FILLER_41_1187 ();
 sg13g2_decap_8 FILLER_41_1194 ();
 sg13g2_decap_8 FILLER_41_1201 ();
 sg13g2_decap_8 FILLER_41_1208 ();
 sg13g2_decap_8 FILLER_41_1215 ();
 sg13g2_decap_8 FILLER_41_1222 ();
 sg13g2_decap_8 FILLER_41_1229 ();
 sg13g2_decap_8 FILLER_41_1236 ();
 sg13g2_decap_8 FILLER_41_1243 ();
 sg13g2_decap_8 FILLER_41_1250 ();
 sg13g2_decap_8 FILLER_41_1257 ();
 sg13g2_decap_8 FILLER_41_1264 ();
 sg13g2_decap_8 FILLER_41_1271 ();
 sg13g2_decap_8 FILLER_41_1278 ();
 sg13g2_decap_8 FILLER_41_1285 ();
 sg13g2_decap_8 FILLER_41_1292 ();
 sg13g2_decap_8 FILLER_41_1299 ();
 sg13g2_decap_8 FILLER_41_1306 ();
 sg13g2_decap_8 FILLER_41_1313 ();
 sg13g2_decap_8 FILLER_41_1320 ();
 sg13g2_decap_8 FILLER_41_1327 ();
 sg13g2_decap_8 FILLER_41_1334 ();
 sg13g2_decap_8 FILLER_41_1341 ();
 sg13g2_decap_8 FILLER_41_1348 ();
 sg13g2_decap_8 FILLER_41_1355 ();
 sg13g2_decap_8 FILLER_41_1362 ();
 sg13g2_decap_8 FILLER_41_1369 ();
 sg13g2_fill_2 FILLER_41_1376 ();
 sg13g2_decap_8 FILLER_41_1383 ();
 sg13g2_decap_8 FILLER_41_1390 ();
 sg13g2_decap_8 FILLER_41_1397 ();
 sg13g2_decap_8 FILLER_41_1404 ();
 sg13g2_decap_8 FILLER_41_1411 ();
 sg13g2_decap_8 FILLER_41_1418 ();
 sg13g2_decap_8 FILLER_41_1425 ();
 sg13g2_fill_2 FILLER_41_1432 ();
 sg13g2_fill_1 FILLER_41_1434 ();
 sg13g2_decap_8 FILLER_41_1440 ();
 sg13g2_decap_8 FILLER_41_1447 ();
 sg13g2_decap_8 FILLER_41_1454 ();
 sg13g2_decap_8 FILLER_41_1461 ();
 sg13g2_decap_8 FILLER_41_1468 ();
 sg13g2_decap_8 FILLER_41_1475 ();
 sg13g2_decap_8 FILLER_41_1482 ();
 sg13g2_decap_8 FILLER_41_1489 ();
 sg13g2_decap_8 FILLER_41_1496 ();
 sg13g2_decap_8 FILLER_41_1503 ();
 sg13g2_decap_8 FILLER_41_1510 ();
 sg13g2_decap_8 FILLER_41_1517 ();
 sg13g2_decap_8 FILLER_41_1524 ();
 sg13g2_decap_8 FILLER_41_1531 ();
 sg13g2_decap_8 FILLER_41_1538 ();
 sg13g2_decap_8 FILLER_41_1545 ();
 sg13g2_decap_8 FILLER_41_1552 ();
 sg13g2_decap_8 FILLER_41_1559 ();
 sg13g2_decap_8 FILLER_41_1566 ();
 sg13g2_decap_8 FILLER_41_1573 ();
 sg13g2_decap_8 FILLER_41_1580 ();
 sg13g2_decap_8 FILLER_41_1587 ();
 sg13g2_decap_8 FILLER_41_1594 ();
 sg13g2_decap_8 FILLER_41_1601 ();
 sg13g2_decap_8 FILLER_41_1608 ();
 sg13g2_decap_8 FILLER_41_1615 ();
 sg13g2_decap_8 FILLER_41_1622 ();
 sg13g2_decap_8 FILLER_41_1629 ();
 sg13g2_decap_8 FILLER_41_1636 ();
 sg13g2_decap_8 FILLER_41_1643 ();
 sg13g2_decap_8 FILLER_41_1650 ();
 sg13g2_decap_8 FILLER_41_1657 ();
 sg13g2_decap_8 FILLER_41_1664 ();
 sg13g2_decap_8 FILLER_41_1671 ();
 sg13g2_decap_8 FILLER_41_1678 ();
 sg13g2_decap_8 FILLER_41_1685 ();
 sg13g2_decap_8 FILLER_41_1692 ();
 sg13g2_decap_8 FILLER_41_1699 ();
 sg13g2_decap_8 FILLER_41_1706 ();
 sg13g2_decap_8 FILLER_41_1713 ();
 sg13g2_decap_8 FILLER_41_1720 ();
 sg13g2_decap_8 FILLER_41_1727 ();
 sg13g2_decap_8 FILLER_41_1734 ();
 sg13g2_decap_8 FILLER_41_1741 ();
 sg13g2_decap_8 FILLER_41_1748 ();
 sg13g2_decap_8 FILLER_41_1755 ();
 sg13g2_decap_4 FILLER_41_1762 ();
 sg13g2_fill_2 FILLER_41_1766 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_fill_1 FILLER_42_345 ();
 sg13g2_decap_8 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_decap_8 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_42_415 ();
 sg13g2_decap_8 FILLER_42_422 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_443 ();
 sg13g2_decap_8 FILLER_42_450 ();
 sg13g2_decap_8 FILLER_42_457 ();
 sg13g2_decap_8 FILLER_42_464 ();
 sg13g2_decap_8 FILLER_42_471 ();
 sg13g2_decap_8 FILLER_42_478 ();
 sg13g2_decap_8 FILLER_42_485 ();
 sg13g2_decap_8 FILLER_42_492 ();
 sg13g2_decap_8 FILLER_42_499 ();
 sg13g2_decap_8 FILLER_42_506 ();
 sg13g2_decap_8 FILLER_42_513 ();
 sg13g2_decap_8 FILLER_42_520 ();
 sg13g2_decap_8 FILLER_42_527 ();
 sg13g2_decap_8 FILLER_42_534 ();
 sg13g2_decap_8 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_548 ();
 sg13g2_decap_8 FILLER_42_555 ();
 sg13g2_decap_8 FILLER_42_562 ();
 sg13g2_decap_8 FILLER_42_569 ();
 sg13g2_decap_8 FILLER_42_576 ();
 sg13g2_decap_8 FILLER_42_583 ();
 sg13g2_decap_8 FILLER_42_590 ();
 sg13g2_decap_8 FILLER_42_597 ();
 sg13g2_decap_8 FILLER_42_604 ();
 sg13g2_decap_8 FILLER_42_611 ();
 sg13g2_decap_8 FILLER_42_618 ();
 sg13g2_decap_8 FILLER_42_625 ();
 sg13g2_decap_8 FILLER_42_632 ();
 sg13g2_decap_8 FILLER_42_639 ();
 sg13g2_decap_8 FILLER_42_646 ();
 sg13g2_decap_8 FILLER_42_653 ();
 sg13g2_decap_8 FILLER_42_660 ();
 sg13g2_decap_8 FILLER_42_667 ();
 sg13g2_decap_8 FILLER_42_674 ();
 sg13g2_decap_8 FILLER_42_681 ();
 sg13g2_decap_8 FILLER_42_688 ();
 sg13g2_decap_8 FILLER_42_695 ();
 sg13g2_fill_1 FILLER_42_702 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_4 FILLER_42_717 ();
 sg13g2_fill_2 FILLER_42_721 ();
 sg13g2_fill_2 FILLER_42_728 ();
 sg13g2_fill_1 FILLER_42_730 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_746 ();
 sg13g2_decap_8 FILLER_42_753 ();
 sg13g2_decap_8 FILLER_42_760 ();
 sg13g2_decap_8 FILLER_42_767 ();
 sg13g2_fill_2 FILLER_42_774 ();
 sg13g2_fill_1 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_799 ();
 sg13g2_decap_8 FILLER_42_806 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_fill_1 FILLER_42_820 ();
 sg13g2_fill_1 FILLER_42_830 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_8 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_865 ();
 sg13g2_decap_4 FILLER_42_872 ();
 sg13g2_fill_1 FILLER_42_876 ();
 sg13g2_fill_1 FILLER_42_893 ();
 sg13g2_fill_1 FILLER_42_902 ();
 sg13g2_decap_8 FILLER_42_917 ();
 sg13g2_decap_4 FILLER_42_924 ();
 sg13g2_fill_2 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_934 ();
 sg13g2_decap_4 FILLER_42_941 ();
 sg13g2_fill_2 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_951 ();
 sg13g2_decap_4 FILLER_42_958 ();
 sg13g2_fill_2 FILLER_42_970 ();
 sg13g2_fill_1 FILLER_42_972 ();
 sg13g2_decap_8 FILLER_42_981 ();
 sg13g2_decap_8 FILLER_42_988 ();
 sg13g2_decap_8 FILLER_42_995 ();
 sg13g2_decap_8 FILLER_42_1002 ();
 sg13g2_decap_8 FILLER_42_1009 ();
 sg13g2_decap_8 FILLER_42_1016 ();
 sg13g2_decap_8 FILLER_42_1023 ();
 sg13g2_decap_8 FILLER_42_1030 ();
 sg13g2_decap_8 FILLER_42_1037 ();
 sg13g2_decap_8 FILLER_42_1044 ();
 sg13g2_decap_8 FILLER_42_1051 ();
 sg13g2_decap_8 FILLER_42_1058 ();
 sg13g2_decap_8 FILLER_42_1065 ();
 sg13g2_decap_8 FILLER_42_1072 ();
 sg13g2_fill_1 FILLER_42_1079 ();
 sg13g2_decap_8 FILLER_42_1083 ();
 sg13g2_decap_8 FILLER_42_1090 ();
 sg13g2_decap_8 FILLER_42_1097 ();
 sg13g2_decap_8 FILLER_42_1104 ();
 sg13g2_decap_8 FILLER_42_1111 ();
 sg13g2_decap_8 FILLER_42_1118 ();
 sg13g2_decap_8 FILLER_42_1125 ();
 sg13g2_decap_8 FILLER_42_1132 ();
 sg13g2_decap_8 FILLER_42_1139 ();
 sg13g2_decap_8 FILLER_42_1146 ();
 sg13g2_decap_8 FILLER_42_1153 ();
 sg13g2_decap_8 FILLER_42_1160 ();
 sg13g2_decap_8 FILLER_42_1167 ();
 sg13g2_decap_8 FILLER_42_1174 ();
 sg13g2_decap_8 FILLER_42_1181 ();
 sg13g2_decap_8 FILLER_42_1188 ();
 sg13g2_decap_8 FILLER_42_1195 ();
 sg13g2_decap_8 FILLER_42_1202 ();
 sg13g2_decap_8 FILLER_42_1209 ();
 sg13g2_decap_8 FILLER_42_1216 ();
 sg13g2_decap_8 FILLER_42_1223 ();
 sg13g2_decap_8 FILLER_42_1230 ();
 sg13g2_decap_8 FILLER_42_1237 ();
 sg13g2_decap_8 FILLER_42_1244 ();
 sg13g2_decap_8 FILLER_42_1251 ();
 sg13g2_decap_8 FILLER_42_1258 ();
 sg13g2_decap_8 FILLER_42_1265 ();
 sg13g2_decap_8 FILLER_42_1272 ();
 sg13g2_decap_8 FILLER_42_1279 ();
 sg13g2_decap_8 FILLER_42_1286 ();
 sg13g2_decap_8 FILLER_42_1293 ();
 sg13g2_decap_8 FILLER_42_1300 ();
 sg13g2_decap_8 FILLER_42_1307 ();
 sg13g2_decap_8 FILLER_42_1314 ();
 sg13g2_decap_8 FILLER_42_1321 ();
 sg13g2_decap_8 FILLER_42_1328 ();
 sg13g2_decap_8 FILLER_42_1335 ();
 sg13g2_decap_8 FILLER_42_1342 ();
 sg13g2_decap_8 FILLER_42_1349 ();
 sg13g2_decap_4 FILLER_42_1356 ();
 sg13g2_decap_4 FILLER_42_1363 ();
 sg13g2_fill_1 FILLER_42_1367 ();
 sg13g2_fill_1 FILLER_42_1375 ();
 sg13g2_decap_8 FILLER_42_1392 ();
 sg13g2_decap_8 FILLER_42_1399 ();
 sg13g2_decap_8 FILLER_42_1406 ();
 sg13g2_decap_8 FILLER_42_1413 ();
 sg13g2_decap_4 FILLER_42_1420 ();
 sg13g2_fill_1 FILLER_42_1424 ();
 sg13g2_decap_8 FILLER_42_1453 ();
 sg13g2_decap_8 FILLER_42_1460 ();
 sg13g2_decap_8 FILLER_42_1467 ();
 sg13g2_decap_8 FILLER_42_1474 ();
 sg13g2_decap_8 FILLER_42_1481 ();
 sg13g2_decap_8 FILLER_42_1488 ();
 sg13g2_decap_8 FILLER_42_1495 ();
 sg13g2_decap_8 FILLER_42_1502 ();
 sg13g2_decap_8 FILLER_42_1509 ();
 sg13g2_decap_8 FILLER_42_1516 ();
 sg13g2_decap_8 FILLER_42_1523 ();
 sg13g2_decap_8 FILLER_42_1530 ();
 sg13g2_decap_8 FILLER_42_1537 ();
 sg13g2_decap_8 FILLER_42_1544 ();
 sg13g2_decap_8 FILLER_42_1551 ();
 sg13g2_decap_8 FILLER_42_1558 ();
 sg13g2_decap_8 FILLER_42_1565 ();
 sg13g2_decap_8 FILLER_42_1572 ();
 sg13g2_decap_8 FILLER_42_1579 ();
 sg13g2_decap_8 FILLER_42_1586 ();
 sg13g2_decap_8 FILLER_42_1593 ();
 sg13g2_decap_8 FILLER_42_1600 ();
 sg13g2_decap_8 FILLER_42_1607 ();
 sg13g2_decap_8 FILLER_42_1614 ();
 sg13g2_decap_8 FILLER_42_1621 ();
 sg13g2_decap_8 FILLER_42_1628 ();
 sg13g2_decap_8 FILLER_42_1635 ();
 sg13g2_decap_8 FILLER_42_1642 ();
 sg13g2_decap_8 FILLER_42_1649 ();
 sg13g2_decap_8 FILLER_42_1656 ();
 sg13g2_decap_8 FILLER_42_1663 ();
 sg13g2_decap_8 FILLER_42_1670 ();
 sg13g2_decap_8 FILLER_42_1677 ();
 sg13g2_decap_8 FILLER_42_1684 ();
 sg13g2_decap_8 FILLER_42_1691 ();
 sg13g2_decap_8 FILLER_42_1698 ();
 sg13g2_decap_8 FILLER_42_1705 ();
 sg13g2_decap_8 FILLER_42_1712 ();
 sg13g2_decap_8 FILLER_42_1719 ();
 sg13g2_decap_8 FILLER_42_1726 ();
 sg13g2_decap_8 FILLER_42_1733 ();
 sg13g2_decap_8 FILLER_42_1740 ();
 sg13g2_decap_8 FILLER_42_1747 ();
 sg13g2_decap_8 FILLER_42_1754 ();
 sg13g2_decap_8 FILLER_42_1761 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_decap_8 FILLER_43_286 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_decap_8 FILLER_43_300 ();
 sg13g2_decap_8 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_314 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_327 ();
 sg13g2_decap_4 FILLER_43_334 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_421 ();
 sg13g2_decap_8 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_43_435 ();
 sg13g2_decap_8 FILLER_43_442 ();
 sg13g2_decap_8 FILLER_43_449 ();
 sg13g2_decap_8 FILLER_43_456 ();
 sg13g2_decap_8 FILLER_43_463 ();
 sg13g2_decap_8 FILLER_43_470 ();
 sg13g2_decap_8 FILLER_43_477 ();
 sg13g2_decap_8 FILLER_43_484 ();
 sg13g2_decap_8 FILLER_43_491 ();
 sg13g2_decap_8 FILLER_43_498 ();
 sg13g2_decap_8 FILLER_43_505 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_decap_8 FILLER_43_519 ();
 sg13g2_decap_8 FILLER_43_526 ();
 sg13g2_decap_8 FILLER_43_533 ();
 sg13g2_decap_8 FILLER_43_540 ();
 sg13g2_decap_8 FILLER_43_547 ();
 sg13g2_decap_8 FILLER_43_554 ();
 sg13g2_decap_8 FILLER_43_561 ();
 sg13g2_decap_8 FILLER_43_568 ();
 sg13g2_decap_8 FILLER_43_575 ();
 sg13g2_decap_8 FILLER_43_582 ();
 sg13g2_decap_8 FILLER_43_589 ();
 sg13g2_decap_8 FILLER_43_596 ();
 sg13g2_decap_8 FILLER_43_603 ();
 sg13g2_decap_8 FILLER_43_610 ();
 sg13g2_decap_8 FILLER_43_617 ();
 sg13g2_decap_8 FILLER_43_624 ();
 sg13g2_decap_8 FILLER_43_631 ();
 sg13g2_decap_8 FILLER_43_638 ();
 sg13g2_decap_8 FILLER_43_645 ();
 sg13g2_decap_8 FILLER_43_652 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_decap_8 FILLER_43_666 ();
 sg13g2_decap_8 FILLER_43_673 ();
 sg13g2_decap_8 FILLER_43_680 ();
 sg13g2_fill_2 FILLER_43_687 ();
 sg13g2_fill_1 FILLER_43_689 ();
 sg13g2_decap_8 FILLER_43_698 ();
 sg13g2_decap_4 FILLER_43_705 ();
 sg13g2_fill_2 FILLER_43_709 ();
 sg13g2_fill_1 FILLER_43_742 ();
 sg13g2_fill_2 FILLER_43_756 ();
 sg13g2_fill_2 FILLER_43_773 ();
 sg13g2_decap_8 FILLER_43_801 ();
 sg13g2_decap_8 FILLER_43_808 ();
 sg13g2_decap_8 FILLER_43_815 ();
 sg13g2_decap_8 FILLER_43_822 ();
 sg13g2_decap_8 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_fill_2 FILLER_43_894 ();
 sg13g2_fill_1 FILLER_43_896 ();
 sg13g2_fill_2 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_916 ();
 sg13g2_decap_4 FILLER_43_923 ();
 sg13g2_fill_1 FILLER_43_927 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_fill_1 FILLER_43_976 ();
 sg13g2_decap_8 FILLER_43_986 ();
 sg13g2_decap_8 FILLER_43_993 ();
 sg13g2_decap_8 FILLER_43_1000 ();
 sg13g2_decap_8 FILLER_43_1031 ();
 sg13g2_decap_8 FILLER_43_1038 ();
 sg13g2_decap_8 FILLER_43_1045 ();
 sg13g2_decap_8 FILLER_43_1052 ();
 sg13g2_decap_8 FILLER_43_1059 ();
 sg13g2_fill_2 FILLER_43_1066 ();
 sg13g2_fill_1 FILLER_43_1068 ();
 sg13g2_decap_8 FILLER_43_1077 ();
 sg13g2_decap_4 FILLER_43_1084 ();
 sg13g2_fill_2 FILLER_43_1088 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_decap_8 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1178 ();
 sg13g2_decap_8 FILLER_43_1185 ();
 sg13g2_decap_8 FILLER_43_1192 ();
 sg13g2_decap_8 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_decap_8 FILLER_43_1213 ();
 sg13g2_decap_8 FILLER_43_1220 ();
 sg13g2_decap_8 FILLER_43_1227 ();
 sg13g2_decap_8 FILLER_43_1234 ();
 sg13g2_decap_8 FILLER_43_1241 ();
 sg13g2_decap_8 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1255 ();
 sg13g2_decap_8 FILLER_43_1262 ();
 sg13g2_decap_8 FILLER_43_1269 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_4 FILLER_43_1304 ();
 sg13g2_fill_2 FILLER_43_1308 ();
 sg13g2_fill_1 FILLER_43_1319 ();
 sg13g2_decap_8 FILLER_43_1329 ();
 sg13g2_decap_8 FILLER_43_1336 ();
 sg13g2_fill_1 FILLER_43_1343 ();
 sg13g2_decap_8 FILLER_43_1394 ();
 sg13g2_decap_4 FILLER_43_1401 ();
 sg13g2_fill_1 FILLER_43_1405 ();
 sg13g2_decap_8 FILLER_43_1422 ();
 sg13g2_fill_2 FILLER_43_1429 ();
 sg13g2_fill_1 FILLER_43_1463 ();
 sg13g2_decap_4 FILLER_43_1471 ();
 sg13g2_decap_8 FILLER_43_1485 ();
 sg13g2_fill_1 FILLER_43_1492 ();
 sg13g2_decap_8 FILLER_43_1497 ();
 sg13g2_decap_8 FILLER_43_1504 ();
 sg13g2_decap_8 FILLER_43_1511 ();
 sg13g2_decap_8 FILLER_43_1518 ();
 sg13g2_decap_8 FILLER_43_1525 ();
 sg13g2_decap_8 FILLER_43_1532 ();
 sg13g2_decap_8 FILLER_43_1539 ();
 sg13g2_decap_8 FILLER_43_1546 ();
 sg13g2_decap_8 FILLER_43_1553 ();
 sg13g2_decap_8 FILLER_43_1560 ();
 sg13g2_decap_8 FILLER_43_1567 ();
 sg13g2_decap_8 FILLER_43_1574 ();
 sg13g2_decap_8 FILLER_43_1581 ();
 sg13g2_decap_8 FILLER_43_1588 ();
 sg13g2_decap_8 FILLER_43_1595 ();
 sg13g2_decap_8 FILLER_43_1602 ();
 sg13g2_decap_8 FILLER_43_1609 ();
 sg13g2_decap_8 FILLER_43_1616 ();
 sg13g2_decap_8 FILLER_43_1623 ();
 sg13g2_decap_8 FILLER_43_1630 ();
 sg13g2_decap_8 FILLER_43_1637 ();
 sg13g2_decap_8 FILLER_43_1644 ();
 sg13g2_decap_8 FILLER_43_1651 ();
 sg13g2_decap_8 FILLER_43_1658 ();
 sg13g2_decap_8 FILLER_43_1665 ();
 sg13g2_decap_8 FILLER_43_1672 ();
 sg13g2_decap_8 FILLER_43_1679 ();
 sg13g2_decap_8 FILLER_43_1686 ();
 sg13g2_decap_8 FILLER_43_1693 ();
 sg13g2_decap_8 FILLER_43_1700 ();
 sg13g2_decap_8 FILLER_43_1707 ();
 sg13g2_decap_8 FILLER_43_1714 ();
 sg13g2_decap_8 FILLER_43_1721 ();
 sg13g2_decap_8 FILLER_43_1728 ();
 sg13g2_decap_8 FILLER_43_1735 ();
 sg13g2_decap_8 FILLER_43_1742 ();
 sg13g2_decap_8 FILLER_43_1749 ();
 sg13g2_decap_8 FILLER_43_1756 ();
 sg13g2_decap_4 FILLER_43_1763 ();
 sg13g2_fill_1 FILLER_43_1767 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_fill_2 FILLER_44_276 ();
 sg13g2_decap_4 FILLER_44_285 ();
 sg13g2_fill_1 FILLER_44_289 ();
 sg13g2_fill_1 FILLER_44_308 ();
 sg13g2_fill_2 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_fill_2 FILLER_44_362 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_fill_2 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_432 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_450 ();
 sg13g2_decap_8 FILLER_44_457 ();
 sg13g2_decap_8 FILLER_44_464 ();
 sg13g2_decap_8 FILLER_44_471 ();
 sg13g2_decap_8 FILLER_44_478 ();
 sg13g2_decap_8 FILLER_44_485 ();
 sg13g2_decap_8 FILLER_44_492 ();
 sg13g2_decap_8 FILLER_44_499 ();
 sg13g2_decap_8 FILLER_44_506 ();
 sg13g2_decap_8 FILLER_44_513 ();
 sg13g2_decap_8 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_527 ();
 sg13g2_decap_8 FILLER_44_534 ();
 sg13g2_decap_8 FILLER_44_541 ();
 sg13g2_decap_8 FILLER_44_548 ();
 sg13g2_decap_8 FILLER_44_555 ();
 sg13g2_decap_8 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_569 ();
 sg13g2_decap_8 FILLER_44_576 ();
 sg13g2_decap_8 FILLER_44_583 ();
 sg13g2_decap_8 FILLER_44_590 ();
 sg13g2_decap_8 FILLER_44_597 ();
 sg13g2_decap_8 FILLER_44_604 ();
 sg13g2_decap_8 FILLER_44_611 ();
 sg13g2_decap_8 FILLER_44_618 ();
 sg13g2_decap_8 FILLER_44_625 ();
 sg13g2_decap_8 FILLER_44_632 ();
 sg13g2_decap_8 FILLER_44_639 ();
 sg13g2_decap_8 FILLER_44_646 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_decap_8 FILLER_44_660 ();
 sg13g2_decap_8 FILLER_44_667 ();
 sg13g2_decap_8 FILLER_44_674 ();
 sg13g2_decap_8 FILLER_44_681 ();
 sg13g2_decap_8 FILLER_44_688 ();
 sg13g2_fill_2 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_697 ();
 sg13g2_fill_2 FILLER_44_724 ();
 sg13g2_fill_2 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_4 FILLER_44_872 ();
 sg13g2_fill_2 FILLER_44_876 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_fill_1 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_44_944 ();
 sg13g2_decap_4 FILLER_44_951 ();
 sg13g2_fill_2 FILLER_44_955 ();
 sg13g2_decap_8 FILLER_44_965 ();
 sg13g2_decap_8 FILLER_44_972 ();
 sg13g2_decap_8 FILLER_44_979 ();
 sg13g2_fill_1 FILLER_44_1000 ();
 sg13g2_decap_8 FILLER_44_1029 ();
 sg13g2_fill_1 FILLER_44_1036 ();
 sg13g2_fill_1 FILLER_44_1049 ();
 sg13g2_fill_2 FILLER_44_1054 ();
 sg13g2_decap_4 FILLER_44_1061 ();
 sg13g2_fill_1 FILLER_44_1090 ();
 sg13g2_decap_8 FILLER_44_1096 ();
 sg13g2_decap_8 FILLER_44_1103 ();
 sg13g2_fill_2 FILLER_44_1110 ();
 sg13g2_fill_1 FILLER_44_1112 ();
 sg13g2_decap_8 FILLER_44_1117 ();
 sg13g2_fill_2 FILLER_44_1124 ();
 sg13g2_decap_8 FILLER_44_1129 ();
 sg13g2_decap_8 FILLER_44_1136 ();
 sg13g2_decap_8 FILLER_44_1143 ();
 sg13g2_decap_8 FILLER_44_1150 ();
 sg13g2_decap_8 FILLER_44_1157 ();
 sg13g2_decap_8 FILLER_44_1164 ();
 sg13g2_decap_8 FILLER_44_1171 ();
 sg13g2_decap_8 FILLER_44_1178 ();
 sg13g2_decap_8 FILLER_44_1185 ();
 sg13g2_decap_8 FILLER_44_1192 ();
 sg13g2_decap_8 FILLER_44_1199 ();
 sg13g2_decap_8 FILLER_44_1206 ();
 sg13g2_decap_8 FILLER_44_1213 ();
 sg13g2_decap_8 FILLER_44_1220 ();
 sg13g2_decap_8 FILLER_44_1227 ();
 sg13g2_decap_8 FILLER_44_1234 ();
 sg13g2_decap_8 FILLER_44_1241 ();
 sg13g2_decap_8 FILLER_44_1248 ();
 sg13g2_decap_8 FILLER_44_1255 ();
 sg13g2_decap_8 FILLER_44_1262 ();
 sg13g2_decap_8 FILLER_44_1269 ();
 sg13g2_decap_8 FILLER_44_1276 ();
 sg13g2_decap_8 FILLER_44_1283 ();
 sg13g2_decap_8 FILLER_44_1290 ();
 sg13g2_fill_2 FILLER_44_1297 ();
 sg13g2_fill_2 FILLER_44_1315 ();
 sg13g2_fill_1 FILLER_44_1317 ();
 sg13g2_decap_8 FILLER_44_1330 ();
 sg13g2_decap_8 FILLER_44_1337 ();
 sg13g2_fill_1 FILLER_44_1344 ();
 sg13g2_decap_8 FILLER_44_1352 ();
 sg13g2_fill_2 FILLER_44_1363 ();
 sg13g2_decap_8 FILLER_44_1380 ();
 sg13g2_decap_8 FILLER_44_1387 ();
 sg13g2_decap_8 FILLER_44_1394 ();
 sg13g2_decap_4 FILLER_44_1401 ();
 sg13g2_fill_1 FILLER_44_1411 ();
 sg13g2_decap_8 FILLER_44_1421 ();
 sg13g2_decap_8 FILLER_44_1428 ();
 sg13g2_decap_8 FILLER_44_1435 ();
 sg13g2_decap_8 FILLER_44_1452 ();
 sg13g2_decap_4 FILLER_44_1459 ();
 sg13g2_fill_2 FILLER_44_1463 ();
 sg13g2_fill_2 FILLER_44_1470 ();
 sg13g2_fill_1 FILLER_44_1472 ();
 sg13g2_decap_8 FILLER_44_1496 ();
 sg13g2_decap_4 FILLER_44_1503 ();
 sg13g2_fill_2 FILLER_44_1507 ();
 sg13g2_decap_8 FILLER_44_1513 ();
 sg13g2_fill_1 FILLER_44_1520 ();
 sg13g2_decap_8 FILLER_44_1534 ();
 sg13g2_decap_8 FILLER_44_1541 ();
 sg13g2_decap_8 FILLER_44_1548 ();
 sg13g2_decap_8 FILLER_44_1555 ();
 sg13g2_decap_8 FILLER_44_1562 ();
 sg13g2_decap_8 FILLER_44_1569 ();
 sg13g2_decap_8 FILLER_44_1576 ();
 sg13g2_decap_8 FILLER_44_1583 ();
 sg13g2_decap_8 FILLER_44_1590 ();
 sg13g2_decap_8 FILLER_44_1597 ();
 sg13g2_decap_8 FILLER_44_1604 ();
 sg13g2_decap_8 FILLER_44_1611 ();
 sg13g2_decap_8 FILLER_44_1618 ();
 sg13g2_decap_8 FILLER_44_1625 ();
 sg13g2_decap_8 FILLER_44_1632 ();
 sg13g2_decap_8 FILLER_44_1639 ();
 sg13g2_decap_8 FILLER_44_1646 ();
 sg13g2_decap_8 FILLER_44_1653 ();
 sg13g2_decap_8 FILLER_44_1660 ();
 sg13g2_decap_8 FILLER_44_1667 ();
 sg13g2_decap_8 FILLER_44_1674 ();
 sg13g2_decap_8 FILLER_44_1681 ();
 sg13g2_decap_8 FILLER_44_1688 ();
 sg13g2_decap_8 FILLER_44_1695 ();
 sg13g2_decap_8 FILLER_44_1702 ();
 sg13g2_decap_8 FILLER_44_1709 ();
 sg13g2_decap_8 FILLER_44_1716 ();
 sg13g2_decap_8 FILLER_44_1723 ();
 sg13g2_decap_8 FILLER_44_1730 ();
 sg13g2_decap_8 FILLER_44_1737 ();
 sg13g2_decap_8 FILLER_44_1744 ();
 sg13g2_decap_8 FILLER_44_1751 ();
 sg13g2_decap_8 FILLER_44_1758 ();
 sg13g2_fill_2 FILLER_44_1765 ();
 sg13g2_fill_1 FILLER_44_1767 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_fill_2 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_decap_8 FILLER_45_291 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_decap_8 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_decap_8 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_4 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_4 FILLER_45_389 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_fill_1 FILLER_45_430 ();
 sg13g2_fill_2 FILLER_45_443 ();
 sg13g2_decap_8 FILLER_45_460 ();
 sg13g2_decap_8 FILLER_45_467 ();
 sg13g2_decap_4 FILLER_45_474 ();
 sg13g2_fill_2 FILLER_45_478 ();
 sg13g2_decap_4 FILLER_45_496 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_507 ();
 sg13g2_decap_8 FILLER_45_514 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_decap_8 FILLER_45_528 ();
 sg13g2_decap_8 FILLER_45_535 ();
 sg13g2_decap_8 FILLER_45_542 ();
 sg13g2_decap_8 FILLER_45_549 ();
 sg13g2_decap_8 FILLER_45_556 ();
 sg13g2_decap_8 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_8 FILLER_45_598 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_8 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_decap_8 FILLER_45_654 ();
 sg13g2_decap_8 FILLER_45_661 ();
 sg13g2_decap_4 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_fill_2 FILLER_45_690 ();
 sg13g2_decap_8 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_decap_8 FILLER_45_711 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_764 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_4 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_4 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_decap_8 FILLER_45_859 ();
 sg13g2_decap_4 FILLER_45_866 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_decap_8 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_decap_4 FILLER_45_952 ();
 sg13g2_fill_1 FILLER_45_956 ();
 sg13g2_decap_8 FILLER_45_971 ();
 sg13g2_decap_8 FILLER_45_978 ();
 sg13g2_decap_8 FILLER_45_985 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_decap_8 FILLER_45_1027 ();
 sg13g2_decap_8 FILLER_45_1034 ();
 sg13g2_decap_4 FILLER_45_1041 ();
 sg13g2_fill_1 FILLER_45_1045 ();
 sg13g2_decap_4 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1086 ();
 sg13g2_decap_8 FILLER_45_1093 ();
 sg13g2_fill_2 FILLER_45_1100 ();
 sg13g2_decap_8 FILLER_45_1110 ();
 sg13g2_fill_1 FILLER_45_1117 ();
 sg13g2_fill_1 FILLER_45_1131 ();
 sg13g2_decap_8 FILLER_45_1153 ();
 sg13g2_decap_8 FILLER_45_1160 ();
 sg13g2_decap_8 FILLER_45_1167 ();
 sg13g2_decap_8 FILLER_45_1174 ();
 sg13g2_decap_8 FILLER_45_1181 ();
 sg13g2_decap_8 FILLER_45_1188 ();
 sg13g2_decap_8 FILLER_45_1195 ();
 sg13g2_decap_8 FILLER_45_1202 ();
 sg13g2_decap_8 FILLER_45_1209 ();
 sg13g2_decap_8 FILLER_45_1216 ();
 sg13g2_decap_8 FILLER_45_1223 ();
 sg13g2_decap_8 FILLER_45_1230 ();
 sg13g2_decap_8 FILLER_45_1237 ();
 sg13g2_decap_8 FILLER_45_1244 ();
 sg13g2_decap_8 FILLER_45_1251 ();
 sg13g2_decap_8 FILLER_45_1258 ();
 sg13g2_decap_8 FILLER_45_1265 ();
 sg13g2_decap_8 FILLER_45_1272 ();
 sg13g2_decap_8 FILLER_45_1279 ();
 sg13g2_decap_4 FILLER_45_1286 ();
 sg13g2_fill_2 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1305 ();
 sg13g2_decap_4 FILLER_45_1312 ();
 sg13g2_decap_8 FILLER_45_1333 ();
 sg13g2_decap_8 FILLER_45_1340 ();
 sg13g2_decap_8 FILLER_45_1347 ();
 sg13g2_decap_8 FILLER_45_1354 ();
 sg13g2_decap_4 FILLER_45_1361 ();
 sg13g2_fill_2 FILLER_45_1365 ();
 sg13g2_decap_8 FILLER_45_1371 ();
 sg13g2_decap_8 FILLER_45_1378 ();
 sg13g2_decap_8 FILLER_45_1385 ();
 sg13g2_decap_8 FILLER_45_1392 ();
 sg13g2_decap_8 FILLER_45_1399 ();
 sg13g2_decap_8 FILLER_45_1422 ();
 sg13g2_decap_8 FILLER_45_1429 ();
 sg13g2_decap_8 FILLER_45_1436 ();
 sg13g2_decap_8 FILLER_45_1443 ();
 sg13g2_decap_8 FILLER_45_1450 ();
 sg13g2_decap_8 FILLER_45_1457 ();
 sg13g2_decap_8 FILLER_45_1464 ();
 sg13g2_decap_4 FILLER_45_1471 ();
 sg13g2_fill_1 FILLER_45_1475 ();
 sg13g2_decap_8 FILLER_45_1480 ();
 sg13g2_decap_8 FILLER_45_1487 ();
 sg13g2_decap_8 FILLER_45_1497 ();
 sg13g2_decap_4 FILLER_45_1504 ();
 sg13g2_decap_8 FILLER_45_1512 ();
 sg13g2_fill_1 FILLER_45_1519 ();
 sg13g2_fill_2 FILLER_45_1527 ();
 sg13g2_decap_8 FILLER_45_1541 ();
 sg13g2_decap_8 FILLER_45_1548 ();
 sg13g2_decap_8 FILLER_45_1555 ();
 sg13g2_decap_8 FILLER_45_1562 ();
 sg13g2_decap_8 FILLER_45_1569 ();
 sg13g2_decap_8 FILLER_45_1576 ();
 sg13g2_decap_8 FILLER_45_1583 ();
 sg13g2_decap_8 FILLER_45_1590 ();
 sg13g2_decap_8 FILLER_45_1597 ();
 sg13g2_decap_8 FILLER_45_1604 ();
 sg13g2_decap_8 FILLER_45_1611 ();
 sg13g2_decap_8 FILLER_45_1618 ();
 sg13g2_decap_8 FILLER_45_1625 ();
 sg13g2_decap_8 FILLER_45_1632 ();
 sg13g2_decap_8 FILLER_45_1639 ();
 sg13g2_decap_8 FILLER_45_1646 ();
 sg13g2_decap_8 FILLER_45_1653 ();
 sg13g2_decap_8 FILLER_45_1660 ();
 sg13g2_decap_8 FILLER_45_1667 ();
 sg13g2_decap_8 FILLER_45_1674 ();
 sg13g2_decap_8 FILLER_45_1681 ();
 sg13g2_decap_8 FILLER_45_1688 ();
 sg13g2_decap_8 FILLER_45_1695 ();
 sg13g2_decap_8 FILLER_45_1702 ();
 sg13g2_decap_8 FILLER_45_1709 ();
 sg13g2_decap_8 FILLER_45_1716 ();
 sg13g2_decap_8 FILLER_45_1723 ();
 sg13g2_decap_8 FILLER_45_1730 ();
 sg13g2_decap_8 FILLER_45_1737 ();
 sg13g2_decap_8 FILLER_45_1744 ();
 sg13g2_decap_8 FILLER_45_1751 ();
 sg13g2_decap_8 FILLER_45_1758 ();
 sg13g2_fill_2 FILLER_45_1765 ();
 sg13g2_fill_1 FILLER_45_1767 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_4 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_decap_4 FILLER_46_260 ();
 sg13g2_decap_8 FILLER_46_277 ();
 sg13g2_decap_8 FILLER_46_284 ();
 sg13g2_decap_8 FILLER_46_291 ();
 sg13g2_decap_8 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_305 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_decap_8 FILLER_46_323 ();
 sg13g2_decap_8 FILLER_46_330 ();
 sg13g2_decap_8 FILLER_46_337 ();
 sg13g2_decap_8 FILLER_46_344 ();
 sg13g2_decap_8 FILLER_46_351 ();
 sg13g2_decap_8 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_46_421 ();
 sg13g2_decap_8 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_46_435 ();
 sg13g2_decap_8 FILLER_46_442 ();
 sg13g2_fill_2 FILLER_46_449 ();
 sg13g2_fill_1 FILLER_46_451 ();
 sg13g2_decap_8 FILLER_46_457 ();
 sg13g2_decap_8 FILLER_46_464 ();
 sg13g2_decap_8 FILLER_46_471 ();
 sg13g2_decap_8 FILLER_46_478 ();
 sg13g2_decap_4 FILLER_46_491 ();
 sg13g2_fill_2 FILLER_46_495 ();
 sg13g2_decap_4 FILLER_46_520 ();
 sg13g2_fill_2 FILLER_46_524 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_fill_2 FILLER_46_651 ();
 sg13g2_fill_1 FILLER_46_653 ();
 sg13g2_decap_8 FILLER_46_657 ();
 sg13g2_fill_2 FILLER_46_664 ();
 sg13g2_fill_2 FILLER_46_679 ();
 sg13g2_fill_2 FILLER_46_702 ();
 sg13g2_decap_8 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_723 ();
 sg13g2_decap_8 FILLER_46_730 ();
 sg13g2_decap_8 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_744 ();
 sg13g2_decap_8 FILLER_46_751 ();
 sg13g2_decap_4 FILLER_46_758 ();
 sg13g2_fill_2 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_fill_2 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_817 ();
 sg13g2_fill_1 FILLER_46_824 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_fill_2 FILLER_46_856 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_4 FILLER_46_889 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_913 ();
 sg13g2_decap_8 FILLER_46_920 ();
 sg13g2_decap_8 FILLER_46_927 ();
 sg13g2_decap_8 FILLER_46_934 ();
 sg13g2_decap_8 FILLER_46_941 ();
 sg13g2_decap_8 FILLER_46_948 ();
 sg13g2_decap_8 FILLER_46_955 ();
 sg13g2_decap_8 FILLER_46_962 ();
 sg13g2_decap_8 FILLER_46_969 ();
 sg13g2_decap_8 FILLER_46_976 ();
 sg13g2_decap_4 FILLER_46_983 ();
 sg13g2_fill_2 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_1014 ();
 sg13g2_decap_8 FILLER_46_1021 ();
 sg13g2_decap_8 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_46_1035 ();
 sg13g2_decap_8 FILLER_46_1042 ();
 sg13g2_decap_8 FILLER_46_1049 ();
 sg13g2_decap_8 FILLER_46_1056 ();
 sg13g2_decap_8 FILLER_46_1063 ();
 sg13g2_decap_8 FILLER_46_1070 ();
 sg13g2_decap_8 FILLER_46_1077 ();
 sg13g2_decap_4 FILLER_46_1084 ();
 sg13g2_decap_8 FILLER_46_1097 ();
 sg13g2_decap_8 FILLER_46_1104 ();
 sg13g2_fill_1 FILLER_46_1111 ();
 sg13g2_fill_2 FILLER_46_1117 ();
 sg13g2_fill_1 FILLER_46_1119 ();
 sg13g2_decap_8 FILLER_46_1124 ();
 sg13g2_decap_8 FILLER_46_1131 ();
 sg13g2_fill_2 FILLER_46_1138 ();
 sg13g2_decap_8 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1155 ();
 sg13g2_decap_8 FILLER_46_1162 ();
 sg13g2_decap_8 FILLER_46_1169 ();
 sg13g2_decap_8 FILLER_46_1176 ();
 sg13g2_decap_8 FILLER_46_1183 ();
 sg13g2_decap_8 FILLER_46_1190 ();
 sg13g2_decap_8 FILLER_46_1197 ();
 sg13g2_decap_8 FILLER_46_1204 ();
 sg13g2_decap_8 FILLER_46_1211 ();
 sg13g2_decap_8 FILLER_46_1218 ();
 sg13g2_decap_8 FILLER_46_1225 ();
 sg13g2_decap_8 FILLER_46_1232 ();
 sg13g2_decap_8 FILLER_46_1239 ();
 sg13g2_decap_8 FILLER_46_1246 ();
 sg13g2_decap_8 FILLER_46_1253 ();
 sg13g2_decap_8 FILLER_46_1260 ();
 sg13g2_decap_8 FILLER_46_1267 ();
 sg13g2_decap_8 FILLER_46_1274 ();
 sg13g2_decap_8 FILLER_46_1281 ();
 sg13g2_decap_8 FILLER_46_1288 ();
 sg13g2_decap_8 FILLER_46_1295 ();
 sg13g2_decap_4 FILLER_46_1302 ();
 sg13g2_fill_1 FILLER_46_1306 ();
 sg13g2_decap_4 FILLER_46_1315 ();
 sg13g2_decap_8 FILLER_46_1322 ();
 sg13g2_decap_8 FILLER_46_1329 ();
 sg13g2_decap_8 FILLER_46_1336 ();
 sg13g2_decap_8 FILLER_46_1343 ();
 sg13g2_decap_8 FILLER_46_1350 ();
 sg13g2_decap_8 FILLER_46_1357 ();
 sg13g2_decap_4 FILLER_46_1364 ();
 sg13g2_fill_1 FILLER_46_1368 ();
 sg13g2_decap_8 FILLER_46_1378 ();
 sg13g2_decap_8 FILLER_46_1385 ();
 sg13g2_decap_8 FILLER_46_1392 ();
 sg13g2_decap_8 FILLER_46_1399 ();
 sg13g2_decap_4 FILLER_46_1406 ();
 sg13g2_fill_2 FILLER_46_1410 ();
 sg13g2_decap_8 FILLER_46_1426 ();
 sg13g2_decap_8 FILLER_46_1433 ();
 sg13g2_decap_8 FILLER_46_1440 ();
 sg13g2_decap_8 FILLER_46_1447 ();
 sg13g2_decap_8 FILLER_46_1454 ();
 sg13g2_fill_2 FILLER_46_1461 ();
 sg13g2_fill_1 FILLER_46_1463 ();
 sg13g2_decap_8 FILLER_46_1480 ();
 sg13g2_decap_8 FILLER_46_1487 ();
 sg13g2_decap_8 FILLER_46_1494 ();
 sg13g2_decap_8 FILLER_46_1501 ();
 sg13g2_decap_8 FILLER_46_1508 ();
 sg13g2_fill_1 FILLER_46_1531 ();
 sg13g2_decap_8 FILLER_46_1537 ();
 sg13g2_decap_8 FILLER_46_1544 ();
 sg13g2_decap_8 FILLER_46_1551 ();
 sg13g2_decap_8 FILLER_46_1558 ();
 sg13g2_decap_8 FILLER_46_1565 ();
 sg13g2_decap_8 FILLER_46_1572 ();
 sg13g2_decap_8 FILLER_46_1579 ();
 sg13g2_decap_8 FILLER_46_1586 ();
 sg13g2_decap_8 FILLER_46_1593 ();
 sg13g2_decap_8 FILLER_46_1600 ();
 sg13g2_decap_8 FILLER_46_1607 ();
 sg13g2_decap_8 FILLER_46_1614 ();
 sg13g2_decap_8 FILLER_46_1621 ();
 sg13g2_decap_8 FILLER_46_1628 ();
 sg13g2_decap_8 FILLER_46_1635 ();
 sg13g2_decap_8 FILLER_46_1642 ();
 sg13g2_decap_8 FILLER_46_1649 ();
 sg13g2_decap_8 FILLER_46_1656 ();
 sg13g2_decap_8 FILLER_46_1663 ();
 sg13g2_decap_8 FILLER_46_1670 ();
 sg13g2_decap_8 FILLER_46_1677 ();
 sg13g2_decap_8 FILLER_46_1684 ();
 sg13g2_decap_8 FILLER_46_1691 ();
 sg13g2_decap_8 FILLER_46_1698 ();
 sg13g2_decap_8 FILLER_46_1705 ();
 sg13g2_decap_8 FILLER_46_1712 ();
 sg13g2_decap_8 FILLER_46_1719 ();
 sg13g2_decap_8 FILLER_46_1726 ();
 sg13g2_decap_8 FILLER_46_1733 ();
 sg13g2_decap_8 FILLER_46_1740 ();
 sg13g2_decap_8 FILLER_46_1747 ();
 sg13g2_decap_8 FILLER_46_1754 ();
 sg13g2_decap_8 FILLER_46_1761 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_fill_2 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_246 ();
 sg13g2_decap_8 FILLER_47_253 ();
 sg13g2_decap_8 FILLER_47_260 ();
 sg13g2_decap_4 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_decap_8 FILLER_47_290 ();
 sg13g2_decap_8 FILLER_47_297 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_decap_8 FILLER_47_337 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_fill_2 FILLER_47_400 ();
 sg13g2_fill_1 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_47_421 ();
 sg13g2_decap_8 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_47_435 ();
 sg13g2_decap_8 FILLER_47_442 ();
 sg13g2_decap_8 FILLER_47_449 ();
 sg13g2_decap_8 FILLER_47_456 ();
 sg13g2_fill_1 FILLER_47_471 ();
 sg13g2_decap_8 FILLER_47_492 ();
 sg13g2_decap_8 FILLER_47_499 ();
 sg13g2_fill_2 FILLER_47_506 ();
 sg13g2_decap_8 FILLER_47_517 ();
 sg13g2_decap_8 FILLER_47_544 ();
 sg13g2_decap_8 FILLER_47_551 ();
 sg13g2_decap_8 FILLER_47_558 ();
 sg13g2_fill_2 FILLER_47_565 ();
 sg13g2_fill_1 FILLER_47_571 ();
 sg13g2_fill_2 FILLER_47_580 ();
 sg13g2_decap_8 FILLER_47_586 ();
 sg13g2_decap_8 FILLER_47_593 ();
 sg13g2_decap_8 FILLER_47_600 ();
 sg13g2_decap_8 FILLER_47_607 ();
 sg13g2_decap_8 FILLER_47_614 ();
 sg13g2_decap_8 FILLER_47_621 ();
 sg13g2_decap_8 FILLER_47_628 ();
 sg13g2_decap_8 FILLER_47_635 ();
 sg13g2_decap_8 FILLER_47_642 ();
 sg13g2_fill_1 FILLER_47_649 ();
 sg13g2_decap_8 FILLER_47_678 ();
 sg13g2_fill_1 FILLER_47_685 ();
 sg13g2_decap_8 FILLER_47_699 ();
 sg13g2_decap_8 FILLER_47_706 ();
 sg13g2_decap_8 FILLER_47_713 ();
 sg13g2_decap_8 FILLER_47_720 ();
 sg13g2_decap_8 FILLER_47_727 ();
 sg13g2_decap_8 FILLER_47_734 ();
 sg13g2_decap_8 FILLER_47_741 ();
 sg13g2_decap_8 FILLER_47_748 ();
 sg13g2_fill_1 FILLER_47_755 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_decap_8 FILLER_47_786 ();
 sg13g2_decap_4 FILLER_47_793 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_fill_2 FILLER_47_849 ();
 sg13g2_fill_1 FILLER_47_851 ();
 sg13g2_decap_8 FILLER_47_876 ();
 sg13g2_decap_8 FILLER_47_883 ();
 sg13g2_decap_8 FILLER_47_890 ();
 sg13g2_fill_2 FILLER_47_897 ();
 sg13g2_fill_1 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_fill_2 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_953 ();
 sg13g2_decap_8 FILLER_47_960 ();
 sg13g2_decap_8 FILLER_47_967 ();
 sg13g2_decap_8 FILLER_47_974 ();
 sg13g2_decap_8 FILLER_47_981 ();
 sg13g2_decap_8 FILLER_47_988 ();
 sg13g2_decap_8 FILLER_47_995 ();
 sg13g2_decap_8 FILLER_47_1002 ();
 sg13g2_decap_8 FILLER_47_1009 ();
 sg13g2_decap_8 FILLER_47_1016 ();
 sg13g2_decap_4 FILLER_47_1023 ();
 sg13g2_fill_2 FILLER_47_1035 ();
 sg13g2_fill_2 FILLER_47_1040 ();
 sg13g2_decap_8 FILLER_47_1051 ();
 sg13g2_decap_8 FILLER_47_1058 ();
 sg13g2_decap_8 FILLER_47_1065 ();
 sg13g2_decap_8 FILLER_47_1072 ();
 sg13g2_decap_8 FILLER_47_1079 ();
 sg13g2_decap_8 FILLER_47_1086 ();
 sg13g2_decap_8 FILLER_47_1093 ();
 sg13g2_decap_8 FILLER_47_1100 ();
 sg13g2_decap_8 FILLER_47_1107 ();
 sg13g2_decap_8 FILLER_47_1114 ();
 sg13g2_decap_8 FILLER_47_1121 ();
 sg13g2_decap_8 FILLER_47_1128 ();
 sg13g2_fill_1 FILLER_47_1135 ();
 sg13g2_decap_8 FILLER_47_1149 ();
 sg13g2_decap_8 FILLER_47_1156 ();
 sg13g2_decap_8 FILLER_47_1163 ();
 sg13g2_decap_8 FILLER_47_1170 ();
 sg13g2_decap_8 FILLER_47_1177 ();
 sg13g2_decap_8 FILLER_47_1184 ();
 sg13g2_decap_8 FILLER_47_1191 ();
 sg13g2_decap_8 FILLER_47_1198 ();
 sg13g2_decap_8 FILLER_47_1205 ();
 sg13g2_decap_8 FILLER_47_1212 ();
 sg13g2_decap_8 FILLER_47_1219 ();
 sg13g2_decap_8 FILLER_47_1226 ();
 sg13g2_decap_8 FILLER_47_1233 ();
 sg13g2_decap_8 FILLER_47_1240 ();
 sg13g2_decap_8 FILLER_47_1247 ();
 sg13g2_decap_8 FILLER_47_1254 ();
 sg13g2_decap_8 FILLER_47_1261 ();
 sg13g2_decap_8 FILLER_47_1268 ();
 sg13g2_decap_8 FILLER_47_1275 ();
 sg13g2_decap_8 FILLER_47_1282 ();
 sg13g2_decap_8 FILLER_47_1289 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_decap_8 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1310 ();
 sg13g2_decap_8 FILLER_47_1317 ();
 sg13g2_decap_8 FILLER_47_1324 ();
 sg13g2_decap_8 FILLER_47_1331 ();
 sg13g2_decap_8 FILLER_47_1338 ();
 sg13g2_decap_8 FILLER_47_1345 ();
 sg13g2_decap_8 FILLER_47_1352 ();
 sg13g2_decap_8 FILLER_47_1359 ();
 sg13g2_decap_8 FILLER_47_1366 ();
 sg13g2_decap_8 FILLER_47_1373 ();
 sg13g2_decap_8 FILLER_47_1380 ();
 sg13g2_decap_8 FILLER_47_1387 ();
 sg13g2_decap_8 FILLER_47_1394 ();
 sg13g2_decap_8 FILLER_47_1401 ();
 sg13g2_decap_8 FILLER_47_1416 ();
 sg13g2_decap_8 FILLER_47_1423 ();
 sg13g2_decap_8 FILLER_47_1430 ();
 sg13g2_decap_8 FILLER_47_1437 ();
 sg13g2_decap_8 FILLER_47_1455 ();
 sg13g2_fill_1 FILLER_47_1462 ();
 sg13g2_decap_8 FILLER_47_1483 ();
 sg13g2_decap_8 FILLER_47_1490 ();
 sg13g2_decap_8 FILLER_47_1497 ();
 sg13g2_decap_8 FILLER_47_1504 ();
 sg13g2_decap_8 FILLER_47_1511 ();
 sg13g2_decap_4 FILLER_47_1518 ();
 sg13g2_fill_1 FILLER_47_1522 ();
 sg13g2_decap_8 FILLER_47_1546 ();
 sg13g2_decap_8 FILLER_47_1553 ();
 sg13g2_fill_1 FILLER_47_1560 ();
 sg13g2_decap_8 FILLER_47_1582 ();
 sg13g2_decap_8 FILLER_47_1589 ();
 sg13g2_decap_8 FILLER_47_1596 ();
 sg13g2_decap_8 FILLER_47_1603 ();
 sg13g2_decap_8 FILLER_47_1610 ();
 sg13g2_decap_8 FILLER_47_1617 ();
 sg13g2_decap_8 FILLER_47_1624 ();
 sg13g2_decap_8 FILLER_47_1631 ();
 sg13g2_decap_8 FILLER_47_1638 ();
 sg13g2_decap_8 FILLER_47_1645 ();
 sg13g2_decap_8 FILLER_47_1652 ();
 sg13g2_decap_8 FILLER_47_1659 ();
 sg13g2_decap_8 FILLER_47_1666 ();
 sg13g2_decap_8 FILLER_47_1673 ();
 sg13g2_decap_8 FILLER_47_1680 ();
 sg13g2_decap_8 FILLER_47_1687 ();
 sg13g2_decap_8 FILLER_47_1694 ();
 sg13g2_decap_8 FILLER_47_1701 ();
 sg13g2_decap_8 FILLER_47_1708 ();
 sg13g2_decap_8 FILLER_47_1715 ();
 sg13g2_decap_8 FILLER_47_1722 ();
 sg13g2_decap_8 FILLER_47_1729 ();
 sg13g2_decap_8 FILLER_47_1736 ();
 sg13g2_decap_8 FILLER_47_1743 ();
 sg13g2_decap_8 FILLER_47_1750 ();
 sg13g2_decap_8 FILLER_47_1757 ();
 sg13g2_decap_4 FILLER_47_1764 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_4 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_decap_4 FILLER_48_358 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_fill_2 FILLER_48_409 ();
 sg13g2_decap_8 FILLER_48_416 ();
 sg13g2_decap_8 FILLER_48_423 ();
 sg13g2_decap_8 FILLER_48_430 ();
 sg13g2_decap_8 FILLER_48_437 ();
 sg13g2_decap_8 FILLER_48_444 ();
 sg13g2_decap_8 FILLER_48_451 ();
 sg13g2_decap_8 FILLER_48_458 ();
 sg13g2_decap_8 FILLER_48_465 ();
 sg13g2_decap_8 FILLER_48_472 ();
 sg13g2_decap_8 FILLER_48_479 ();
 sg13g2_decap_8 FILLER_48_486 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_fill_1 FILLER_48_495 ();
 sg13g2_fill_1 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_514 ();
 sg13g2_decap_8 FILLER_48_521 ();
 sg13g2_decap_8 FILLER_48_528 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_8 FILLER_48_542 ();
 sg13g2_decap_4 FILLER_48_549 ();
 sg13g2_fill_2 FILLER_48_553 ();
 sg13g2_fill_2 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_586 ();
 sg13g2_decap_8 FILLER_48_593 ();
 sg13g2_decap_8 FILLER_48_600 ();
 sg13g2_decap_8 FILLER_48_607 ();
 sg13g2_decap_8 FILLER_48_614 ();
 sg13g2_decap_8 FILLER_48_621 ();
 sg13g2_decap_8 FILLER_48_628 ();
 sg13g2_fill_1 FILLER_48_635 ();
 sg13g2_fill_1 FILLER_48_656 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_4 FILLER_48_728 ();
 sg13g2_fill_1 FILLER_48_732 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_decap_8 FILLER_48_759 ();
 sg13g2_decap_8 FILLER_48_766 ();
 sg13g2_decap_8 FILLER_48_773 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_decap_8 FILLER_48_787 ();
 sg13g2_decap_8 FILLER_48_794 ();
 sg13g2_decap_8 FILLER_48_801 ();
 sg13g2_decap_8 FILLER_48_808 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_fill_2 FILLER_48_850 ();
 sg13g2_fill_1 FILLER_48_852 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_4 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_919 ();
 sg13g2_decap_8 FILLER_48_926 ();
 sg13g2_decap_8 FILLER_48_933 ();
 sg13g2_decap_8 FILLER_48_940 ();
 sg13g2_decap_4 FILLER_48_955 ();
 sg13g2_decap_4 FILLER_48_980 ();
 sg13g2_fill_2 FILLER_48_984 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_48_1029 ();
 sg13g2_decap_8 FILLER_48_1036 ();
 sg13g2_decap_8 FILLER_48_1043 ();
 sg13g2_decap_8 FILLER_48_1050 ();
 sg13g2_decap_8 FILLER_48_1057 ();
 sg13g2_decap_4 FILLER_48_1064 ();
 sg13g2_fill_2 FILLER_48_1068 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_4 FILLER_48_1092 ();
 sg13g2_fill_2 FILLER_48_1096 ();
 sg13g2_decap_8 FILLER_48_1111 ();
 sg13g2_decap_4 FILLER_48_1118 ();
 sg13g2_fill_1 FILLER_48_1122 ();
 sg13g2_fill_1 FILLER_48_1128 ();
 sg13g2_fill_2 FILLER_48_1137 ();
 sg13g2_decap_8 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1154 ();
 sg13g2_decap_8 FILLER_48_1161 ();
 sg13g2_fill_1 FILLER_48_1168 ();
 sg13g2_decap_8 FILLER_48_1221 ();
 sg13g2_decap_8 FILLER_48_1228 ();
 sg13g2_decap_8 FILLER_48_1235 ();
 sg13g2_decap_8 FILLER_48_1242 ();
 sg13g2_decap_8 FILLER_48_1249 ();
 sg13g2_decap_8 FILLER_48_1256 ();
 sg13g2_decap_8 FILLER_48_1263 ();
 sg13g2_decap_8 FILLER_48_1270 ();
 sg13g2_decap_8 FILLER_48_1277 ();
 sg13g2_decap_8 FILLER_48_1284 ();
 sg13g2_decap_8 FILLER_48_1291 ();
 sg13g2_decap_8 FILLER_48_1298 ();
 sg13g2_decap_8 FILLER_48_1305 ();
 sg13g2_decap_8 FILLER_48_1312 ();
 sg13g2_decap_8 FILLER_48_1319 ();
 sg13g2_decap_8 FILLER_48_1326 ();
 sg13g2_decap_8 FILLER_48_1346 ();
 sg13g2_decap_8 FILLER_48_1353 ();
 sg13g2_decap_4 FILLER_48_1360 ();
 sg13g2_fill_1 FILLER_48_1364 ();
 sg13g2_decap_8 FILLER_48_1383 ();
 sg13g2_decap_8 FILLER_48_1390 ();
 sg13g2_decap_8 FILLER_48_1397 ();
 sg13g2_fill_1 FILLER_48_1404 ();
 sg13g2_decap_8 FILLER_48_1415 ();
 sg13g2_decap_8 FILLER_48_1422 ();
 sg13g2_decap_8 FILLER_48_1429 ();
 sg13g2_decap_8 FILLER_48_1436 ();
 sg13g2_fill_2 FILLER_48_1443 ();
 sg13g2_decap_8 FILLER_48_1464 ();
 sg13g2_fill_2 FILLER_48_1471 ();
 sg13g2_decap_8 FILLER_48_1481 ();
 sg13g2_decap_8 FILLER_48_1488 ();
 sg13g2_decap_8 FILLER_48_1495 ();
 sg13g2_decap_8 FILLER_48_1502 ();
 sg13g2_decap_8 FILLER_48_1509 ();
 sg13g2_fill_2 FILLER_48_1516 ();
 sg13g2_fill_1 FILLER_48_1518 ();
 sg13g2_fill_2 FILLER_48_1537 ();
 sg13g2_fill_2 FILLER_48_1551 ();
 sg13g2_fill_2 FILLER_48_1558 ();
 sg13g2_decap_8 FILLER_48_1584 ();
 sg13g2_decap_8 FILLER_48_1591 ();
 sg13g2_decap_8 FILLER_48_1598 ();
 sg13g2_decap_8 FILLER_48_1605 ();
 sg13g2_decap_8 FILLER_48_1612 ();
 sg13g2_decap_8 FILLER_48_1619 ();
 sg13g2_decap_8 FILLER_48_1626 ();
 sg13g2_decap_8 FILLER_48_1633 ();
 sg13g2_decap_8 FILLER_48_1640 ();
 sg13g2_decap_8 FILLER_48_1647 ();
 sg13g2_decap_8 FILLER_48_1654 ();
 sg13g2_decap_8 FILLER_48_1661 ();
 sg13g2_decap_8 FILLER_48_1668 ();
 sg13g2_decap_8 FILLER_48_1675 ();
 sg13g2_decap_8 FILLER_48_1682 ();
 sg13g2_decap_8 FILLER_48_1689 ();
 sg13g2_decap_8 FILLER_48_1696 ();
 sg13g2_decap_8 FILLER_48_1703 ();
 sg13g2_decap_8 FILLER_48_1710 ();
 sg13g2_decap_8 FILLER_48_1717 ();
 sg13g2_decap_8 FILLER_48_1724 ();
 sg13g2_decap_8 FILLER_48_1731 ();
 sg13g2_decap_8 FILLER_48_1738 ();
 sg13g2_decap_8 FILLER_48_1745 ();
 sg13g2_decap_8 FILLER_48_1752 ();
 sg13g2_decap_8 FILLER_48_1759 ();
 sg13g2_fill_2 FILLER_48_1766 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_4 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_225 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_4 FILLER_49_259 ();
 sg13g2_fill_2 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_293 ();
 sg13g2_decap_8 FILLER_49_300 ();
 sg13g2_decap_4 FILLER_49_307 ();
 sg13g2_fill_1 FILLER_49_311 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_330 ();
 sg13g2_fill_1 FILLER_49_335 ();
 sg13g2_decap_8 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_351 ();
 sg13g2_decap_8 FILLER_49_358 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_fill_2 FILLER_49_417 ();
 sg13g2_fill_1 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_435 ();
 sg13g2_decap_8 FILLER_49_442 ();
 sg13g2_fill_2 FILLER_49_449 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_fill_1 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_fill_1 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_521 ();
 sg13g2_fill_2 FILLER_49_528 ();
 sg13g2_fill_1 FILLER_49_530 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_4 FILLER_49_560 ();
 sg13g2_fill_1 FILLER_49_564 ();
 sg13g2_decap_4 FILLER_49_581 ();
 sg13g2_fill_1 FILLER_49_585 ();
 sg13g2_decap_8 FILLER_49_607 ();
 sg13g2_decap_8 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_621 ();
 sg13g2_decap_8 FILLER_49_628 ();
 sg13g2_decap_8 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_decap_8 FILLER_49_657 ();
 sg13g2_decap_8 FILLER_49_664 ();
 sg13g2_decap_8 FILLER_49_671 ();
 sg13g2_decap_8 FILLER_49_678 ();
 sg13g2_decap_8 FILLER_49_685 ();
 sg13g2_decap_8 FILLER_49_692 ();
 sg13g2_decap_8 FILLER_49_699 ();
 sg13g2_decap_4 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_715 ();
 sg13g2_decap_8 FILLER_49_722 ();
 sg13g2_fill_2 FILLER_49_729 ();
 sg13g2_fill_1 FILLER_49_731 ();
 sg13g2_decap_8 FILLER_49_751 ();
 sg13g2_decap_8 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_765 ();
 sg13g2_decap_8 FILLER_49_772 ();
 sg13g2_decap_8 FILLER_49_779 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_decap_4 FILLER_49_793 ();
 sg13g2_fill_1 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_807 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_8 FILLER_49_856 ();
 sg13g2_decap_8 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_870 ();
 sg13g2_decap_8 FILLER_49_877 ();
 sg13g2_decap_8 FILLER_49_884 ();
 sg13g2_decap_8 FILLER_49_891 ();
 sg13g2_decap_8 FILLER_49_898 ();
 sg13g2_fill_2 FILLER_49_912 ();
 sg13g2_fill_1 FILLER_49_914 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_4 FILLER_49_959 ();
 sg13g2_fill_1 FILLER_49_963 ();
 sg13g2_fill_2 FILLER_49_984 ();
 sg13g2_fill_1 FILLER_49_986 ();
 sg13g2_decap_8 FILLER_49_999 ();
 sg13g2_decap_8 FILLER_49_1006 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_decap_8 FILLER_49_1020 ();
 sg13g2_decap_8 FILLER_49_1027 ();
 sg13g2_decap_8 FILLER_49_1034 ();
 sg13g2_fill_1 FILLER_49_1041 ();
 sg13g2_decap_4 FILLER_49_1046 ();
 sg13g2_decap_8 FILLER_49_1055 ();
 sg13g2_decap_8 FILLER_49_1062 ();
 sg13g2_decap_8 FILLER_49_1069 ();
 sg13g2_fill_2 FILLER_49_1097 ();
 sg13g2_fill_1 FILLER_49_1099 ();
 sg13g2_decap_8 FILLER_49_1150 ();
 sg13g2_decap_8 FILLER_49_1157 ();
 sg13g2_decap_8 FILLER_49_1164 ();
 sg13g2_decap_8 FILLER_49_1171 ();
 sg13g2_fill_2 FILLER_49_1178 ();
 sg13g2_decap_4 FILLER_49_1184 ();
 sg13g2_fill_1 FILLER_49_1188 ();
 sg13g2_fill_1 FILLER_49_1214 ();
 sg13g2_decap_8 FILLER_49_1240 ();
 sg13g2_decap_4 FILLER_49_1247 ();
 sg13g2_decap_8 FILLER_49_1259 ();
 sg13g2_decap_8 FILLER_49_1266 ();
 sg13g2_decap_4 FILLER_49_1273 ();
 sg13g2_fill_1 FILLER_49_1280 ();
 sg13g2_fill_1 FILLER_49_1286 ();
 sg13g2_decap_4 FILLER_49_1312 ();
 sg13g2_fill_1 FILLER_49_1316 ();
 sg13g2_decap_4 FILLER_49_1329 ();
 sg13g2_fill_1 FILLER_49_1333 ();
 sg13g2_decap_8 FILLER_49_1350 ();
 sg13g2_fill_1 FILLER_49_1357 ();
 sg13g2_fill_2 FILLER_49_1377 ();
 sg13g2_fill_1 FILLER_49_1379 ();
 sg13g2_decap_8 FILLER_49_1388 ();
 sg13g2_decap_4 FILLER_49_1395 ();
 sg13g2_decap_8 FILLER_49_1407 ();
 sg13g2_decap_4 FILLER_49_1414 ();
 sg13g2_fill_1 FILLER_49_1418 ();
 sg13g2_decap_8 FILLER_49_1422 ();
 sg13g2_decap_8 FILLER_49_1429 ();
 sg13g2_decap_8 FILLER_49_1436 ();
 sg13g2_fill_1 FILLER_49_1443 ();
 sg13g2_decap_8 FILLER_49_1454 ();
 sg13g2_decap_8 FILLER_49_1461 ();
 sg13g2_fill_1 FILLER_49_1468 ();
 sg13g2_decap_8 FILLER_49_1474 ();
 sg13g2_decap_8 FILLER_49_1481 ();
 sg13g2_decap_8 FILLER_49_1488 ();
 sg13g2_fill_1 FILLER_49_1495 ();
 sg13g2_decap_8 FILLER_49_1513 ();
 sg13g2_decap_8 FILLER_49_1520 ();
 sg13g2_decap_8 FILLER_49_1527 ();
 sg13g2_decap_8 FILLER_49_1534 ();
 sg13g2_decap_8 FILLER_49_1541 ();
 sg13g2_decap_8 FILLER_49_1548 ();
 sg13g2_fill_1 FILLER_49_1555 ();
 sg13g2_fill_2 FILLER_49_1560 ();
 sg13g2_fill_2 FILLER_49_1566 ();
 sg13g2_decap_8 FILLER_49_1576 ();
 sg13g2_decap_8 FILLER_49_1583 ();
 sg13g2_decap_8 FILLER_49_1590 ();
 sg13g2_decap_8 FILLER_49_1597 ();
 sg13g2_decap_8 FILLER_49_1604 ();
 sg13g2_decap_8 FILLER_49_1611 ();
 sg13g2_decap_8 FILLER_49_1618 ();
 sg13g2_decap_8 FILLER_49_1625 ();
 sg13g2_decap_8 FILLER_49_1632 ();
 sg13g2_decap_8 FILLER_49_1639 ();
 sg13g2_decap_8 FILLER_49_1646 ();
 sg13g2_decap_8 FILLER_49_1653 ();
 sg13g2_decap_8 FILLER_49_1660 ();
 sg13g2_decap_8 FILLER_49_1667 ();
 sg13g2_decap_8 FILLER_49_1674 ();
 sg13g2_decap_8 FILLER_49_1681 ();
 sg13g2_decap_8 FILLER_49_1688 ();
 sg13g2_decap_8 FILLER_49_1695 ();
 sg13g2_decap_8 FILLER_49_1702 ();
 sg13g2_decap_8 FILLER_49_1709 ();
 sg13g2_decap_8 FILLER_49_1716 ();
 sg13g2_decap_8 FILLER_49_1723 ();
 sg13g2_decap_8 FILLER_49_1730 ();
 sg13g2_decap_8 FILLER_49_1737 ();
 sg13g2_decap_8 FILLER_49_1744 ();
 sg13g2_decap_8 FILLER_49_1751 ();
 sg13g2_decap_8 FILLER_49_1758 ();
 sg13g2_fill_2 FILLER_49_1765 ();
 sg13g2_fill_1 FILLER_49_1767 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_4 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_212 ();
 sg13g2_decap_8 FILLER_50_230 ();
 sg13g2_decap_8 FILLER_50_237 ();
 sg13g2_decap_8 FILLER_50_244 ();
 sg13g2_decap_8 FILLER_50_251 ();
 sg13g2_decap_8 FILLER_50_258 ();
 sg13g2_decap_8 FILLER_50_272 ();
 sg13g2_decap_8 FILLER_50_279 ();
 sg13g2_decap_8 FILLER_50_286 ();
 sg13g2_decap_8 FILLER_50_293 ();
 sg13g2_decap_8 FILLER_50_300 ();
 sg13g2_decap_8 FILLER_50_307 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_decap_8 FILLER_50_353 ();
 sg13g2_decap_4 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_372 ();
 sg13g2_decap_4 FILLER_50_382 ();
 sg13g2_fill_1 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_8 FILLER_50_405 ();
 sg13g2_fill_2 FILLER_50_412 ();
 sg13g2_fill_1 FILLER_50_414 ();
 sg13g2_decap_8 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_50_435 ();
 sg13g2_decap_8 FILLER_50_442 ();
 sg13g2_decap_4 FILLER_50_449 ();
 sg13g2_fill_1 FILLER_50_453 ();
 sg13g2_decap_8 FILLER_50_472 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_decap_8 FILLER_50_486 ();
 sg13g2_decap_8 FILLER_50_493 ();
 sg13g2_decap_8 FILLER_50_500 ();
 sg13g2_decap_8 FILLER_50_507 ();
 sg13g2_fill_2 FILLER_50_514 ();
 sg13g2_fill_1 FILLER_50_516 ();
 sg13g2_decap_4 FILLER_50_521 ();
 sg13g2_fill_2 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_545 ();
 sg13g2_decap_8 FILLER_50_552 ();
 sg13g2_decap_8 FILLER_50_559 ();
 sg13g2_decap_4 FILLER_50_566 ();
 sg13g2_fill_1 FILLER_50_570 ();
 sg13g2_fill_2 FILLER_50_593 ();
 sg13g2_decap_8 FILLER_50_603 ();
 sg13g2_decap_4 FILLER_50_610 ();
 sg13g2_fill_1 FILLER_50_614 ();
 sg13g2_decap_8 FILLER_50_632 ();
 sg13g2_decap_8 FILLER_50_639 ();
 sg13g2_decap_8 FILLER_50_646 ();
 sg13g2_decap_8 FILLER_50_653 ();
 sg13g2_decap_8 FILLER_50_660 ();
 sg13g2_decap_8 FILLER_50_667 ();
 sg13g2_decap_8 FILLER_50_674 ();
 sg13g2_decap_8 FILLER_50_681 ();
 sg13g2_decap_8 FILLER_50_688 ();
 sg13g2_decap_8 FILLER_50_695 ();
 sg13g2_decap_4 FILLER_50_702 ();
 sg13g2_fill_1 FILLER_50_714 ();
 sg13g2_decap_8 FILLER_50_723 ();
 sg13g2_fill_2 FILLER_50_730 ();
 sg13g2_fill_1 FILLER_50_732 ();
 sg13g2_decap_4 FILLER_50_746 ();
 sg13g2_fill_1 FILLER_50_750 ();
 sg13g2_decap_8 FILLER_50_761 ();
 sg13g2_decap_8 FILLER_50_768 ();
 sg13g2_decap_4 FILLER_50_775 ();
 sg13g2_fill_2 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_797 ();
 sg13g2_decap_8 FILLER_50_804 ();
 sg13g2_decap_8 FILLER_50_811 ();
 sg13g2_decap_8 FILLER_50_818 ();
 sg13g2_fill_1 FILLER_50_825 ();
 sg13g2_decap_4 FILLER_50_831 ();
 sg13g2_fill_2 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_857 ();
 sg13g2_decap_8 FILLER_50_864 ();
 sg13g2_decap_8 FILLER_50_871 ();
 sg13g2_decap_8 FILLER_50_878 ();
 sg13g2_decap_8 FILLER_50_885 ();
 sg13g2_decap_8 FILLER_50_892 ();
 sg13g2_decap_8 FILLER_50_899 ();
 sg13g2_decap_4 FILLER_50_906 ();
 sg13g2_fill_2 FILLER_50_910 ();
 sg13g2_decap_8 FILLER_50_932 ();
 sg13g2_decap_8 FILLER_50_939 ();
 sg13g2_decap_8 FILLER_50_946 ();
 sg13g2_decap_8 FILLER_50_953 ();
 sg13g2_fill_2 FILLER_50_960 ();
 sg13g2_decap_4 FILLER_50_967 ();
 sg13g2_decap_8 FILLER_50_994 ();
 sg13g2_decap_8 FILLER_50_1001 ();
 sg13g2_decap_8 FILLER_50_1008 ();
 sg13g2_decap_8 FILLER_50_1015 ();
 sg13g2_decap_8 FILLER_50_1022 ();
 sg13g2_decap_8 FILLER_50_1029 ();
 sg13g2_fill_1 FILLER_50_1036 ();
 sg13g2_fill_1 FILLER_50_1049 ();
 sg13g2_decap_8 FILLER_50_1058 ();
 sg13g2_decap_8 FILLER_50_1065 ();
 sg13g2_decap_8 FILLER_50_1072 ();
 sg13g2_decap_8 FILLER_50_1079 ();
 sg13g2_decap_8 FILLER_50_1086 ();
 sg13g2_fill_2 FILLER_50_1093 ();
 sg13g2_decap_8 FILLER_50_1104 ();
 sg13g2_decap_8 FILLER_50_1111 ();
 sg13g2_decap_8 FILLER_50_1118 ();
 sg13g2_decap_8 FILLER_50_1125 ();
 sg13g2_decap_4 FILLER_50_1132 ();
 sg13g2_decap_8 FILLER_50_1146 ();
 sg13g2_decap_8 FILLER_50_1153 ();
 sg13g2_decap_8 FILLER_50_1160 ();
 sg13g2_decap_8 FILLER_50_1167 ();
 sg13g2_decap_8 FILLER_50_1174 ();
 sg13g2_fill_2 FILLER_50_1181 ();
 sg13g2_fill_1 FILLER_50_1183 ();
 sg13g2_decap_8 FILLER_50_1189 ();
 sg13g2_decap_4 FILLER_50_1213 ();
 sg13g2_fill_2 FILLER_50_1217 ();
 sg13g2_decap_8 FILLER_50_1228 ();
 sg13g2_decap_4 FILLER_50_1235 ();
 sg13g2_fill_2 FILLER_50_1244 ();
 sg13g2_fill_1 FILLER_50_1246 ();
 sg13g2_decap_8 FILLER_50_1259 ();
 sg13g2_decap_4 FILLER_50_1266 ();
 sg13g2_decap_8 FILLER_50_1338 ();
 sg13g2_decap_8 FILLER_50_1345 ();
 sg13g2_decap_8 FILLER_50_1352 ();
 sg13g2_fill_2 FILLER_50_1359 ();
 sg13g2_fill_1 FILLER_50_1361 ();
 sg13g2_decap_4 FILLER_50_1366 ();
 sg13g2_fill_1 FILLER_50_1370 ();
 sg13g2_fill_2 FILLER_50_1383 ();
 sg13g2_decap_8 FILLER_50_1398 ();
 sg13g2_decap_8 FILLER_50_1405 ();
 sg13g2_decap_8 FILLER_50_1412 ();
 sg13g2_decap_8 FILLER_50_1419 ();
 sg13g2_decap_8 FILLER_50_1426 ();
 sg13g2_fill_1 FILLER_50_1433 ();
 sg13g2_fill_1 FILLER_50_1442 ();
 sg13g2_decap_4 FILLER_50_1465 ();
 sg13g2_decap_8 FILLER_50_1484 ();
 sg13g2_decap_8 FILLER_50_1491 ();
 sg13g2_fill_1 FILLER_50_1498 ();
 sg13g2_fill_2 FILLER_50_1503 ();
 sg13g2_fill_1 FILLER_50_1505 ();
 sg13g2_decap_8 FILLER_50_1514 ();
 sg13g2_decap_8 FILLER_50_1521 ();
 sg13g2_decap_4 FILLER_50_1528 ();
 sg13g2_decap_4 FILLER_50_1537 ();
 sg13g2_fill_2 FILLER_50_1541 ();
 sg13g2_decap_8 FILLER_50_1551 ();
 sg13g2_decap_8 FILLER_50_1558 ();
 sg13g2_decap_8 FILLER_50_1565 ();
 sg13g2_decap_8 FILLER_50_1572 ();
 sg13g2_decap_8 FILLER_50_1579 ();
 sg13g2_decap_8 FILLER_50_1586 ();
 sg13g2_decap_8 FILLER_50_1593 ();
 sg13g2_decap_8 FILLER_50_1600 ();
 sg13g2_decap_8 FILLER_50_1607 ();
 sg13g2_decap_8 FILLER_50_1614 ();
 sg13g2_decap_8 FILLER_50_1621 ();
 sg13g2_decap_8 FILLER_50_1628 ();
 sg13g2_decap_8 FILLER_50_1635 ();
 sg13g2_decap_8 FILLER_50_1642 ();
 sg13g2_decap_8 FILLER_50_1649 ();
 sg13g2_decap_8 FILLER_50_1656 ();
 sg13g2_decap_8 FILLER_50_1663 ();
 sg13g2_decap_8 FILLER_50_1670 ();
 sg13g2_decap_8 FILLER_50_1677 ();
 sg13g2_decap_8 FILLER_50_1684 ();
 sg13g2_decap_8 FILLER_50_1691 ();
 sg13g2_decap_8 FILLER_50_1698 ();
 sg13g2_decap_8 FILLER_50_1705 ();
 sg13g2_decap_8 FILLER_50_1712 ();
 sg13g2_decap_8 FILLER_50_1719 ();
 sg13g2_decap_8 FILLER_50_1726 ();
 sg13g2_decap_8 FILLER_50_1733 ();
 sg13g2_decap_8 FILLER_50_1740 ();
 sg13g2_decap_8 FILLER_50_1747 ();
 sg13g2_decap_8 FILLER_50_1754 ();
 sg13g2_decap_8 FILLER_50_1761 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_fill_2 FILLER_51_196 ();
 sg13g2_fill_2 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_205 ();
 sg13g2_decap_8 FILLER_51_221 ();
 sg13g2_decap_8 FILLER_51_228 ();
 sg13g2_decap_8 FILLER_51_235 ();
 sg13g2_decap_8 FILLER_51_242 ();
 sg13g2_decap_8 FILLER_51_249 ();
 sg13g2_decap_8 FILLER_51_256 ();
 sg13g2_decap_8 FILLER_51_263 ();
 sg13g2_decap_4 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_274 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_decap_8 FILLER_51_288 ();
 sg13g2_decap_8 FILLER_51_295 ();
 sg13g2_decap_4 FILLER_51_302 ();
 sg13g2_decap_8 FILLER_51_310 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_fill_1 FILLER_51_330 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_337 ();
 sg13g2_fill_2 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_349 ();
 sg13g2_decap_8 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_377 ();
 sg13g2_decap_8 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_391 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_decap_8 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_51_415 ();
 sg13g2_decap_4 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_51_432 ();
 sg13g2_fill_1 FILLER_51_434 ();
 sg13g2_fill_1 FILLER_51_439 ();
 sg13g2_decap_8 FILLER_51_457 ();
 sg13g2_decap_8 FILLER_51_464 ();
 sg13g2_decap_8 FILLER_51_471 ();
 sg13g2_decap_4 FILLER_51_478 ();
 sg13g2_decap_8 FILLER_51_486 ();
 sg13g2_decap_8 FILLER_51_493 ();
 sg13g2_decap_8 FILLER_51_500 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_decap_4 FILLER_51_514 ();
 sg13g2_decap_4 FILLER_51_541 ();
 sg13g2_fill_1 FILLER_51_545 ();
 sg13g2_decap_8 FILLER_51_554 ();
 sg13g2_decap_8 FILLER_51_569 ();
 sg13g2_decap_8 FILLER_51_576 ();
 sg13g2_decap_8 FILLER_51_583 ();
 sg13g2_decap_8 FILLER_51_590 ();
 sg13g2_decap_8 FILLER_51_597 ();
 sg13g2_decap_8 FILLER_51_636 ();
 sg13g2_decap_8 FILLER_51_643 ();
 sg13g2_decap_8 FILLER_51_650 ();
 sg13g2_decap_8 FILLER_51_657 ();
 sg13g2_decap_8 FILLER_51_664 ();
 sg13g2_decap_8 FILLER_51_671 ();
 sg13g2_decap_8 FILLER_51_682 ();
 sg13g2_decap_8 FILLER_51_689 ();
 sg13g2_decap_8 FILLER_51_696 ();
 sg13g2_decap_4 FILLER_51_703 ();
 sg13g2_decap_8 FILLER_51_714 ();
 sg13g2_decap_8 FILLER_51_721 ();
 sg13g2_decap_8 FILLER_51_728 ();
 sg13g2_decap_8 FILLER_51_735 ();
 sg13g2_decap_8 FILLER_51_742 ();
 sg13g2_decap_8 FILLER_51_749 ();
 sg13g2_decap_8 FILLER_51_756 ();
 sg13g2_decap_8 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_770 ();
 sg13g2_decap_8 FILLER_51_777 ();
 sg13g2_decap_8 FILLER_51_784 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_decap_8 FILLER_51_812 ();
 sg13g2_fill_2 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_863 ();
 sg13g2_decap_8 FILLER_51_870 ();
 sg13g2_decap_8 FILLER_51_877 ();
 sg13g2_fill_1 FILLER_51_884 ();
 sg13g2_decap_8 FILLER_51_901 ();
 sg13g2_fill_2 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_921 ();
 sg13g2_fill_1 FILLER_51_931 ();
 sg13g2_decap_8 FILLER_51_935 ();
 sg13g2_decap_8 FILLER_51_942 ();
 sg13g2_decap_8 FILLER_51_949 ();
 sg13g2_decap_4 FILLER_51_956 ();
 sg13g2_fill_1 FILLER_51_960 ();
 sg13g2_decap_8 FILLER_51_965 ();
 sg13g2_decap_8 FILLER_51_977 ();
 sg13g2_decap_8 FILLER_51_984 ();
 sg13g2_decap_8 FILLER_51_991 ();
 sg13g2_decap_8 FILLER_51_998 ();
 sg13g2_decap_8 FILLER_51_1013 ();
 sg13g2_decap_8 FILLER_51_1020 ();
 sg13g2_decap_4 FILLER_51_1027 ();
 sg13g2_fill_2 FILLER_51_1031 ();
 sg13g2_decap_8 FILLER_51_1057 ();
 sg13g2_decap_8 FILLER_51_1064 ();
 sg13g2_decap_8 FILLER_51_1071 ();
 sg13g2_decap_8 FILLER_51_1078 ();
 sg13g2_decap_8 FILLER_51_1085 ();
 sg13g2_decap_8 FILLER_51_1092 ();
 sg13g2_decap_4 FILLER_51_1099 ();
 sg13g2_fill_1 FILLER_51_1103 ();
 sg13g2_decap_8 FILLER_51_1113 ();
 sg13g2_decap_8 FILLER_51_1120 ();
 sg13g2_decap_8 FILLER_51_1127 ();
 sg13g2_fill_1 FILLER_51_1134 ();
 sg13g2_fill_2 FILLER_51_1143 ();
 sg13g2_decap_8 FILLER_51_1150 ();
 sg13g2_decap_8 FILLER_51_1157 ();
 sg13g2_decap_8 FILLER_51_1164 ();
 sg13g2_decap_8 FILLER_51_1171 ();
 sg13g2_decap_8 FILLER_51_1178 ();
 sg13g2_decap_8 FILLER_51_1185 ();
 sg13g2_decap_8 FILLER_51_1192 ();
 sg13g2_decap_8 FILLER_51_1199 ();
 sg13g2_decap_8 FILLER_51_1206 ();
 sg13g2_decap_8 FILLER_51_1213 ();
 sg13g2_decap_8 FILLER_51_1220 ();
 sg13g2_fill_2 FILLER_51_1227 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1271 ();
 sg13g2_decap_4 FILLER_51_1282 ();
 sg13g2_fill_2 FILLER_51_1286 ();
 sg13g2_decap_8 FILLER_51_1307 ();
 sg13g2_decap_8 FILLER_51_1314 ();
 sg13g2_decap_4 FILLER_51_1321 ();
 sg13g2_decap_8 FILLER_51_1329 ();
 sg13g2_decap_8 FILLER_51_1336 ();
 sg13g2_decap_8 FILLER_51_1343 ();
 sg13g2_decap_8 FILLER_51_1350 ();
 sg13g2_decap_8 FILLER_51_1357 ();
 sg13g2_decap_8 FILLER_51_1364 ();
 sg13g2_decap_4 FILLER_51_1371 ();
 sg13g2_fill_2 FILLER_51_1375 ();
 sg13g2_decap_8 FILLER_51_1384 ();
 sg13g2_decap_8 FILLER_51_1391 ();
 sg13g2_decap_8 FILLER_51_1398 ();
 sg13g2_decap_8 FILLER_51_1405 ();
 sg13g2_decap_8 FILLER_51_1412 ();
 sg13g2_decap_8 FILLER_51_1419 ();
 sg13g2_decap_8 FILLER_51_1426 ();
 sg13g2_decap_8 FILLER_51_1433 ();
 sg13g2_decap_4 FILLER_51_1440 ();
 sg13g2_fill_2 FILLER_51_1444 ();
 sg13g2_decap_8 FILLER_51_1450 ();
 sg13g2_decap_8 FILLER_51_1457 ();
 sg13g2_decap_4 FILLER_51_1464 ();
 sg13g2_fill_2 FILLER_51_1468 ();
 sg13g2_decap_8 FILLER_51_1479 ();
 sg13g2_fill_2 FILLER_51_1486 ();
 sg13g2_fill_1 FILLER_51_1488 ();
 sg13g2_decap_8 FILLER_51_1493 ();
 sg13g2_decap_8 FILLER_51_1500 ();
 sg13g2_decap_8 FILLER_51_1507 ();
 sg13g2_decap_8 FILLER_51_1514 ();
 sg13g2_decap_8 FILLER_51_1521 ();
 sg13g2_fill_1 FILLER_51_1528 ();
 sg13g2_decap_8 FILLER_51_1555 ();
 sg13g2_decap_8 FILLER_51_1562 ();
 sg13g2_decap_8 FILLER_51_1569 ();
 sg13g2_decap_8 FILLER_51_1576 ();
 sg13g2_decap_8 FILLER_51_1583 ();
 sg13g2_decap_8 FILLER_51_1590 ();
 sg13g2_decap_8 FILLER_51_1597 ();
 sg13g2_decap_8 FILLER_51_1604 ();
 sg13g2_decap_8 FILLER_51_1611 ();
 sg13g2_decap_8 FILLER_51_1618 ();
 sg13g2_decap_8 FILLER_51_1625 ();
 sg13g2_decap_8 FILLER_51_1632 ();
 sg13g2_decap_8 FILLER_51_1639 ();
 sg13g2_decap_8 FILLER_51_1646 ();
 sg13g2_decap_8 FILLER_51_1653 ();
 sg13g2_decap_8 FILLER_51_1660 ();
 sg13g2_decap_8 FILLER_51_1667 ();
 sg13g2_decap_8 FILLER_51_1674 ();
 sg13g2_decap_8 FILLER_51_1681 ();
 sg13g2_decap_8 FILLER_51_1688 ();
 sg13g2_decap_8 FILLER_51_1695 ();
 sg13g2_decap_8 FILLER_51_1702 ();
 sg13g2_decap_8 FILLER_51_1709 ();
 sg13g2_decap_8 FILLER_51_1716 ();
 sg13g2_decap_8 FILLER_51_1723 ();
 sg13g2_decap_8 FILLER_51_1730 ();
 sg13g2_decap_8 FILLER_51_1737 ();
 sg13g2_decap_8 FILLER_51_1744 ();
 sg13g2_decap_8 FILLER_51_1751 ();
 sg13g2_decap_8 FILLER_51_1758 ();
 sg13g2_fill_2 FILLER_51_1765 ();
 sg13g2_fill_1 FILLER_51_1767 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_276 ();
 sg13g2_decap_8 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_290 ();
 sg13g2_decap_8 FILLER_52_297 ();
 sg13g2_decap_8 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_decap_8 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_decap_8 FILLER_52_332 ();
 sg13g2_decap_8 FILLER_52_339 ();
 sg13g2_decap_8 FILLER_52_346 ();
 sg13g2_decap_8 FILLER_52_353 ();
 sg13g2_decap_8 FILLER_52_360 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_374 ();
 sg13g2_decap_4 FILLER_52_379 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_4 FILLER_52_420 ();
 sg13g2_fill_1 FILLER_52_447 ();
 sg13g2_decap_8 FILLER_52_456 ();
 sg13g2_decap_8 FILLER_52_463 ();
 sg13g2_fill_2 FILLER_52_470 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_fill_2 FILLER_52_504 ();
 sg13g2_decap_8 FILLER_52_510 ();
 sg13g2_decap_8 FILLER_52_517 ();
 sg13g2_decap_8 FILLER_52_524 ();
 sg13g2_decap_8 FILLER_52_531 ();
 sg13g2_decap_8 FILLER_52_538 ();
 sg13g2_decap_8 FILLER_52_545 ();
 sg13g2_decap_8 FILLER_52_552 ();
 sg13g2_decap_8 FILLER_52_559 ();
 sg13g2_decap_4 FILLER_52_566 ();
 sg13g2_fill_1 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_576 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_fill_2 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_fill_1 FILLER_52_614 ();
 sg13g2_fill_2 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_624 ();
 sg13g2_decap_8 FILLER_52_631 ();
 sg13g2_decap_8 FILLER_52_638 ();
 sg13g2_decap_8 FILLER_52_645 ();
 sg13g2_decap_8 FILLER_52_652 ();
 sg13g2_decap_8 FILLER_52_659 ();
 sg13g2_decap_8 FILLER_52_699 ();
 sg13g2_decap_8 FILLER_52_706 ();
 sg13g2_decap_8 FILLER_52_713 ();
 sg13g2_decap_8 FILLER_52_720 ();
 sg13g2_decap_8 FILLER_52_727 ();
 sg13g2_decap_4 FILLER_52_734 ();
 sg13g2_fill_2 FILLER_52_738 ();
 sg13g2_decap_8 FILLER_52_744 ();
 sg13g2_decap_8 FILLER_52_751 ();
 sg13g2_decap_8 FILLER_52_758 ();
 sg13g2_decap_8 FILLER_52_765 ();
 sg13g2_decap_4 FILLER_52_772 ();
 sg13g2_fill_2 FILLER_52_776 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_decap_8 FILLER_52_793 ();
 sg13g2_fill_1 FILLER_52_800 ();
 sg13g2_decap_8 FILLER_52_810 ();
 sg13g2_decap_8 FILLER_52_817 ();
 sg13g2_decap_8 FILLER_52_824 ();
 sg13g2_fill_2 FILLER_52_831 ();
 sg13g2_fill_1 FILLER_52_833 ();
 sg13g2_fill_2 FILLER_52_838 ();
 sg13g2_decap_8 FILLER_52_856 ();
 sg13g2_decap_8 FILLER_52_863 ();
 sg13g2_decap_8 FILLER_52_870 ();
 sg13g2_decap_8 FILLER_52_877 ();
 sg13g2_fill_2 FILLER_52_884 ();
 sg13g2_decap_4 FILLER_52_890 ();
 sg13g2_fill_2 FILLER_52_902 ();
 sg13g2_fill_1 FILLER_52_904 ();
 sg13g2_decap_8 FILLER_52_913 ();
 sg13g2_decap_8 FILLER_52_920 ();
 sg13g2_decap_8 FILLER_52_927 ();
 sg13g2_decap_4 FILLER_52_934 ();
 sg13g2_fill_1 FILLER_52_938 ();
 sg13g2_decap_8 FILLER_52_943 ();
 sg13g2_decap_8 FILLER_52_950 ();
 sg13g2_decap_8 FILLER_52_957 ();
 sg13g2_decap_8 FILLER_52_964 ();
 sg13g2_decap_8 FILLER_52_971 ();
 sg13g2_decap_8 FILLER_52_978 ();
 sg13g2_decap_8 FILLER_52_985 ();
 sg13g2_decap_8 FILLER_52_992 ();
 sg13g2_decap_4 FILLER_52_999 ();
 sg13g2_fill_2 FILLER_52_1003 ();
 sg13g2_decap_8 FILLER_52_1025 ();
 sg13g2_fill_2 FILLER_52_1032 ();
 sg13g2_fill_1 FILLER_52_1034 ();
 sg13g2_decap_4 FILLER_52_1039 ();
 sg13g2_fill_2 FILLER_52_1048 ();
 sg13g2_decap_8 FILLER_52_1058 ();
 sg13g2_decap_8 FILLER_52_1065 ();
 sg13g2_decap_8 FILLER_52_1072 ();
 sg13g2_decap_4 FILLER_52_1079 ();
 sg13g2_fill_2 FILLER_52_1083 ();
 sg13g2_decap_8 FILLER_52_1093 ();
 sg13g2_decap_8 FILLER_52_1100 ();
 sg13g2_decap_8 FILLER_52_1107 ();
 sg13g2_decap_8 FILLER_52_1114 ();
 sg13g2_decap_4 FILLER_52_1121 ();
 sg13g2_decap_8 FILLER_52_1129 ();
 sg13g2_fill_1 FILLER_52_1136 ();
 sg13g2_decap_8 FILLER_52_1161 ();
 sg13g2_decap_8 FILLER_52_1168 ();
 sg13g2_decap_8 FILLER_52_1175 ();
 sg13g2_decap_8 FILLER_52_1182 ();
 sg13g2_decap_8 FILLER_52_1197 ();
 sg13g2_decap_8 FILLER_52_1204 ();
 sg13g2_decap_8 FILLER_52_1211 ();
 sg13g2_decap_8 FILLER_52_1218 ();
 sg13g2_decap_8 FILLER_52_1225 ();
 sg13g2_fill_2 FILLER_52_1232 ();
 sg13g2_fill_1 FILLER_52_1234 ();
 sg13g2_decap_4 FILLER_52_1243 ();
 sg13g2_decap_8 FILLER_52_1262 ();
 sg13g2_decap_8 FILLER_52_1269 ();
 sg13g2_decap_8 FILLER_52_1276 ();
 sg13g2_decap_8 FILLER_52_1283 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_decap_8 FILLER_52_1297 ();
 sg13g2_decap_8 FILLER_52_1304 ();
 sg13g2_decap_8 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_decap_8 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_52_1332 ();
 sg13g2_decap_8 FILLER_52_1339 ();
 sg13g2_decap_8 FILLER_52_1346 ();
 sg13g2_decap_8 FILLER_52_1353 ();
 sg13g2_decap_8 FILLER_52_1360 ();
 sg13g2_decap_8 FILLER_52_1367 ();
 sg13g2_decap_8 FILLER_52_1374 ();
 sg13g2_decap_4 FILLER_52_1381 ();
 sg13g2_fill_2 FILLER_52_1385 ();
 sg13g2_decap_4 FILLER_52_1392 ();
 sg13g2_fill_1 FILLER_52_1401 ();
 sg13g2_decap_8 FILLER_52_1406 ();
 sg13g2_decap_8 FILLER_52_1413 ();
 sg13g2_decap_8 FILLER_52_1420 ();
 sg13g2_decap_4 FILLER_52_1427 ();
 sg13g2_decap_8 FILLER_52_1440 ();
 sg13g2_decap_8 FILLER_52_1447 ();
 sg13g2_decap_8 FILLER_52_1454 ();
 sg13g2_decap_8 FILLER_52_1461 ();
 sg13g2_decap_8 FILLER_52_1468 ();
 sg13g2_decap_8 FILLER_52_1475 ();
 sg13g2_fill_1 FILLER_52_1482 ();
 sg13g2_decap_8 FILLER_52_1503 ();
 sg13g2_decap_8 FILLER_52_1510 ();
 sg13g2_decap_8 FILLER_52_1517 ();
 sg13g2_decap_8 FILLER_52_1524 ();
 sg13g2_decap_8 FILLER_52_1531 ();
 sg13g2_decap_8 FILLER_52_1538 ();
 sg13g2_decap_4 FILLER_52_1545 ();
 sg13g2_fill_2 FILLER_52_1549 ();
 sg13g2_fill_2 FILLER_52_1563 ();
 sg13g2_fill_1 FILLER_52_1565 ();
 sg13g2_decap_8 FILLER_52_1571 ();
 sg13g2_decap_8 FILLER_52_1578 ();
 sg13g2_decap_8 FILLER_52_1585 ();
 sg13g2_decap_8 FILLER_52_1592 ();
 sg13g2_decap_8 FILLER_52_1599 ();
 sg13g2_decap_8 FILLER_52_1606 ();
 sg13g2_decap_8 FILLER_52_1613 ();
 sg13g2_decap_8 FILLER_52_1620 ();
 sg13g2_decap_8 FILLER_52_1627 ();
 sg13g2_decap_8 FILLER_52_1634 ();
 sg13g2_decap_8 FILLER_52_1641 ();
 sg13g2_decap_8 FILLER_52_1648 ();
 sg13g2_decap_8 FILLER_52_1655 ();
 sg13g2_decap_8 FILLER_52_1662 ();
 sg13g2_decap_8 FILLER_52_1669 ();
 sg13g2_decap_8 FILLER_52_1676 ();
 sg13g2_decap_8 FILLER_52_1683 ();
 sg13g2_decap_8 FILLER_52_1690 ();
 sg13g2_decap_8 FILLER_52_1697 ();
 sg13g2_decap_8 FILLER_52_1704 ();
 sg13g2_decap_8 FILLER_52_1711 ();
 sg13g2_decap_8 FILLER_52_1718 ();
 sg13g2_decap_8 FILLER_52_1725 ();
 sg13g2_decap_8 FILLER_52_1732 ();
 sg13g2_decap_8 FILLER_52_1739 ();
 sg13g2_decap_8 FILLER_52_1746 ();
 sg13g2_decap_8 FILLER_52_1753 ();
 sg13g2_decap_8 FILLER_52_1760 ();
 sg13g2_fill_1 FILLER_52_1767 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_4 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_8 FILLER_53_218 ();
 sg13g2_decap_8 FILLER_53_225 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_8 FILLER_53_246 ();
 sg13g2_decap_8 FILLER_53_253 ();
 sg13g2_decap_8 FILLER_53_260 ();
 sg13g2_decap_4 FILLER_53_267 ();
 sg13g2_fill_2 FILLER_53_271 ();
 sg13g2_decap_4 FILLER_53_277 ();
 sg13g2_decap_8 FILLER_53_284 ();
 sg13g2_fill_2 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_decap_8 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_decap_8 FILLER_53_337 ();
 sg13g2_decap_8 FILLER_53_344 ();
 sg13g2_decap_8 FILLER_53_351 ();
 sg13g2_decap_8 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_decap_8 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_decap_8 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_53_414 ();
 sg13g2_decap_8 FILLER_53_421 ();
 sg13g2_decap_8 FILLER_53_428 ();
 sg13g2_fill_2 FILLER_53_435 ();
 sg13g2_decap_8 FILLER_53_449 ();
 sg13g2_decap_8 FILLER_53_456 ();
 sg13g2_fill_1 FILLER_53_463 ();
 sg13g2_decap_8 FILLER_53_473 ();
 sg13g2_decap_8 FILLER_53_480 ();
 sg13g2_fill_2 FILLER_53_487 ();
 sg13g2_fill_1 FILLER_53_489 ();
 sg13g2_decap_4 FILLER_53_495 ();
 sg13g2_fill_1 FILLER_53_499 ();
 sg13g2_decap_8 FILLER_53_516 ();
 sg13g2_decap_8 FILLER_53_523 ();
 sg13g2_decap_8 FILLER_53_530 ();
 sg13g2_decap_8 FILLER_53_537 ();
 sg13g2_decap_8 FILLER_53_544 ();
 sg13g2_decap_4 FILLER_53_551 ();
 sg13g2_fill_1 FILLER_53_555 ();
 sg13g2_decap_4 FILLER_53_559 ();
 sg13g2_fill_1 FILLER_53_563 ();
 sg13g2_decap_8 FILLER_53_567 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_581 ();
 sg13g2_decap_8 FILLER_53_588 ();
 sg13g2_decap_8 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_602 ();
 sg13g2_fill_2 FILLER_53_609 ();
 sg13g2_fill_2 FILLER_53_619 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_8 FILLER_53_651 ();
 sg13g2_decap_4 FILLER_53_658 ();
 sg13g2_decap_4 FILLER_53_670 ();
 sg13g2_fill_2 FILLER_53_674 ();
 sg13g2_decap_8 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_693 ();
 sg13g2_decap_8 FILLER_53_700 ();
 sg13g2_decap_4 FILLER_53_707 ();
 sg13g2_fill_1 FILLER_53_711 ();
 sg13g2_fill_2 FILLER_53_717 ();
 sg13g2_fill_1 FILLER_53_719 ();
 sg13g2_fill_1 FILLER_53_728 ();
 sg13g2_decap_4 FILLER_53_751 ();
 sg13g2_fill_2 FILLER_53_755 ();
 sg13g2_fill_1 FILLER_53_778 ();
 sg13g2_decap_8 FILLER_53_799 ();
 sg13g2_decap_8 FILLER_53_806 ();
 sg13g2_fill_2 FILLER_53_813 ();
 sg13g2_fill_1 FILLER_53_815 ();
 sg13g2_fill_2 FILLER_53_824 ();
 sg13g2_fill_1 FILLER_53_826 ();
 sg13g2_decap_4 FILLER_53_833 ();
 sg13g2_fill_2 FILLER_53_837 ();
 sg13g2_decap_8 FILLER_53_856 ();
 sg13g2_decap_8 FILLER_53_863 ();
 sg13g2_decap_8 FILLER_53_870 ();
 sg13g2_decap_8 FILLER_53_877 ();
 sg13g2_decap_8 FILLER_53_884 ();
 sg13g2_decap_8 FILLER_53_918 ();
 sg13g2_decap_8 FILLER_53_925 ();
 sg13g2_decap_4 FILLER_53_932 ();
 sg13g2_fill_2 FILLER_53_936 ();
 sg13g2_decap_8 FILLER_53_942 ();
 sg13g2_decap_4 FILLER_53_949 ();
 sg13g2_decap_4 FILLER_53_961 ();
 sg13g2_decap_8 FILLER_53_969 ();
 sg13g2_decap_8 FILLER_53_976 ();
 sg13g2_decap_8 FILLER_53_983 ();
 sg13g2_decap_8 FILLER_53_990 ();
 sg13g2_decap_8 FILLER_53_997 ();
 sg13g2_decap_8 FILLER_53_1004 ();
 sg13g2_decap_8 FILLER_53_1016 ();
 sg13g2_decap_8 FILLER_53_1023 ();
 sg13g2_decap_8 FILLER_53_1030 ();
 sg13g2_decap_8 FILLER_53_1037 ();
 sg13g2_decap_8 FILLER_53_1044 ();
 sg13g2_decap_8 FILLER_53_1051 ();
 sg13g2_decap_8 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_decap_4 FILLER_53_1072 ();
 sg13g2_fill_2 FILLER_53_1076 ();
 sg13g2_decap_8 FILLER_53_1099 ();
 sg13g2_decap_8 FILLER_53_1106 ();
 sg13g2_decap_8 FILLER_53_1113 ();
 sg13g2_decap_8 FILLER_53_1120 ();
 sg13g2_decap_8 FILLER_53_1127 ();
 sg13g2_decap_8 FILLER_53_1134 ();
 sg13g2_decap_4 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1150 ();
 sg13g2_decap_8 FILLER_53_1157 ();
 sg13g2_decap_8 FILLER_53_1164 ();
 sg13g2_fill_2 FILLER_53_1171 ();
 sg13g2_fill_1 FILLER_53_1173 ();
 sg13g2_decap_8 FILLER_53_1200 ();
 sg13g2_decap_8 FILLER_53_1207 ();
 sg13g2_decap_8 FILLER_53_1214 ();
 sg13g2_fill_2 FILLER_53_1221 ();
 sg13g2_fill_1 FILLER_53_1223 ();
 sg13g2_fill_2 FILLER_53_1233 ();
 sg13g2_fill_1 FILLER_53_1240 ();
 sg13g2_decap_8 FILLER_53_1255 ();
 sg13g2_decap_8 FILLER_53_1262 ();
 sg13g2_decap_8 FILLER_53_1269 ();
 sg13g2_decap_8 FILLER_53_1276 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_decap_8 FILLER_53_1290 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_decap_8 FILLER_53_1304 ();
 sg13g2_decap_4 FILLER_53_1311 ();
 sg13g2_fill_2 FILLER_53_1315 ();
 sg13g2_decap_8 FILLER_53_1321 ();
 sg13g2_decap_8 FILLER_53_1333 ();
 sg13g2_decap_8 FILLER_53_1340 ();
 sg13g2_decap_8 FILLER_53_1347 ();
 sg13g2_decap_8 FILLER_53_1354 ();
 sg13g2_decap_8 FILLER_53_1361 ();
 sg13g2_decap_8 FILLER_53_1368 ();
 sg13g2_fill_2 FILLER_53_1375 ();
 sg13g2_fill_1 FILLER_53_1377 ();
 sg13g2_decap_8 FILLER_53_1412 ();
 sg13g2_decap_8 FILLER_53_1419 ();
 sg13g2_decap_8 FILLER_53_1426 ();
 sg13g2_decap_4 FILLER_53_1433 ();
 sg13g2_fill_2 FILLER_53_1437 ();
 sg13g2_decap_8 FILLER_53_1447 ();
 sg13g2_decap_8 FILLER_53_1454 ();
 sg13g2_decap_8 FILLER_53_1461 ();
 sg13g2_fill_2 FILLER_53_1468 ();
 sg13g2_fill_2 FILLER_53_1479 ();
 sg13g2_decap_8 FILLER_53_1491 ();
 sg13g2_decap_8 FILLER_53_1498 ();
 sg13g2_decap_8 FILLER_53_1505 ();
 sg13g2_fill_2 FILLER_53_1512 ();
 sg13g2_fill_1 FILLER_53_1514 ();
 sg13g2_decap_8 FILLER_53_1520 ();
 sg13g2_fill_1 FILLER_53_1527 ();
 sg13g2_decap_8 FILLER_53_1541 ();
 sg13g2_decap_8 FILLER_53_1548 ();
 sg13g2_decap_4 FILLER_53_1555 ();
 sg13g2_decap_8 FILLER_53_1579 ();
 sg13g2_decap_8 FILLER_53_1586 ();
 sg13g2_decap_8 FILLER_53_1593 ();
 sg13g2_decap_8 FILLER_53_1600 ();
 sg13g2_decap_8 FILLER_53_1607 ();
 sg13g2_decap_8 FILLER_53_1614 ();
 sg13g2_decap_8 FILLER_53_1621 ();
 sg13g2_decap_8 FILLER_53_1628 ();
 sg13g2_decap_8 FILLER_53_1635 ();
 sg13g2_decap_8 FILLER_53_1642 ();
 sg13g2_decap_8 FILLER_53_1649 ();
 sg13g2_decap_8 FILLER_53_1656 ();
 sg13g2_decap_8 FILLER_53_1663 ();
 sg13g2_decap_8 FILLER_53_1670 ();
 sg13g2_decap_8 FILLER_53_1677 ();
 sg13g2_decap_8 FILLER_53_1684 ();
 sg13g2_decap_8 FILLER_53_1691 ();
 sg13g2_decap_8 FILLER_53_1698 ();
 sg13g2_decap_8 FILLER_53_1705 ();
 sg13g2_decap_8 FILLER_53_1712 ();
 sg13g2_decap_8 FILLER_53_1719 ();
 sg13g2_decap_8 FILLER_53_1726 ();
 sg13g2_decap_8 FILLER_53_1733 ();
 sg13g2_decap_8 FILLER_53_1740 ();
 sg13g2_decap_8 FILLER_53_1747 ();
 sg13g2_decap_8 FILLER_53_1754 ();
 sg13g2_decap_8 FILLER_53_1761 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_decap_4 FILLER_54_222 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_8 FILLER_54_246 ();
 sg13g2_decap_8 FILLER_54_253 ();
 sg13g2_fill_2 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_262 ();
 sg13g2_decap_4 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_316 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_decap_8 FILLER_54_330 ();
 sg13g2_decap_8 FILLER_54_337 ();
 sg13g2_decap_8 FILLER_54_344 ();
 sg13g2_decap_8 FILLER_54_351 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_fill_2 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_8 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_441 ();
 sg13g2_decap_8 FILLER_54_456 ();
 sg13g2_decap_8 FILLER_54_463 ();
 sg13g2_decap_8 FILLER_54_470 ();
 sg13g2_decap_8 FILLER_54_477 ();
 sg13g2_decap_8 FILLER_54_484 ();
 sg13g2_decap_8 FILLER_54_491 ();
 sg13g2_decap_8 FILLER_54_498 ();
 sg13g2_decap_4 FILLER_54_505 ();
 sg13g2_fill_1 FILLER_54_509 ();
 sg13g2_decap_8 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_526 ();
 sg13g2_decap_8 FILLER_54_540 ();
 sg13g2_decap_4 FILLER_54_547 ();
 sg13g2_fill_1 FILLER_54_551 ();
 sg13g2_decap_8 FILLER_54_556 ();
 sg13g2_decap_8 FILLER_54_563 ();
 sg13g2_decap_8 FILLER_54_570 ();
 sg13g2_decap_8 FILLER_54_577 ();
 sg13g2_decap_8 FILLER_54_584 ();
 sg13g2_decap_8 FILLER_54_591 ();
 sg13g2_decap_8 FILLER_54_615 ();
 sg13g2_decap_8 FILLER_54_622 ();
 sg13g2_decap_8 FILLER_54_637 ();
 sg13g2_decap_8 FILLER_54_644 ();
 sg13g2_decap_8 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_decap_8 FILLER_54_672 ();
 sg13g2_decap_8 FILLER_54_679 ();
 sg13g2_fill_1 FILLER_54_686 ();
 sg13g2_decap_8 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_708 ();
 sg13g2_decap_8 FILLER_54_729 ();
 sg13g2_decap_8 FILLER_54_736 ();
 sg13g2_decap_8 FILLER_54_743 ();
 sg13g2_decap_8 FILLER_54_750 ();
 sg13g2_fill_1 FILLER_54_757 ();
 sg13g2_decap_8 FILLER_54_774 ();
 sg13g2_fill_1 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_fill_1 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_8 FILLER_54_856 ();
 sg13g2_decap_8 FILLER_54_863 ();
 sg13g2_decap_8 FILLER_54_870 ();
 sg13g2_decap_8 FILLER_54_877 ();
 sg13g2_decap_8 FILLER_54_884 ();
 sg13g2_decap_8 FILLER_54_891 ();
 sg13g2_fill_2 FILLER_54_898 ();
 sg13g2_decap_8 FILLER_54_905 ();
 sg13g2_decap_8 FILLER_54_912 ();
 sg13g2_decap_8 FILLER_54_919 ();
 sg13g2_decap_8 FILLER_54_926 ();
 sg13g2_decap_8 FILLER_54_933 ();
 sg13g2_decap_8 FILLER_54_940 ();
 sg13g2_fill_2 FILLER_54_947 ();
 sg13g2_fill_2 FILLER_54_952 ();
 sg13g2_fill_2 FILLER_54_963 ();
 sg13g2_decap_8 FILLER_54_970 ();
 sg13g2_decap_8 FILLER_54_977 ();
 sg13g2_decap_8 FILLER_54_984 ();
 sg13g2_fill_2 FILLER_54_991 ();
 sg13g2_decap_8 FILLER_54_1001 ();
 sg13g2_decap_8 FILLER_54_1008 ();
 sg13g2_decap_8 FILLER_54_1015 ();
 sg13g2_decap_8 FILLER_54_1022 ();
 sg13g2_decap_8 FILLER_54_1029 ();
 sg13g2_decap_8 FILLER_54_1036 ();
 sg13g2_fill_2 FILLER_54_1043 ();
 sg13g2_fill_1 FILLER_54_1045 ();
 sg13g2_decap_8 FILLER_54_1064 ();
 sg13g2_decap_4 FILLER_54_1071 ();
 sg13g2_decap_4 FILLER_54_1080 ();
 sg13g2_fill_2 FILLER_54_1084 ();
 sg13g2_decap_8 FILLER_54_1094 ();
 sg13g2_decap_8 FILLER_54_1101 ();
 sg13g2_decap_8 FILLER_54_1108 ();
 sg13g2_decap_8 FILLER_54_1115 ();
 sg13g2_decap_8 FILLER_54_1122 ();
 sg13g2_decap_8 FILLER_54_1137 ();
 sg13g2_fill_2 FILLER_54_1149 ();
 sg13g2_fill_1 FILLER_54_1151 ();
 sg13g2_decap_8 FILLER_54_1164 ();
 sg13g2_decap_8 FILLER_54_1171 ();
 sg13g2_decap_8 FILLER_54_1178 ();
 sg13g2_decap_8 FILLER_54_1211 ();
 sg13g2_decap_8 FILLER_54_1218 ();
 sg13g2_decap_4 FILLER_54_1225 ();
 sg13g2_fill_1 FILLER_54_1229 ();
 sg13g2_decap_8 FILLER_54_1238 ();
 sg13g2_fill_1 FILLER_54_1245 ();
 sg13g2_decap_8 FILLER_54_1250 ();
 sg13g2_decap_8 FILLER_54_1257 ();
 sg13g2_decap_8 FILLER_54_1264 ();
 sg13g2_decap_4 FILLER_54_1271 ();
 sg13g2_decap_4 FILLER_54_1279 ();
 sg13g2_fill_1 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1288 ();
 sg13g2_decap_8 FILLER_54_1295 ();
 sg13g2_decap_8 FILLER_54_1302 ();
 sg13g2_fill_2 FILLER_54_1330 ();
 sg13g2_fill_1 FILLER_54_1332 ();
 sg13g2_fill_1 FILLER_54_1345 ();
 sg13g2_decap_8 FILLER_54_1354 ();
 sg13g2_decap_8 FILLER_54_1361 ();
 sg13g2_decap_4 FILLER_54_1368 ();
 sg13g2_decap_8 FILLER_54_1398 ();
 sg13g2_decap_8 FILLER_54_1405 ();
 sg13g2_decap_8 FILLER_54_1412 ();
 sg13g2_decap_8 FILLER_54_1419 ();
 sg13g2_decap_8 FILLER_54_1426 ();
 sg13g2_fill_2 FILLER_54_1433 ();
 sg13g2_fill_1 FILLER_54_1435 ();
 sg13g2_decap_8 FILLER_54_1448 ();
 sg13g2_decap_8 FILLER_54_1455 ();
 sg13g2_fill_1 FILLER_54_1462 ();
 sg13g2_fill_2 FILLER_54_1475 ();
 sg13g2_decap_8 FILLER_54_1493 ();
 sg13g2_decap_8 FILLER_54_1500 ();
 sg13g2_fill_2 FILLER_54_1507 ();
 sg13g2_decap_8 FILLER_54_1517 ();
 sg13g2_decap_8 FILLER_54_1524 ();
 sg13g2_decap_8 FILLER_54_1531 ();
 sg13g2_decap_8 FILLER_54_1538 ();
 sg13g2_decap_8 FILLER_54_1545 ();
 sg13g2_fill_1 FILLER_54_1552 ();
 sg13g2_fill_1 FILLER_54_1562 ();
 sg13g2_decap_8 FILLER_54_1587 ();
 sg13g2_decap_8 FILLER_54_1594 ();
 sg13g2_decap_8 FILLER_54_1601 ();
 sg13g2_decap_8 FILLER_54_1608 ();
 sg13g2_decap_8 FILLER_54_1615 ();
 sg13g2_decap_8 FILLER_54_1622 ();
 sg13g2_decap_8 FILLER_54_1629 ();
 sg13g2_decap_8 FILLER_54_1636 ();
 sg13g2_decap_8 FILLER_54_1643 ();
 sg13g2_decap_8 FILLER_54_1650 ();
 sg13g2_decap_8 FILLER_54_1657 ();
 sg13g2_decap_8 FILLER_54_1664 ();
 sg13g2_decap_8 FILLER_54_1671 ();
 sg13g2_decap_8 FILLER_54_1678 ();
 sg13g2_decap_8 FILLER_54_1685 ();
 sg13g2_decap_8 FILLER_54_1692 ();
 sg13g2_decap_8 FILLER_54_1699 ();
 sg13g2_decap_8 FILLER_54_1706 ();
 sg13g2_decap_8 FILLER_54_1713 ();
 sg13g2_decap_8 FILLER_54_1720 ();
 sg13g2_decap_8 FILLER_54_1727 ();
 sg13g2_decap_8 FILLER_54_1734 ();
 sg13g2_decap_8 FILLER_54_1741 ();
 sg13g2_decap_8 FILLER_54_1748 ();
 sg13g2_decap_8 FILLER_54_1755 ();
 sg13g2_decap_4 FILLER_54_1762 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_220 ();
 sg13g2_decap_8 FILLER_55_227 ();
 sg13g2_decap_8 FILLER_55_234 ();
 sg13g2_decap_8 FILLER_55_241 ();
 sg13g2_decap_8 FILLER_55_248 ();
 sg13g2_fill_2 FILLER_55_255 ();
 sg13g2_fill_1 FILLER_55_257 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_decap_8 FILLER_55_282 ();
 sg13g2_decap_8 FILLER_55_289 ();
 sg13g2_decap_8 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_311 ();
 sg13g2_decap_8 FILLER_55_318 ();
 sg13g2_decap_8 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_332 ();
 sg13g2_decap_4 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_356 ();
 sg13g2_fill_1 FILLER_55_363 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_fill_1 FILLER_55_404 ();
 sg13g2_fill_2 FILLER_55_413 ();
 sg13g2_fill_1 FILLER_55_419 ();
 sg13g2_fill_1 FILLER_55_424 ();
 sg13g2_decap_8 FILLER_55_437 ();
 sg13g2_fill_1 FILLER_55_444 ();
 sg13g2_fill_2 FILLER_55_449 ();
 sg13g2_decap_8 FILLER_55_456 ();
 sg13g2_decap_8 FILLER_55_463 ();
 sg13g2_decap_8 FILLER_55_470 ();
 sg13g2_decap_8 FILLER_55_477 ();
 sg13g2_fill_2 FILLER_55_484 ();
 sg13g2_decap_8 FILLER_55_494 ();
 sg13g2_decap_8 FILLER_55_501 ();
 sg13g2_decap_8 FILLER_55_508 ();
 sg13g2_decap_8 FILLER_55_515 ();
 sg13g2_decap_4 FILLER_55_522 ();
 sg13g2_fill_2 FILLER_55_550 ();
 sg13g2_fill_1 FILLER_55_552 ();
 sg13g2_fill_2 FILLER_55_557 ();
 sg13g2_fill_2 FILLER_55_564 ();
 sg13g2_fill_2 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_574 ();
 sg13g2_decap_4 FILLER_55_581 ();
 sg13g2_decap_4 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_601 ();
 sg13g2_decap_8 FILLER_55_606 ();
 sg13g2_decap_8 FILLER_55_613 ();
 sg13g2_decap_8 FILLER_55_620 ();
 sg13g2_decap_8 FILLER_55_627 ();
 sg13g2_decap_8 FILLER_55_634 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_decap_8 FILLER_55_648 ();
 sg13g2_decap_8 FILLER_55_655 ();
 sg13g2_fill_2 FILLER_55_662 ();
 sg13g2_decap_8 FILLER_55_672 ();
 sg13g2_decap_4 FILLER_55_679 ();
 sg13g2_fill_1 FILLER_55_683 ();
 sg13g2_decap_8 FILLER_55_692 ();
 sg13g2_decap_8 FILLER_55_699 ();
 sg13g2_decap_8 FILLER_55_706 ();
 sg13g2_decap_8 FILLER_55_713 ();
 sg13g2_fill_1 FILLER_55_720 ();
 sg13g2_fill_2 FILLER_55_732 ();
 sg13g2_fill_1 FILLER_55_734 ();
 sg13g2_decap_8 FILLER_55_747 ();
 sg13g2_fill_2 FILLER_55_754 ();
 sg13g2_fill_1 FILLER_55_756 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_771 ();
 sg13g2_decap_8 FILLER_55_778 ();
 sg13g2_decap_8 FILLER_55_785 ();
 sg13g2_decap_8 FILLER_55_792 ();
 sg13g2_decap_8 FILLER_55_799 ();
 sg13g2_decap_8 FILLER_55_806 ();
 sg13g2_decap_8 FILLER_55_813 ();
 sg13g2_fill_2 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_834 ();
 sg13g2_decap_8 FILLER_55_841 ();
 sg13g2_decap_8 FILLER_55_848 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_55_862 ();
 sg13g2_decap_8 FILLER_55_869 ();
 sg13g2_decap_8 FILLER_55_876 ();
 sg13g2_decap_8 FILLER_55_883 ();
 sg13g2_decap_4 FILLER_55_890 ();
 sg13g2_decap_8 FILLER_55_912 ();
 sg13g2_decap_8 FILLER_55_925 ();
 sg13g2_decap_8 FILLER_55_932 ();
 sg13g2_decap_8 FILLER_55_939 ();
 sg13g2_decap_8 FILLER_55_946 ();
 sg13g2_decap_8 FILLER_55_974 ();
 sg13g2_decap_8 FILLER_55_981 ();
 sg13g2_decap_8 FILLER_55_1017 ();
 sg13g2_decap_8 FILLER_55_1024 ();
 sg13g2_decap_8 FILLER_55_1031 ();
 sg13g2_decap_8 FILLER_55_1038 ();
 sg13g2_fill_2 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1047 ();
 sg13g2_fill_1 FILLER_55_1069 ();
 sg13g2_decap_8 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1098 ();
 sg13g2_decap_8 FILLER_55_1105 ();
 sg13g2_fill_2 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1122 ();
 sg13g2_decap_8 FILLER_55_1129 ();
 sg13g2_fill_2 FILLER_55_1136 ();
 sg13g2_fill_1 FILLER_55_1138 ();
 sg13g2_decap_8 FILLER_55_1169 ();
 sg13g2_decap_8 FILLER_55_1176 ();
 sg13g2_decap_8 FILLER_55_1183 ();
 sg13g2_decap_8 FILLER_55_1190 ();
 sg13g2_decap_8 FILLER_55_1197 ();
 sg13g2_decap_8 FILLER_55_1204 ();
 sg13g2_decap_8 FILLER_55_1211 ();
 sg13g2_decap_8 FILLER_55_1218 ();
 sg13g2_decap_4 FILLER_55_1225 ();
 sg13g2_fill_1 FILLER_55_1229 ();
 sg13g2_decap_8 FILLER_55_1233 ();
 sg13g2_decap_8 FILLER_55_1240 ();
 sg13g2_fill_1 FILLER_55_1247 ();
 sg13g2_fill_2 FILLER_55_1252 ();
 sg13g2_fill_1 FILLER_55_1254 ();
 sg13g2_decap_4 FILLER_55_1263 ();
 sg13g2_fill_2 FILLER_55_1267 ();
 sg13g2_decap_8 FILLER_55_1290 ();
 sg13g2_decap_4 FILLER_55_1297 ();
 sg13g2_decap_4 FILLER_55_1312 ();
 sg13g2_fill_2 FILLER_55_1316 ();
 sg13g2_decap_8 FILLER_55_1322 ();
 sg13g2_decap_8 FILLER_55_1333 ();
 sg13g2_decap_8 FILLER_55_1340 ();
 sg13g2_decap_8 FILLER_55_1347 ();
 sg13g2_decap_8 FILLER_55_1354 ();
 sg13g2_decap_8 FILLER_55_1361 ();
 sg13g2_decap_8 FILLER_55_1368 ();
 sg13g2_decap_8 FILLER_55_1375 ();
 sg13g2_decap_4 FILLER_55_1382 ();
 sg13g2_decap_8 FILLER_55_1394 ();
 sg13g2_fill_2 FILLER_55_1401 ();
 sg13g2_decap_8 FILLER_55_1412 ();
 sg13g2_decap_8 FILLER_55_1419 ();
 sg13g2_decap_4 FILLER_55_1426 ();
 sg13g2_fill_1 FILLER_55_1430 ();
 sg13g2_fill_2 FILLER_55_1437 ();
 sg13g2_decap_8 FILLER_55_1447 ();
 sg13g2_decap_8 FILLER_55_1454 ();
 sg13g2_decap_8 FILLER_55_1461 ();
 sg13g2_decap_8 FILLER_55_1468 ();
 sg13g2_decap_8 FILLER_55_1475 ();
 sg13g2_fill_2 FILLER_55_1482 ();
 sg13g2_fill_1 FILLER_55_1484 ();
 sg13g2_fill_2 FILLER_55_1490 ();
 sg13g2_fill_1 FILLER_55_1492 ();
 sg13g2_decap_4 FILLER_55_1501 ();
 sg13g2_fill_2 FILLER_55_1513 ();
 sg13g2_fill_1 FILLER_55_1515 ();
 sg13g2_decap_8 FILLER_55_1524 ();
 sg13g2_decap_8 FILLER_55_1531 ();
 sg13g2_decap_8 FILLER_55_1538 ();
 sg13g2_decap_8 FILLER_55_1545 ();
 sg13g2_decap_8 FILLER_55_1552 ();
 sg13g2_fill_1 FILLER_55_1559 ();
 sg13g2_fill_2 FILLER_55_1564 ();
 sg13g2_fill_1 FILLER_55_1566 ();
 sg13g2_decap_8 FILLER_55_1580 ();
 sg13g2_decap_8 FILLER_55_1587 ();
 sg13g2_decap_8 FILLER_55_1594 ();
 sg13g2_decap_8 FILLER_55_1601 ();
 sg13g2_decap_8 FILLER_55_1608 ();
 sg13g2_decap_8 FILLER_55_1615 ();
 sg13g2_decap_8 FILLER_55_1622 ();
 sg13g2_decap_8 FILLER_55_1629 ();
 sg13g2_decap_8 FILLER_55_1636 ();
 sg13g2_decap_8 FILLER_55_1643 ();
 sg13g2_decap_8 FILLER_55_1650 ();
 sg13g2_decap_8 FILLER_55_1657 ();
 sg13g2_decap_8 FILLER_55_1664 ();
 sg13g2_decap_8 FILLER_55_1671 ();
 sg13g2_decap_8 FILLER_55_1678 ();
 sg13g2_decap_8 FILLER_55_1685 ();
 sg13g2_decap_8 FILLER_55_1692 ();
 sg13g2_decap_8 FILLER_55_1699 ();
 sg13g2_decap_8 FILLER_55_1706 ();
 sg13g2_decap_8 FILLER_55_1713 ();
 sg13g2_decap_8 FILLER_55_1720 ();
 sg13g2_decap_8 FILLER_55_1727 ();
 sg13g2_decap_8 FILLER_55_1734 ();
 sg13g2_decap_8 FILLER_55_1741 ();
 sg13g2_decap_8 FILLER_55_1748 ();
 sg13g2_decap_8 FILLER_55_1755 ();
 sg13g2_decap_4 FILLER_55_1762 ();
 sg13g2_fill_2 FILLER_55_1766 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_4 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_205 ();
 sg13g2_decap_8 FILLER_56_212 ();
 sg13g2_decap_8 FILLER_56_219 ();
 sg13g2_decap_8 FILLER_56_226 ();
 sg13g2_decap_4 FILLER_56_233 ();
 sg13g2_fill_2 FILLER_56_237 ();
 sg13g2_fill_2 FILLER_56_244 ();
 sg13g2_decap_8 FILLER_56_282 ();
 sg13g2_decap_8 FILLER_56_289 ();
 sg13g2_decap_8 FILLER_56_296 ();
 sg13g2_decap_8 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_310 ();
 sg13g2_decap_8 FILLER_56_317 ();
 sg13g2_decap_8 FILLER_56_324 ();
 sg13g2_fill_2 FILLER_56_331 ();
 sg13g2_decap_8 FILLER_56_355 ();
 sg13g2_decap_8 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_56_409 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_8 FILLER_56_430 ();
 sg13g2_decap_8 FILLER_56_437 ();
 sg13g2_decap_8 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_451 ();
 sg13g2_fill_2 FILLER_56_458 ();
 sg13g2_decap_4 FILLER_56_468 ();
 sg13g2_fill_2 FILLER_56_472 ();
 sg13g2_decap_8 FILLER_56_495 ();
 sg13g2_decap_8 FILLER_56_502 ();
 sg13g2_decap_4 FILLER_56_509 ();
 sg13g2_fill_1 FILLER_56_513 ();
 sg13g2_decap_4 FILLER_56_520 ();
 sg13g2_decap_8 FILLER_56_536 ();
 sg13g2_decap_8 FILLER_56_543 ();
 sg13g2_decap_8 FILLER_56_550 ();
 sg13g2_decap_8 FILLER_56_557 ();
 sg13g2_decap_8 FILLER_56_564 ();
 sg13g2_decap_4 FILLER_56_571 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_decap_8 FILLER_56_609 ();
 sg13g2_fill_2 FILLER_56_616 ();
 sg13g2_decap_8 FILLER_56_626 ();
 sg13g2_decap_8 FILLER_56_633 ();
 sg13g2_decap_8 FILLER_56_640 ();
 sg13g2_decap_8 FILLER_56_647 ();
 sg13g2_decap_8 FILLER_56_654 ();
 sg13g2_decap_8 FILLER_56_661 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_decap_8 FILLER_56_675 ();
 sg13g2_decap_8 FILLER_56_682 ();
 sg13g2_decap_8 FILLER_56_689 ();
 sg13g2_decap_8 FILLER_56_696 ();
 sg13g2_fill_1 FILLER_56_703 ();
 sg13g2_decap_8 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_4 FILLER_56_726 ();
 sg13g2_fill_2 FILLER_56_730 ();
 sg13g2_decap_8 FILLER_56_736 ();
 sg13g2_decap_8 FILLER_56_743 ();
 sg13g2_fill_2 FILLER_56_750 ();
 sg13g2_fill_1 FILLER_56_752 ();
 sg13g2_decap_8 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_decap_8 FILLER_56_774 ();
 sg13g2_decap_8 FILLER_56_781 ();
 sg13g2_decap_8 FILLER_56_788 ();
 sg13g2_decap_8 FILLER_56_795 ();
 sg13g2_decap_8 FILLER_56_802 ();
 sg13g2_fill_2 FILLER_56_809 ();
 sg13g2_fill_1 FILLER_56_811 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_8 FILLER_56_856 ();
 sg13g2_decap_8 FILLER_56_863 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_decap_8 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_56_884 ();
 sg13g2_fill_1 FILLER_56_891 ();
 sg13g2_decap_8 FILLER_56_926 ();
 sg13g2_decap_8 FILLER_56_933 ();
 sg13g2_decap_8 FILLER_56_940 ();
 sg13g2_decap_8 FILLER_56_947 ();
 sg13g2_decap_8 FILLER_56_954 ();
 sg13g2_decap_8 FILLER_56_966 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_decap_8 FILLER_56_980 ();
 sg13g2_decap_4 FILLER_56_987 ();
 sg13g2_decap_4 FILLER_56_995 ();
 sg13g2_fill_2 FILLER_56_999 ();
 sg13g2_decap_8 FILLER_56_1020 ();
 sg13g2_decap_8 FILLER_56_1027 ();
 sg13g2_decap_8 FILLER_56_1034 ();
 sg13g2_decap_8 FILLER_56_1041 ();
 sg13g2_decap_4 FILLER_56_1048 ();
 sg13g2_fill_2 FILLER_56_1052 ();
 sg13g2_decap_8 FILLER_56_1065 ();
 sg13g2_decap_8 FILLER_56_1072 ();
 sg13g2_decap_8 FILLER_56_1079 ();
 sg13g2_decap_8 FILLER_56_1086 ();
 sg13g2_decap_8 FILLER_56_1093 ();
 sg13g2_decap_8 FILLER_56_1100 ();
 sg13g2_decap_8 FILLER_56_1107 ();
 sg13g2_decap_8 FILLER_56_1114 ();
 sg13g2_decap_8 FILLER_56_1121 ();
 sg13g2_decap_8 FILLER_56_1128 ();
 sg13g2_fill_2 FILLER_56_1135 ();
 sg13g2_decap_8 FILLER_56_1145 ();
 sg13g2_decap_8 FILLER_56_1152 ();
 sg13g2_decap_8 FILLER_56_1159 ();
 sg13g2_decap_8 FILLER_56_1166 ();
 sg13g2_decap_8 FILLER_56_1173 ();
 sg13g2_decap_8 FILLER_56_1180 ();
 sg13g2_decap_8 FILLER_56_1187 ();
 sg13g2_decap_8 FILLER_56_1194 ();
 sg13g2_decap_8 FILLER_56_1201 ();
 sg13g2_fill_2 FILLER_56_1208 ();
 sg13g2_fill_1 FILLER_56_1218 ();
 sg13g2_decap_8 FILLER_56_1227 ();
 sg13g2_decap_4 FILLER_56_1234 ();
 sg13g2_fill_2 FILLER_56_1238 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1267 ();
 sg13g2_decap_8 FILLER_56_1274 ();
 sg13g2_decap_8 FILLER_56_1281 ();
 sg13g2_fill_1 FILLER_56_1288 ();
 sg13g2_fill_2 FILLER_56_1293 ();
 sg13g2_decap_4 FILLER_56_1303 ();
 sg13g2_fill_1 FILLER_56_1307 ();
 sg13g2_decap_8 FILLER_56_1319 ();
 sg13g2_decap_8 FILLER_56_1326 ();
 sg13g2_decap_8 FILLER_56_1333 ();
 sg13g2_decap_8 FILLER_56_1340 ();
 sg13g2_decap_8 FILLER_56_1347 ();
 sg13g2_fill_2 FILLER_56_1354 ();
 sg13g2_fill_2 FILLER_56_1360 ();
 sg13g2_fill_2 FILLER_56_1375 ();
 sg13g2_decap_8 FILLER_56_1389 ();
 sg13g2_decap_8 FILLER_56_1396 ();
 sg13g2_decap_8 FILLER_56_1403 ();
 sg13g2_decap_8 FILLER_56_1410 ();
 sg13g2_decap_4 FILLER_56_1417 ();
 sg13g2_fill_2 FILLER_56_1421 ();
 sg13g2_fill_1 FILLER_56_1435 ();
 sg13g2_decap_8 FILLER_56_1449 ();
 sg13g2_decap_8 FILLER_56_1456 ();
 sg13g2_decap_8 FILLER_56_1463 ();
 sg13g2_decap_8 FILLER_56_1470 ();
 sg13g2_decap_4 FILLER_56_1477 ();
 sg13g2_decap_8 FILLER_56_1497 ();
 sg13g2_decap_8 FILLER_56_1504 ();
 sg13g2_decap_8 FILLER_56_1511 ();
 sg13g2_decap_8 FILLER_56_1518 ();
 sg13g2_decap_8 FILLER_56_1525 ();
 sg13g2_decap_8 FILLER_56_1532 ();
 sg13g2_decap_8 FILLER_56_1539 ();
 sg13g2_decap_8 FILLER_56_1546 ();
 sg13g2_fill_2 FILLER_56_1553 ();
 sg13g2_fill_1 FILLER_56_1555 ();
 sg13g2_decap_4 FILLER_56_1564 ();
 sg13g2_fill_2 FILLER_56_1568 ();
 sg13g2_decap_8 FILLER_56_1579 ();
 sg13g2_decap_8 FILLER_56_1586 ();
 sg13g2_decap_8 FILLER_56_1593 ();
 sg13g2_decap_8 FILLER_56_1600 ();
 sg13g2_decap_8 FILLER_56_1607 ();
 sg13g2_decap_8 FILLER_56_1614 ();
 sg13g2_decap_8 FILLER_56_1621 ();
 sg13g2_decap_8 FILLER_56_1628 ();
 sg13g2_decap_8 FILLER_56_1635 ();
 sg13g2_decap_8 FILLER_56_1642 ();
 sg13g2_decap_8 FILLER_56_1649 ();
 sg13g2_decap_8 FILLER_56_1656 ();
 sg13g2_decap_8 FILLER_56_1663 ();
 sg13g2_decap_8 FILLER_56_1670 ();
 sg13g2_decap_8 FILLER_56_1677 ();
 sg13g2_decap_8 FILLER_56_1684 ();
 sg13g2_decap_8 FILLER_56_1691 ();
 sg13g2_decap_8 FILLER_56_1698 ();
 sg13g2_decap_8 FILLER_56_1705 ();
 sg13g2_decap_8 FILLER_56_1712 ();
 sg13g2_decap_8 FILLER_56_1719 ();
 sg13g2_decap_8 FILLER_56_1726 ();
 sg13g2_decap_8 FILLER_56_1733 ();
 sg13g2_decap_8 FILLER_56_1740 ();
 sg13g2_decap_8 FILLER_56_1747 ();
 sg13g2_decap_8 FILLER_56_1754 ();
 sg13g2_decap_8 FILLER_56_1761 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_fill_1 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_340 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_4 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_decap_4 FILLER_57_393 ();
 sg13g2_fill_2 FILLER_57_397 ();
 sg13g2_decap_8 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_414 ();
 sg13g2_fill_2 FILLER_57_421 ();
 sg13g2_fill_1 FILLER_57_423 ();
 sg13g2_decap_4 FILLER_57_436 ();
 sg13g2_decap_4 FILLER_57_448 ();
 sg13g2_fill_1 FILLER_57_452 ();
 sg13g2_decap_8 FILLER_57_474 ();
 sg13g2_decap_8 FILLER_57_481 ();
 sg13g2_decap_8 FILLER_57_488 ();
 sg13g2_decap_8 FILLER_57_495 ();
 sg13g2_decap_8 FILLER_57_502 ();
 sg13g2_decap_4 FILLER_57_509 ();
 sg13g2_fill_1 FILLER_57_513 ();
 sg13g2_decap_8 FILLER_57_546 ();
 sg13g2_decap_8 FILLER_57_553 ();
 sg13g2_decap_8 FILLER_57_560 ();
 sg13g2_fill_2 FILLER_57_567 ();
 sg13g2_fill_1 FILLER_57_569 ();
 sg13g2_decap_8 FILLER_57_578 ();
 sg13g2_fill_2 FILLER_57_585 ();
 sg13g2_decap_8 FILLER_57_592 ();
 sg13g2_decap_8 FILLER_57_599 ();
 sg13g2_decap_8 FILLER_57_606 ();
 sg13g2_fill_1 FILLER_57_613 ();
 sg13g2_decap_8 FILLER_57_635 ();
 sg13g2_decap_8 FILLER_57_642 ();
 sg13g2_decap_8 FILLER_57_649 ();
 sg13g2_decap_8 FILLER_57_656 ();
 sg13g2_decap_8 FILLER_57_663 ();
 sg13g2_decap_8 FILLER_57_670 ();
 sg13g2_decap_8 FILLER_57_677 ();
 sg13g2_decap_8 FILLER_57_684 ();
 sg13g2_decap_8 FILLER_57_691 ();
 sg13g2_decap_8 FILLER_57_714 ();
 sg13g2_decap_8 FILLER_57_721 ();
 sg13g2_decap_8 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_735 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_749 ();
 sg13g2_decap_8 FILLER_57_756 ();
 sg13g2_decap_8 FILLER_57_763 ();
 sg13g2_decap_8 FILLER_57_770 ();
 sg13g2_decap_8 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_784 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_fill_2 FILLER_57_798 ();
 sg13g2_fill_1 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_809 ();
 sg13g2_fill_1 FILLER_57_816 ();
 sg13g2_decap_4 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_848 ();
 sg13g2_decap_8 FILLER_57_855 ();
 sg13g2_decap_8 FILLER_57_862 ();
 sg13g2_decap_4 FILLER_57_869 ();
 sg13g2_fill_1 FILLER_57_873 ();
 sg13g2_decap_4 FILLER_57_880 ();
 sg13g2_fill_1 FILLER_57_884 ();
 sg13g2_decap_4 FILLER_57_893 ();
 sg13g2_fill_1 FILLER_57_897 ();
 sg13g2_fill_1 FILLER_57_905 ();
 sg13g2_decap_8 FILLER_57_914 ();
 sg13g2_decap_4 FILLER_57_921 ();
 sg13g2_fill_2 FILLER_57_925 ();
 sg13g2_decap_8 FILLER_57_930 ();
 sg13g2_decap_8 FILLER_57_937 ();
 sg13g2_fill_1 FILLER_57_944 ();
 sg13g2_decap_8 FILLER_57_953 ();
 sg13g2_decap_8 FILLER_57_960 ();
 sg13g2_decap_8 FILLER_57_967 ();
 sg13g2_decap_8 FILLER_57_974 ();
 sg13g2_decap_8 FILLER_57_981 ();
 sg13g2_decap_8 FILLER_57_988 ();
 sg13g2_decap_8 FILLER_57_995 ();
 sg13g2_decap_8 FILLER_57_1002 ();
 sg13g2_fill_2 FILLER_57_1009 ();
 sg13g2_decap_8 FILLER_57_1031 ();
 sg13g2_decap_8 FILLER_57_1038 ();
 sg13g2_decap_8 FILLER_57_1045 ();
 sg13g2_decap_8 FILLER_57_1052 ();
 sg13g2_decap_8 FILLER_57_1059 ();
 sg13g2_decap_8 FILLER_57_1066 ();
 sg13g2_decap_8 FILLER_57_1073 ();
 sg13g2_decap_4 FILLER_57_1080 ();
 sg13g2_fill_2 FILLER_57_1084 ();
 sg13g2_decap_8 FILLER_57_1094 ();
 sg13g2_fill_1 FILLER_57_1101 ();
 sg13g2_decap_8 FILLER_57_1110 ();
 sg13g2_decap_8 FILLER_57_1117 ();
 sg13g2_decap_8 FILLER_57_1124 ();
 sg13g2_decap_4 FILLER_57_1131 ();
 sg13g2_fill_2 FILLER_57_1143 ();
 sg13g2_decap_8 FILLER_57_1155 ();
 sg13g2_decap_8 FILLER_57_1162 ();
 sg13g2_decap_8 FILLER_57_1169 ();
 sg13g2_decap_8 FILLER_57_1176 ();
 sg13g2_decap_8 FILLER_57_1183 ();
 sg13g2_decap_8 FILLER_57_1190 ();
 sg13g2_decap_8 FILLER_57_1197 ();
 sg13g2_fill_1 FILLER_57_1218 ();
 sg13g2_decap_8 FILLER_57_1227 ();
 sg13g2_decap_8 FILLER_57_1234 ();
 sg13g2_decap_8 FILLER_57_1241 ();
 sg13g2_decap_8 FILLER_57_1248 ();
 sg13g2_decap_8 FILLER_57_1255 ();
 sg13g2_decap_8 FILLER_57_1262 ();
 sg13g2_decap_4 FILLER_57_1269 ();
 sg13g2_fill_2 FILLER_57_1273 ();
 sg13g2_decap_8 FILLER_57_1283 ();
 sg13g2_fill_1 FILLER_57_1290 ();
 sg13g2_decap_8 FILLER_57_1296 ();
 sg13g2_decap_4 FILLER_57_1303 ();
 sg13g2_fill_1 FILLER_57_1307 ();
 sg13g2_decap_8 FILLER_57_1316 ();
 sg13g2_decap_8 FILLER_57_1323 ();
 sg13g2_decap_8 FILLER_57_1330 ();
 sg13g2_decap_8 FILLER_57_1337 ();
 sg13g2_fill_1 FILLER_57_1344 ();
 sg13g2_decap_8 FILLER_57_1371 ();
 sg13g2_decap_8 FILLER_57_1378 ();
 sg13g2_decap_8 FILLER_57_1385 ();
 sg13g2_decap_8 FILLER_57_1392 ();
 sg13g2_decap_8 FILLER_57_1399 ();
 sg13g2_decap_8 FILLER_57_1406 ();
 sg13g2_decap_8 FILLER_57_1413 ();
 sg13g2_decap_8 FILLER_57_1420 ();
 sg13g2_decap_8 FILLER_57_1427 ();
 sg13g2_fill_1 FILLER_57_1434 ();
 sg13g2_decap_8 FILLER_57_1439 ();
 sg13g2_decap_4 FILLER_57_1446 ();
 sg13g2_fill_2 FILLER_57_1450 ();
 sg13g2_decap_8 FILLER_57_1460 ();
 sg13g2_decap_8 FILLER_57_1467 ();
 sg13g2_decap_8 FILLER_57_1474 ();
 sg13g2_decap_8 FILLER_57_1481 ();
 sg13g2_decap_8 FILLER_57_1488 ();
 sg13g2_decap_8 FILLER_57_1495 ();
 sg13g2_decap_8 FILLER_57_1502 ();
 sg13g2_decap_8 FILLER_57_1509 ();
 sg13g2_decap_8 FILLER_57_1516 ();
 sg13g2_decap_4 FILLER_57_1523 ();
 sg13g2_fill_2 FILLER_57_1527 ();
 sg13g2_decap_8 FILLER_57_1545 ();
 sg13g2_decap_8 FILLER_57_1552 ();
 sg13g2_decap_8 FILLER_57_1559 ();
 sg13g2_fill_1 FILLER_57_1566 ();
 sg13g2_decap_8 FILLER_57_1571 ();
 sg13g2_decap_8 FILLER_57_1578 ();
 sg13g2_decap_8 FILLER_57_1585 ();
 sg13g2_decap_8 FILLER_57_1592 ();
 sg13g2_decap_8 FILLER_57_1599 ();
 sg13g2_decap_8 FILLER_57_1606 ();
 sg13g2_decap_8 FILLER_57_1613 ();
 sg13g2_decap_8 FILLER_57_1620 ();
 sg13g2_decap_8 FILLER_57_1627 ();
 sg13g2_decap_8 FILLER_57_1634 ();
 sg13g2_decap_8 FILLER_57_1641 ();
 sg13g2_decap_8 FILLER_57_1648 ();
 sg13g2_decap_8 FILLER_57_1655 ();
 sg13g2_decap_8 FILLER_57_1662 ();
 sg13g2_decap_8 FILLER_57_1669 ();
 sg13g2_decap_8 FILLER_57_1676 ();
 sg13g2_decap_8 FILLER_57_1683 ();
 sg13g2_decap_8 FILLER_57_1690 ();
 sg13g2_decap_8 FILLER_57_1697 ();
 sg13g2_decap_8 FILLER_57_1704 ();
 sg13g2_decap_8 FILLER_57_1711 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_8 FILLER_57_1725 ();
 sg13g2_decap_8 FILLER_57_1732 ();
 sg13g2_decap_8 FILLER_57_1739 ();
 sg13g2_decap_8 FILLER_57_1746 ();
 sg13g2_decap_8 FILLER_57_1753 ();
 sg13g2_decap_8 FILLER_57_1760 ();
 sg13g2_fill_1 FILLER_57_1767 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_180 ();
 sg13g2_decap_8 FILLER_58_214 ();
 sg13g2_decap_8 FILLER_58_221 ();
 sg13g2_decap_8 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_239 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_fill_1 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_291 ();
 sg13g2_decap_8 FILLER_58_298 ();
 sg13g2_decap_8 FILLER_58_305 ();
 sg13g2_decap_8 FILLER_58_312 ();
 sg13g2_decap_8 FILLER_58_319 ();
 sg13g2_decap_8 FILLER_58_347 ();
 sg13g2_decap_8 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_361 ();
 sg13g2_decap_8 FILLER_58_368 ();
 sg13g2_decap_8 FILLER_58_375 ();
 sg13g2_decap_8 FILLER_58_382 ();
 sg13g2_decap_4 FILLER_58_389 ();
 sg13g2_fill_2 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_405 ();
 sg13g2_decap_8 FILLER_58_412 ();
 sg13g2_decap_4 FILLER_58_419 ();
 sg13g2_fill_1 FILLER_58_423 ();
 sg13g2_decap_8 FILLER_58_445 ();
 sg13g2_decap_8 FILLER_58_452 ();
 sg13g2_decap_8 FILLER_58_459 ();
 sg13g2_decap_8 FILLER_58_466 ();
 sg13g2_decap_8 FILLER_58_473 ();
 sg13g2_decap_8 FILLER_58_480 ();
 sg13g2_decap_8 FILLER_58_487 ();
 sg13g2_decap_8 FILLER_58_494 ();
 sg13g2_decap_8 FILLER_58_501 ();
 sg13g2_decap_8 FILLER_58_516 ();
 sg13g2_decap_4 FILLER_58_523 ();
 sg13g2_fill_2 FILLER_58_527 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_decap_4 FILLER_58_553 ();
 sg13g2_fill_2 FILLER_58_557 ();
 sg13g2_decap_8 FILLER_58_571 ();
 sg13g2_decap_4 FILLER_58_578 ();
 sg13g2_fill_2 FILLER_58_582 ();
 sg13g2_decap_8 FILLER_58_592 ();
 sg13g2_decap_8 FILLER_58_599 ();
 sg13g2_decap_8 FILLER_58_606 ();
 sg13g2_decap_8 FILLER_58_613 ();
 sg13g2_decap_4 FILLER_58_620 ();
 sg13g2_fill_2 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_631 ();
 sg13g2_decap_8 FILLER_58_640 ();
 sg13g2_decap_8 FILLER_58_647 ();
 sg13g2_decap_8 FILLER_58_654 ();
 sg13g2_decap_8 FILLER_58_661 ();
 sg13g2_decap_4 FILLER_58_668 ();
 sg13g2_fill_1 FILLER_58_672 ();
 sg13g2_fill_2 FILLER_58_686 ();
 sg13g2_fill_1 FILLER_58_688 ();
 sg13g2_fill_2 FILLER_58_705 ();
 sg13g2_decap_8 FILLER_58_711 ();
 sg13g2_decap_8 FILLER_58_718 ();
 sg13g2_fill_2 FILLER_58_725 ();
 sg13g2_fill_1 FILLER_58_727 ();
 sg13g2_decap_8 FILLER_58_750 ();
 sg13g2_decap_8 FILLER_58_757 ();
 sg13g2_decap_8 FILLER_58_764 ();
 sg13g2_decap_4 FILLER_58_771 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_decap_8 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_decap_8 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_847 ();
 sg13g2_decap_8 FILLER_58_854 ();
 sg13g2_decap_8 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_58_868 ();
 sg13g2_fill_2 FILLER_58_883 ();
 sg13g2_fill_1 FILLER_58_885 ();
 sg13g2_decap_8 FILLER_58_902 ();
 sg13g2_decap_8 FILLER_58_909 ();
 sg13g2_decap_8 FILLER_58_916 ();
 sg13g2_decap_8 FILLER_58_923 ();
 sg13g2_decap_8 FILLER_58_930 ();
 sg13g2_fill_2 FILLER_58_937 ();
 sg13g2_decap_8 FILLER_58_961 ();
 sg13g2_decap_8 FILLER_58_968 ();
 sg13g2_decap_8 FILLER_58_975 ();
 sg13g2_decap_4 FILLER_58_982 ();
 sg13g2_decap_8 FILLER_58_1003 ();
 sg13g2_decap_8 FILLER_58_1010 ();
 sg13g2_fill_1 FILLER_58_1017 ();
 sg13g2_decap_8 FILLER_58_1022 ();
 sg13g2_fill_1 FILLER_58_1029 ();
 sg13g2_decap_8 FILLER_58_1038 ();
 sg13g2_decap_8 FILLER_58_1045 ();
 sg13g2_decap_8 FILLER_58_1052 ();
 sg13g2_decap_8 FILLER_58_1059 ();
 sg13g2_decap_8 FILLER_58_1066 ();
 sg13g2_decap_8 FILLER_58_1073 ();
 sg13g2_fill_2 FILLER_58_1080 ();
 sg13g2_fill_1 FILLER_58_1082 ();
 sg13g2_decap_4 FILLER_58_1086 ();
 sg13g2_decap_8 FILLER_58_1108 ();
 sg13g2_decap_4 FILLER_58_1115 ();
 sg13g2_decap_8 FILLER_58_1124 ();
 sg13g2_decap_4 FILLER_58_1131 ();
 sg13g2_decap_8 FILLER_58_1159 ();
 sg13g2_decap_8 FILLER_58_1176 ();
 sg13g2_decap_8 FILLER_58_1183 ();
 sg13g2_decap_8 FILLER_58_1190 ();
 sg13g2_decap_4 FILLER_58_1197 ();
 sg13g2_fill_1 FILLER_58_1201 ();
 sg13g2_decap_8 FILLER_58_1223 ();
 sg13g2_decap_4 FILLER_58_1230 ();
 sg13g2_decap_8 FILLER_58_1255 ();
 sg13g2_decap_8 FILLER_58_1262 ();
 sg13g2_fill_1 FILLER_58_1269 ();
 sg13g2_decap_8 FILLER_58_1292 ();
 sg13g2_decap_8 FILLER_58_1299 ();
 sg13g2_decap_8 FILLER_58_1306 ();
 sg13g2_decap_8 FILLER_58_1313 ();
 sg13g2_fill_2 FILLER_58_1320 ();
 sg13g2_decap_8 FILLER_58_1326 ();
 sg13g2_decap_8 FILLER_58_1333 ();
 sg13g2_decap_8 FILLER_58_1340 ();
 sg13g2_fill_1 FILLER_58_1347 ();
 sg13g2_decap_8 FILLER_58_1356 ();
 sg13g2_decap_8 FILLER_58_1363 ();
 sg13g2_decap_8 FILLER_58_1370 ();
 sg13g2_decap_8 FILLER_58_1377 ();
 sg13g2_fill_2 FILLER_58_1384 ();
 sg13g2_fill_1 FILLER_58_1386 ();
 sg13g2_fill_2 FILLER_58_1392 ();
 sg13g2_decap_8 FILLER_58_1402 ();
 sg13g2_decap_8 FILLER_58_1409 ();
 sg13g2_decap_8 FILLER_58_1416 ();
 sg13g2_decap_8 FILLER_58_1423 ();
 sg13g2_fill_2 FILLER_58_1430 ();
 sg13g2_decap_8 FILLER_58_1453 ();
 sg13g2_decap_8 FILLER_58_1460 ();
 sg13g2_decap_8 FILLER_58_1467 ();
 sg13g2_decap_8 FILLER_58_1474 ();
 sg13g2_decap_8 FILLER_58_1481 ();
 sg13g2_fill_2 FILLER_58_1488 ();
 sg13g2_fill_1 FILLER_58_1490 ();
 sg13g2_decap_8 FILLER_58_1499 ();
 sg13g2_decap_8 FILLER_58_1506 ();
 sg13g2_decap_8 FILLER_58_1513 ();
 sg13g2_fill_2 FILLER_58_1520 ();
 sg13g2_decap_8 FILLER_58_1546 ();
 sg13g2_decap_8 FILLER_58_1553 ();
 sg13g2_decap_4 FILLER_58_1560 ();
 sg13g2_fill_1 FILLER_58_1564 ();
 sg13g2_fill_2 FILLER_58_1573 ();
 sg13g2_decap_8 FILLER_58_1591 ();
 sg13g2_decap_8 FILLER_58_1598 ();
 sg13g2_decap_8 FILLER_58_1605 ();
 sg13g2_decap_8 FILLER_58_1612 ();
 sg13g2_decap_8 FILLER_58_1619 ();
 sg13g2_decap_8 FILLER_58_1626 ();
 sg13g2_decap_8 FILLER_58_1633 ();
 sg13g2_decap_8 FILLER_58_1640 ();
 sg13g2_decap_8 FILLER_58_1647 ();
 sg13g2_decap_8 FILLER_58_1654 ();
 sg13g2_decap_8 FILLER_58_1661 ();
 sg13g2_decap_8 FILLER_58_1668 ();
 sg13g2_decap_8 FILLER_58_1675 ();
 sg13g2_decap_8 FILLER_58_1682 ();
 sg13g2_decap_8 FILLER_58_1689 ();
 sg13g2_decap_8 FILLER_58_1696 ();
 sg13g2_decap_8 FILLER_58_1703 ();
 sg13g2_decap_8 FILLER_58_1710 ();
 sg13g2_decap_8 FILLER_58_1717 ();
 sg13g2_decap_8 FILLER_58_1724 ();
 sg13g2_decap_8 FILLER_58_1731 ();
 sg13g2_decap_8 FILLER_58_1738 ();
 sg13g2_decap_8 FILLER_58_1745 ();
 sg13g2_decap_8 FILLER_58_1752 ();
 sg13g2_decap_8 FILLER_58_1759 ();
 sg13g2_fill_2 FILLER_58_1766 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_fill_2 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_decap_8 FILLER_59_134 ();
 sg13g2_decap_8 FILLER_59_171 ();
 sg13g2_decap_4 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_182 ();
 sg13g2_decap_4 FILLER_59_187 ();
 sg13g2_fill_2 FILLER_59_191 ();
 sg13g2_decap_8 FILLER_59_219 ();
 sg13g2_decap_8 FILLER_59_239 ();
 sg13g2_decap_8 FILLER_59_246 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_4 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_decap_8 FILLER_59_288 ();
 sg13g2_decap_8 FILLER_59_295 ();
 sg13g2_decap_8 FILLER_59_302 ();
 sg13g2_decap_8 FILLER_59_309 ();
 sg13g2_decap_4 FILLER_59_316 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_decap_4 FILLER_59_340 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_4 FILLER_59_388 ();
 sg13g2_fill_2 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_409 ();
 sg13g2_decap_8 FILLER_59_416 ();
 sg13g2_decap_8 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_59_430 ();
 sg13g2_decap_8 FILLER_59_437 ();
 sg13g2_decap_8 FILLER_59_444 ();
 sg13g2_decap_8 FILLER_59_451 ();
 sg13g2_decap_8 FILLER_59_458 ();
 sg13g2_decap_8 FILLER_59_465 ();
 sg13g2_decap_4 FILLER_59_472 ();
 sg13g2_decap_8 FILLER_59_484 ();
 sg13g2_decap_8 FILLER_59_491 ();
 sg13g2_decap_8 FILLER_59_498 ();
 sg13g2_decap_8 FILLER_59_505 ();
 sg13g2_decap_8 FILLER_59_512 ();
 sg13g2_decap_4 FILLER_59_519 ();
 sg13g2_fill_1 FILLER_59_523 ();
 sg13g2_decap_8 FILLER_59_542 ();
 sg13g2_decap_8 FILLER_59_549 ();
 sg13g2_fill_2 FILLER_59_556 ();
 sg13g2_decap_8 FILLER_59_566 ();
 sg13g2_decap_8 FILLER_59_573 ();
 sg13g2_decap_8 FILLER_59_580 ();
 sg13g2_decap_8 FILLER_59_587 ();
 sg13g2_decap_8 FILLER_59_594 ();
 sg13g2_decap_8 FILLER_59_601 ();
 sg13g2_decap_8 FILLER_59_608 ();
 sg13g2_decap_8 FILLER_59_615 ();
 sg13g2_decap_8 FILLER_59_622 ();
 sg13g2_fill_1 FILLER_59_629 ();
 sg13g2_decap_4 FILLER_59_634 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_decap_4 FILLER_59_643 ();
 sg13g2_decap_8 FILLER_59_686 ();
 sg13g2_decap_4 FILLER_59_693 ();
 sg13g2_fill_2 FILLER_59_697 ();
 sg13g2_decap_8 FILLER_59_707 ();
 sg13g2_decap_8 FILLER_59_714 ();
 sg13g2_decap_8 FILLER_59_721 ();
 sg13g2_decap_4 FILLER_59_736 ();
 sg13g2_fill_1 FILLER_59_740 ();
 sg13g2_decap_8 FILLER_59_750 ();
 sg13g2_decap_8 FILLER_59_757 ();
 sg13g2_decap_8 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_771 ();
 sg13g2_decap_8 FILLER_59_778 ();
 sg13g2_fill_1 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_8 FILLER_59_797 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_856 ();
 sg13g2_decap_8 FILLER_59_863 ();
 sg13g2_decap_8 FILLER_59_870 ();
 sg13g2_fill_2 FILLER_59_877 ();
 sg13g2_fill_1 FILLER_59_879 ();
 sg13g2_decap_8 FILLER_59_893 ();
 sg13g2_decap_8 FILLER_59_900 ();
 sg13g2_decap_8 FILLER_59_907 ();
 sg13g2_decap_8 FILLER_59_914 ();
 sg13g2_decap_8 FILLER_59_921 ();
 sg13g2_decap_8 FILLER_59_928 ();
 sg13g2_decap_4 FILLER_59_935 ();
 sg13g2_fill_1 FILLER_59_939 ();
 sg13g2_fill_2 FILLER_59_958 ();
 sg13g2_fill_1 FILLER_59_960 ();
 sg13g2_decap_8 FILLER_59_973 ();
 sg13g2_decap_8 FILLER_59_980 ();
 sg13g2_decap_8 FILLER_59_987 ();
 sg13g2_decap_8 FILLER_59_994 ();
 sg13g2_decap_8 FILLER_59_1001 ();
 sg13g2_decap_8 FILLER_59_1008 ();
 sg13g2_decap_8 FILLER_59_1023 ();
 sg13g2_decap_8 FILLER_59_1030 ();
 sg13g2_decap_8 FILLER_59_1037 ();
 sg13g2_fill_2 FILLER_59_1044 ();
 sg13g2_decap_4 FILLER_59_1052 ();
 sg13g2_decap_8 FILLER_59_1064 ();
 sg13g2_decap_8 FILLER_59_1071 ();
 sg13g2_decap_8 FILLER_59_1078 ();
 sg13g2_decap_8 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1120 ();
 sg13g2_decap_8 FILLER_59_1127 ();
 sg13g2_fill_2 FILLER_59_1134 ();
 sg13g2_decap_8 FILLER_59_1153 ();
 sg13g2_decap_8 FILLER_59_1160 ();
 sg13g2_decap_8 FILLER_59_1167 ();
 sg13g2_decap_8 FILLER_59_1174 ();
 sg13g2_fill_1 FILLER_59_1181 ();
 sg13g2_fill_2 FILLER_59_1192 ();
 sg13g2_fill_1 FILLER_59_1194 ();
 sg13g2_fill_2 FILLER_59_1208 ();
 sg13g2_decap_8 FILLER_59_1221 ();
 sg13g2_decap_8 FILLER_59_1228 ();
 sg13g2_decap_8 FILLER_59_1235 ();
 sg13g2_decap_8 FILLER_59_1242 ();
 sg13g2_decap_8 FILLER_59_1249 ();
 sg13g2_decap_8 FILLER_59_1256 ();
 sg13g2_decap_8 FILLER_59_1263 ();
 sg13g2_decap_4 FILLER_59_1270 ();
 sg13g2_decap_8 FILLER_59_1286 ();
 sg13g2_decap_8 FILLER_59_1293 ();
 sg13g2_decap_8 FILLER_59_1300 ();
 sg13g2_decap_8 FILLER_59_1307 ();
 sg13g2_fill_1 FILLER_59_1314 ();
 sg13g2_decap_8 FILLER_59_1340 ();
 sg13g2_decap_4 FILLER_59_1347 ();
 sg13g2_fill_2 FILLER_59_1356 ();
 sg13g2_fill_1 FILLER_59_1358 ();
 sg13g2_decap_8 FILLER_59_1367 ();
 sg13g2_decap_8 FILLER_59_1374 ();
 sg13g2_fill_1 FILLER_59_1381 ();
 sg13g2_decap_8 FILLER_59_1402 ();
 sg13g2_decap_8 FILLER_59_1409 ();
 sg13g2_decap_8 FILLER_59_1416 ();
 sg13g2_decap_8 FILLER_59_1423 ();
 sg13g2_fill_1 FILLER_59_1442 ();
 sg13g2_decap_8 FILLER_59_1451 ();
 sg13g2_decap_8 FILLER_59_1458 ();
 sg13g2_decap_8 FILLER_59_1465 ();
 sg13g2_decap_8 FILLER_59_1472 ();
 sg13g2_fill_1 FILLER_59_1479 ();
 sg13g2_decap_4 FILLER_59_1488 ();
 sg13g2_fill_2 FILLER_59_1492 ();
 sg13g2_fill_1 FILLER_59_1502 ();
 sg13g2_decap_8 FILLER_59_1508 ();
 sg13g2_decap_8 FILLER_59_1515 ();
 sg13g2_decap_8 FILLER_59_1522 ();
 sg13g2_decap_8 FILLER_59_1541 ();
 sg13g2_decap_8 FILLER_59_1548 ();
 sg13g2_decap_4 FILLER_59_1555 ();
 sg13g2_fill_1 FILLER_59_1559 ();
 sg13g2_decap_4 FILLER_59_1575 ();
 sg13g2_fill_2 FILLER_59_1579 ();
 sg13g2_decap_8 FILLER_59_1597 ();
 sg13g2_decap_8 FILLER_59_1604 ();
 sg13g2_decap_8 FILLER_59_1611 ();
 sg13g2_decap_8 FILLER_59_1618 ();
 sg13g2_decap_8 FILLER_59_1625 ();
 sg13g2_decap_8 FILLER_59_1632 ();
 sg13g2_decap_8 FILLER_59_1639 ();
 sg13g2_decap_8 FILLER_59_1646 ();
 sg13g2_decap_8 FILLER_59_1653 ();
 sg13g2_decap_8 FILLER_59_1660 ();
 sg13g2_decap_8 FILLER_59_1667 ();
 sg13g2_decap_8 FILLER_59_1674 ();
 sg13g2_decap_8 FILLER_59_1681 ();
 sg13g2_decap_8 FILLER_59_1688 ();
 sg13g2_decap_8 FILLER_59_1695 ();
 sg13g2_decap_8 FILLER_59_1702 ();
 sg13g2_decap_8 FILLER_59_1709 ();
 sg13g2_decap_8 FILLER_59_1716 ();
 sg13g2_decap_8 FILLER_59_1723 ();
 sg13g2_decap_8 FILLER_59_1730 ();
 sg13g2_decap_8 FILLER_59_1737 ();
 sg13g2_decap_8 FILLER_59_1744 ();
 sg13g2_decap_8 FILLER_59_1751 ();
 sg13g2_decap_8 FILLER_59_1758 ();
 sg13g2_fill_2 FILLER_59_1765 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_110 ();
 sg13g2_decap_4 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_134 ();
 sg13g2_decap_4 FILLER_60_141 ();
 sg13g2_fill_2 FILLER_60_145 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_decap_8 FILLER_60_167 ();
 sg13g2_decap_8 FILLER_60_174 ();
 sg13g2_decap_8 FILLER_60_181 ();
 sg13g2_decap_8 FILLER_60_188 ();
 sg13g2_decap_4 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_199 ();
 sg13g2_decap_8 FILLER_60_215 ();
 sg13g2_decap_8 FILLER_60_222 ();
 sg13g2_decap_8 FILLER_60_229 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_decap_8 FILLER_60_243 ();
 sg13g2_decap_8 FILLER_60_250 ();
 sg13g2_decap_8 FILLER_60_257 ();
 sg13g2_decap_8 FILLER_60_264 ();
 sg13g2_decap_8 FILLER_60_271 ();
 sg13g2_decap_8 FILLER_60_278 ();
 sg13g2_fill_2 FILLER_60_285 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_302 ();
 sg13g2_decap_8 FILLER_60_309 ();
 sg13g2_decap_4 FILLER_60_316 ();
 sg13g2_fill_2 FILLER_60_320 ();
 sg13g2_decap_8 FILLER_60_330 ();
 sg13g2_decap_8 FILLER_60_337 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_60_380 ();
 sg13g2_decap_4 FILLER_60_387 ();
 sg13g2_fill_1 FILLER_60_391 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_decap_8 FILLER_60_407 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_434 ();
 sg13g2_fill_1 FILLER_60_436 ();
 sg13g2_decap_8 FILLER_60_445 ();
 sg13g2_decap_8 FILLER_60_452 ();
 sg13g2_decap_8 FILLER_60_459 ();
 sg13g2_decap_8 FILLER_60_466 ();
 sg13g2_decap_4 FILLER_60_473 ();
 sg13g2_decap_4 FILLER_60_485 ();
 sg13g2_fill_1 FILLER_60_497 ();
 sg13g2_decap_8 FILLER_60_503 ();
 sg13g2_decap_8 FILLER_60_510 ();
 sg13g2_decap_8 FILLER_60_517 ();
 sg13g2_decap_8 FILLER_60_524 ();
 sg13g2_decap_8 FILLER_60_531 ();
 sg13g2_decap_8 FILLER_60_538 ();
 sg13g2_decap_8 FILLER_60_545 ();
 sg13g2_fill_2 FILLER_60_552 ();
 sg13g2_decap_8 FILLER_60_562 ();
 sg13g2_decap_8 FILLER_60_569 ();
 sg13g2_decap_8 FILLER_60_576 ();
 sg13g2_decap_8 FILLER_60_583 ();
 sg13g2_decap_8 FILLER_60_606 ();
 sg13g2_decap_8 FILLER_60_613 ();
 sg13g2_decap_8 FILLER_60_620 ();
 sg13g2_decap_8 FILLER_60_627 ();
 sg13g2_decap_8 FILLER_60_634 ();
 sg13g2_decap_8 FILLER_60_641 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_decap_8 FILLER_60_683 ();
 sg13g2_decap_8 FILLER_60_690 ();
 sg13g2_decap_8 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_4 FILLER_60_711 ();
 sg13g2_fill_1 FILLER_60_715 ();
 sg13g2_decap_8 FILLER_60_734 ();
 sg13g2_decap_8 FILLER_60_741 ();
 sg13g2_decap_8 FILLER_60_748 ();
 sg13g2_decap_8 FILLER_60_755 ();
 sg13g2_decap_4 FILLER_60_762 ();
 sg13g2_fill_1 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_785 ();
 sg13g2_decap_8 FILLER_60_792 ();
 sg13g2_decap_8 FILLER_60_799 ();
 sg13g2_decap_8 FILLER_60_806 ();
 sg13g2_decap_8 FILLER_60_813 ();
 sg13g2_decap_8 FILLER_60_820 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_decap_8 FILLER_60_834 ();
 sg13g2_fill_2 FILLER_60_841 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_decap_4 FILLER_60_869 ();
 sg13g2_fill_2 FILLER_60_873 ();
 sg13g2_decap_8 FILLER_60_889 ();
 sg13g2_decap_8 FILLER_60_901 ();
 sg13g2_decap_8 FILLER_60_908 ();
 sg13g2_decap_8 FILLER_60_915 ();
 sg13g2_decap_8 FILLER_60_922 ();
 sg13g2_decap_8 FILLER_60_929 ();
 sg13g2_decap_8 FILLER_60_936 ();
 sg13g2_fill_1 FILLER_60_943 ();
 sg13g2_decap_4 FILLER_60_949 ();
 sg13g2_fill_2 FILLER_60_953 ();
 sg13g2_decap_8 FILLER_60_959 ();
 sg13g2_fill_2 FILLER_60_966 ();
 sg13g2_decap_8 FILLER_60_971 ();
 sg13g2_decap_8 FILLER_60_978 ();
 sg13g2_decap_8 FILLER_60_985 ();
 sg13g2_decap_8 FILLER_60_992 ();
 sg13g2_decap_8 FILLER_60_999 ();
 sg13g2_fill_1 FILLER_60_1006 ();
 sg13g2_decap_8 FILLER_60_1013 ();
 sg13g2_decap_8 FILLER_60_1028 ();
 sg13g2_decap_8 FILLER_60_1035 ();
 sg13g2_fill_2 FILLER_60_1050 ();
 sg13g2_decap_8 FILLER_60_1068 ();
 sg13g2_decap_8 FILLER_60_1075 ();
 sg13g2_decap_8 FILLER_60_1082 ();
 sg13g2_decap_4 FILLER_60_1089 ();
 sg13g2_decap_8 FILLER_60_1096 ();
 sg13g2_decap_8 FILLER_60_1103 ();
 sg13g2_decap_8 FILLER_60_1110 ();
 sg13g2_decap_8 FILLER_60_1117 ();
 sg13g2_decap_8 FILLER_60_1124 ();
 sg13g2_decap_8 FILLER_60_1131 ();
 sg13g2_decap_8 FILLER_60_1138 ();
 sg13g2_fill_2 FILLER_60_1145 ();
 sg13g2_fill_1 FILLER_60_1147 ();
 sg13g2_fill_2 FILLER_60_1159 ();
 sg13g2_decap_8 FILLER_60_1166 ();
 sg13g2_decap_8 FILLER_60_1173 ();
 sg13g2_decap_8 FILLER_60_1180 ();
 sg13g2_fill_2 FILLER_60_1187 ();
 sg13g2_decap_4 FILLER_60_1205 ();
 sg13g2_fill_1 FILLER_60_1209 ();
 sg13g2_decap_8 FILLER_60_1213 ();
 sg13g2_decap_8 FILLER_60_1220 ();
 sg13g2_decap_8 FILLER_60_1227 ();
 sg13g2_fill_1 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1239 ();
 sg13g2_decap_8 FILLER_60_1246 ();
 sg13g2_decap_4 FILLER_60_1253 ();
 sg13g2_decap_4 FILLER_60_1272 ();
 sg13g2_decap_8 FILLER_60_1284 ();
 sg13g2_decap_8 FILLER_60_1291 ();
 sg13g2_decap_8 FILLER_60_1298 ();
 sg13g2_decap_8 FILLER_60_1305 ();
 sg13g2_decap_8 FILLER_60_1312 ();
 sg13g2_fill_2 FILLER_60_1319 ();
 sg13g2_fill_1 FILLER_60_1321 ();
 sg13g2_decap_8 FILLER_60_1335 ();
 sg13g2_decap_8 FILLER_60_1342 ();
 sg13g2_fill_2 FILLER_60_1349 ();
 sg13g2_decap_8 FILLER_60_1360 ();
 sg13g2_decap_8 FILLER_60_1367 ();
 sg13g2_decap_8 FILLER_60_1374 ();
 sg13g2_decap_8 FILLER_60_1381 ();
 sg13g2_fill_1 FILLER_60_1388 ();
 sg13g2_decap_8 FILLER_60_1397 ();
 sg13g2_decap_8 FILLER_60_1404 ();
 sg13g2_decap_8 FILLER_60_1411 ();
 sg13g2_decap_8 FILLER_60_1418 ();
 sg13g2_decap_4 FILLER_60_1425 ();
 sg13g2_fill_2 FILLER_60_1437 ();
 sg13g2_decap_8 FILLER_60_1452 ();
 sg13g2_decap_8 FILLER_60_1459 ();
 sg13g2_decap_8 FILLER_60_1466 ();
 sg13g2_decap_8 FILLER_60_1473 ();
 sg13g2_decap_8 FILLER_60_1480 ();
 sg13g2_decap_8 FILLER_60_1487 ();
 sg13g2_decap_4 FILLER_60_1494 ();
 sg13g2_fill_2 FILLER_60_1498 ();
 sg13g2_decap_8 FILLER_60_1510 ();
 sg13g2_decap_8 FILLER_60_1517 ();
 sg13g2_decap_8 FILLER_60_1524 ();
 sg13g2_decap_8 FILLER_60_1531 ();
 sg13g2_decap_8 FILLER_60_1538 ();
 sg13g2_fill_2 FILLER_60_1545 ();
 sg13g2_decap_8 FILLER_60_1555 ();
 sg13g2_fill_1 FILLER_60_1562 ();
 sg13g2_decap_8 FILLER_60_1568 ();
 sg13g2_fill_2 FILLER_60_1575 ();
 sg13g2_fill_1 FILLER_60_1577 ();
 sg13g2_decap_8 FILLER_60_1599 ();
 sg13g2_decap_8 FILLER_60_1606 ();
 sg13g2_decap_8 FILLER_60_1613 ();
 sg13g2_decap_8 FILLER_60_1620 ();
 sg13g2_decap_8 FILLER_60_1627 ();
 sg13g2_decap_8 FILLER_60_1634 ();
 sg13g2_decap_8 FILLER_60_1641 ();
 sg13g2_decap_8 FILLER_60_1648 ();
 sg13g2_decap_8 FILLER_60_1655 ();
 sg13g2_decap_8 FILLER_60_1662 ();
 sg13g2_decap_8 FILLER_60_1669 ();
 sg13g2_decap_8 FILLER_60_1676 ();
 sg13g2_decap_8 FILLER_60_1683 ();
 sg13g2_decap_8 FILLER_60_1690 ();
 sg13g2_decap_8 FILLER_60_1697 ();
 sg13g2_decap_8 FILLER_60_1704 ();
 sg13g2_decap_8 FILLER_60_1711 ();
 sg13g2_decap_8 FILLER_60_1718 ();
 sg13g2_decap_8 FILLER_60_1725 ();
 sg13g2_decap_8 FILLER_60_1732 ();
 sg13g2_decap_8 FILLER_60_1739 ();
 sg13g2_decap_8 FILLER_60_1746 ();
 sg13g2_decap_8 FILLER_60_1753 ();
 sg13g2_decap_8 FILLER_60_1760 ();
 sg13g2_fill_1 FILLER_60_1767 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_75 ();
 sg13g2_decap_8 FILLER_61_82 ();
 sg13g2_decap_4 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_93 ();
 sg13g2_decap_8 FILLER_61_99 ();
 sg13g2_decap_8 FILLER_61_106 ();
 sg13g2_fill_2 FILLER_61_113 ();
 sg13g2_decap_8 FILLER_61_120 ();
 sg13g2_decap_8 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_134 ();
 sg13g2_decap_8 FILLER_61_141 ();
 sg13g2_decap_8 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_155 ();
 sg13g2_decap_8 FILLER_61_162 ();
 sg13g2_decap_8 FILLER_61_169 ();
 sg13g2_decap_8 FILLER_61_176 ();
 sg13g2_decap_8 FILLER_61_183 ();
 sg13g2_decap_8 FILLER_61_190 ();
 sg13g2_fill_1 FILLER_61_197 ();
 sg13g2_decap_8 FILLER_61_208 ();
 sg13g2_decap_8 FILLER_61_215 ();
 sg13g2_decap_8 FILLER_61_222 ();
 sg13g2_decap_8 FILLER_61_229 ();
 sg13g2_decap_8 FILLER_61_236 ();
 sg13g2_decap_8 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_decap_8 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_278 ();
 sg13g2_decap_8 FILLER_61_285 ();
 sg13g2_decap_4 FILLER_61_292 ();
 sg13g2_fill_2 FILLER_61_296 ();
 sg13g2_decap_8 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_decap_8 FILLER_61_328 ();
 sg13g2_decap_8 FILLER_61_335 ();
 sg13g2_decap_8 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_2 FILLER_61_433 ();
 sg13g2_decap_8 FILLER_61_447 ();
 sg13g2_decap_8 FILLER_61_454 ();
 sg13g2_fill_2 FILLER_61_461 ();
 sg13g2_fill_1 FILLER_61_463 ();
 sg13g2_fill_2 FILLER_61_487 ();
 sg13g2_decap_8 FILLER_61_506 ();
 sg13g2_decap_8 FILLER_61_513 ();
 sg13g2_decap_8 FILLER_61_520 ();
 sg13g2_decap_4 FILLER_61_527 ();
 sg13g2_decap_8 FILLER_61_543 ();
 sg13g2_decap_8 FILLER_61_550 ();
 sg13g2_decap_8 FILLER_61_557 ();
 sg13g2_decap_8 FILLER_61_564 ();
 sg13g2_decap_8 FILLER_61_571 ();
 sg13g2_decap_8 FILLER_61_578 ();
 sg13g2_decap_4 FILLER_61_585 ();
 sg13g2_decap_8 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_617 ();
 sg13g2_decap_8 FILLER_61_626 ();
 sg13g2_decap_8 FILLER_61_633 ();
 sg13g2_decap_8 FILLER_61_640 ();
 sg13g2_decap_8 FILLER_61_647 ();
 sg13g2_decap_8 FILLER_61_654 ();
 sg13g2_decap_8 FILLER_61_661 ();
 sg13g2_decap_8 FILLER_61_668 ();
 sg13g2_decap_8 FILLER_61_675 ();
 sg13g2_decap_8 FILLER_61_682 ();
 sg13g2_decap_8 FILLER_61_689 ();
 sg13g2_decap_8 FILLER_61_696 ();
 sg13g2_decap_8 FILLER_61_703 ();
 sg13g2_decap_8 FILLER_61_710 ();
 sg13g2_decap_8 FILLER_61_717 ();
 sg13g2_decap_8 FILLER_61_724 ();
 sg13g2_decap_8 FILLER_61_731 ();
 sg13g2_decap_8 FILLER_61_738 ();
 sg13g2_decap_8 FILLER_61_745 ();
 sg13g2_decap_4 FILLER_61_752 ();
 sg13g2_fill_1 FILLER_61_756 ();
 sg13g2_decap_8 FILLER_61_777 ();
 sg13g2_decap_8 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_791 ();
 sg13g2_decap_8 FILLER_61_798 ();
 sg13g2_fill_1 FILLER_61_805 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_fill_2 FILLER_61_838 ();
 sg13g2_fill_1 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_61_857 ();
 sg13g2_decap_8 FILLER_61_864 ();
 sg13g2_decap_8 FILLER_61_871 ();
 sg13g2_decap_8 FILLER_61_878 ();
 sg13g2_decap_8 FILLER_61_885 ();
 sg13g2_fill_1 FILLER_61_892 ();
 sg13g2_decap_8 FILLER_61_917 ();
 sg13g2_decap_8 FILLER_61_924 ();
 sg13g2_decap_4 FILLER_61_931 ();
 sg13g2_decap_8 FILLER_61_948 ();
 sg13g2_decap_8 FILLER_61_955 ();
 sg13g2_decap_4 FILLER_61_962 ();
 sg13g2_fill_2 FILLER_61_966 ();
 sg13g2_decap_8 FILLER_61_980 ();
 sg13g2_decap_8 FILLER_61_987 ();
 sg13g2_decap_4 FILLER_61_994 ();
 sg13g2_fill_2 FILLER_61_1008 ();
 sg13g2_fill_2 FILLER_61_1023 ();
 sg13g2_decap_4 FILLER_61_1046 ();
 sg13g2_fill_1 FILLER_61_1050 ();
 sg13g2_decap_8 FILLER_61_1062 ();
 sg13g2_decap_4 FILLER_61_1077 ();
 sg13g2_decap_4 FILLER_61_1094 ();
 sg13g2_fill_1 FILLER_61_1098 ();
 sg13g2_fill_2 FILLER_61_1125 ();
 sg13g2_decap_8 FILLER_61_1135 ();
 sg13g2_fill_1 FILLER_61_1142 ();
 sg13g2_decap_4 FILLER_61_1148 ();
 sg13g2_fill_1 FILLER_61_1152 ();
 sg13g2_decap_8 FILLER_61_1157 ();
 sg13g2_decap_8 FILLER_61_1164 ();
 sg13g2_decap_8 FILLER_61_1171 ();
 sg13g2_decap_8 FILLER_61_1178 ();
 sg13g2_fill_2 FILLER_61_1193 ();
 sg13g2_decap_8 FILLER_61_1217 ();
 sg13g2_decap_8 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1236 ();
 sg13g2_decap_4 FILLER_61_1243 ();
 sg13g2_fill_1 FILLER_61_1247 ();
 sg13g2_fill_1 FILLER_61_1262 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_8 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_decap_8 FILLER_61_1299 ();
 sg13g2_decap_4 FILLER_61_1306 ();
 sg13g2_fill_1 FILLER_61_1310 ();
 sg13g2_decap_8 FILLER_61_1327 ();
 sg13g2_decap_8 FILLER_61_1334 ();
 sg13g2_decap_8 FILLER_61_1341 ();
 sg13g2_decap_8 FILLER_61_1348 ();
 sg13g2_decap_8 FILLER_61_1355 ();
 sg13g2_decap_8 FILLER_61_1362 ();
 sg13g2_decap_8 FILLER_61_1369 ();
 sg13g2_decap_8 FILLER_61_1376 ();
 sg13g2_decap_8 FILLER_61_1383 ();
 sg13g2_decap_4 FILLER_61_1390 ();
 sg13g2_decap_8 FILLER_61_1414 ();
 sg13g2_decap_8 FILLER_61_1421 ();
 sg13g2_decap_8 FILLER_61_1428 ();
 sg13g2_decap_8 FILLER_61_1435 ();
 sg13g2_fill_2 FILLER_61_1442 ();
 sg13g2_fill_2 FILLER_61_1448 ();
 sg13g2_decap_8 FILLER_61_1454 ();
 sg13g2_fill_1 FILLER_61_1461 ();
 sg13g2_fill_2 FILLER_61_1467 ();
 sg13g2_decap_8 FILLER_61_1474 ();
 sg13g2_fill_2 FILLER_61_1481 ();
 sg13g2_fill_1 FILLER_61_1483 ();
 sg13g2_decap_8 FILLER_61_1489 ();
 sg13g2_decap_8 FILLER_61_1496 ();
 sg13g2_decap_8 FILLER_61_1503 ();
 sg13g2_decap_8 FILLER_61_1510 ();
 sg13g2_decap_8 FILLER_61_1517 ();
 sg13g2_fill_2 FILLER_61_1524 ();
 sg13g2_fill_1 FILLER_61_1526 ();
 sg13g2_decap_8 FILLER_61_1557 ();
 sg13g2_decap_8 FILLER_61_1564 ();
 sg13g2_fill_2 FILLER_61_1571 ();
 sg13g2_fill_1 FILLER_61_1573 ();
 sg13g2_decap_8 FILLER_61_1579 ();
 sg13g2_decap_4 FILLER_61_1586 ();
 sg13g2_fill_1 FILLER_61_1590 ();
 sg13g2_decap_8 FILLER_61_1599 ();
 sg13g2_decap_8 FILLER_61_1606 ();
 sg13g2_decap_8 FILLER_61_1613 ();
 sg13g2_decap_8 FILLER_61_1620 ();
 sg13g2_decap_8 FILLER_61_1627 ();
 sg13g2_decap_8 FILLER_61_1634 ();
 sg13g2_decap_4 FILLER_61_1641 ();
 sg13g2_decap_8 FILLER_61_1654 ();
 sg13g2_decap_8 FILLER_61_1661 ();
 sg13g2_decap_8 FILLER_61_1668 ();
 sg13g2_decap_8 FILLER_61_1675 ();
 sg13g2_decap_8 FILLER_61_1682 ();
 sg13g2_decap_8 FILLER_61_1689 ();
 sg13g2_decap_8 FILLER_61_1696 ();
 sg13g2_decap_8 FILLER_61_1703 ();
 sg13g2_decap_8 FILLER_61_1710 ();
 sg13g2_decap_8 FILLER_61_1717 ();
 sg13g2_decap_8 FILLER_61_1724 ();
 sg13g2_decap_8 FILLER_61_1731 ();
 sg13g2_decap_8 FILLER_61_1738 ();
 sg13g2_decap_8 FILLER_61_1745 ();
 sg13g2_decap_8 FILLER_61_1752 ();
 sg13g2_decap_8 FILLER_61_1759 ();
 sg13g2_fill_2 FILLER_61_1766 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_128 ();
 sg13g2_decap_8 FILLER_62_135 ();
 sg13g2_decap_4 FILLER_62_142 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_decap_8 FILLER_62_155 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_decap_8 FILLER_62_169 ();
 sg13g2_decap_8 FILLER_62_176 ();
 sg13g2_decap_8 FILLER_62_183 ();
 sg13g2_decap_8 FILLER_62_190 ();
 sg13g2_decap_8 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_204 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_239 ();
 sg13g2_decap_8 FILLER_62_246 ();
 sg13g2_decap_8 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_260 ();
 sg13g2_decap_8 FILLER_62_267 ();
 sg13g2_fill_2 FILLER_62_274 ();
 sg13g2_fill_1 FILLER_62_276 ();
 sg13g2_decap_8 FILLER_62_285 ();
 sg13g2_decap_8 FILLER_62_292 ();
 sg13g2_decap_8 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_306 ();
 sg13g2_decap_8 FILLER_62_317 ();
 sg13g2_decap_4 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_328 ();
 sg13g2_decap_8 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_decap_4 FILLER_62_351 ();
 sg13g2_fill_1 FILLER_62_355 ();
 sg13g2_decap_8 FILLER_62_360 ();
 sg13g2_fill_2 FILLER_62_367 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_decap_8 FILLER_62_409 ();
 sg13g2_decap_8 FILLER_62_416 ();
 sg13g2_decap_8 FILLER_62_423 ();
 sg13g2_decap_8 FILLER_62_430 ();
 sg13g2_decap_8 FILLER_62_437 ();
 sg13g2_decap_4 FILLER_62_444 ();
 sg13g2_fill_1 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_457 ();
 sg13g2_decap_8 FILLER_62_464 ();
 sg13g2_decap_8 FILLER_62_471 ();
 sg13g2_decap_8 FILLER_62_478 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_fill_1 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_decap_8 FILLER_62_531 ();
 sg13g2_decap_8 FILLER_62_538 ();
 sg13g2_decap_8 FILLER_62_545 ();
 sg13g2_decap_4 FILLER_62_552 ();
 sg13g2_fill_2 FILLER_62_556 ();
 sg13g2_fill_1 FILLER_62_562 ();
 sg13g2_decap_8 FILLER_62_571 ();
 sg13g2_decap_8 FILLER_62_578 ();
 sg13g2_decap_8 FILLER_62_585 ();
 sg13g2_fill_1 FILLER_62_592 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_1 FILLER_62_619 ();
 sg13g2_decap_8 FILLER_62_634 ();
 sg13g2_decap_8 FILLER_62_641 ();
 sg13g2_decap_8 FILLER_62_648 ();
 sg13g2_decap_8 FILLER_62_655 ();
 sg13g2_decap_4 FILLER_62_662 ();
 sg13g2_decap_8 FILLER_62_677 ();
 sg13g2_decap_8 FILLER_62_684 ();
 sg13g2_decap_8 FILLER_62_691 ();
 sg13g2_fill_2 FILLER_62_698 ();
 sg13g2_fill_1 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_709 ();
 sg13g2_decap_8 FILLER_62_716 ();
 sg13g2_decap_8 FILLER_62_723 ();
 sg13g2_decap_8 FILLER_62_730 ();
 sg13g2_decap_8 FILLER_62_737 ();
 sg13g2_decap_4 FILLER_62_744 ();
 sg13g2_fill_2 FILLER_62_748 ();
 sg13g2_decap_8 FILLER_62_780 ();
 sg13g2_decap_8 FILLER_62_787 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_decap_4 FILLER_62_801 ();
 sg13g2_fill_2 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_815 ();
 sg13g2_decap_4 FILLER_62_822 ();
 sg13g2_fill_1 FILLER_62_826 ();
 sg13g2_decap_4 FILLER_62_835 ();
 sg13g2_fill_2 FILLER_62_839 ();
 sg13g2_decap_8 FILLER_62_853 ();
 sg13g2_decap_8 FILLER_62_860 ();
 sg13g2_decap_8 FILLER_62_867 ();
 sg13g2_decap_8 FILLER_62_874 ();
 sg13g2_decap_8 FILLER_62_881 ();
 sg13g2_decap_8 FILLER_62_914 ();
 sg13g2_decap_8 FILLER_62_921 ();
 sg13g2_decap_8 FILLER_62_928 ();
 sg13g2_fill_1 FILLER_62_935 ();
 sg13g2_decap_8 FILLER_62_953 ();
 sg13g2_fill_1 FILLER_62_960 ();
 sg13g2_decap_8 FILLER_62_977 ();
 sg13g2_decap_8 FILLER_62_984 ();
 sg13g2_decap_8 FILLER_62_991 ();
 sg13g2_decap_8 FILLER_62_998 ();
 sg13g2_decap_4 FILLER_62_1005 ();
 sg13g2_fill_1 FILLER_62_1009 ();
 sg13g2_decap_8 FILLER_62_1027 ();
 sg13g2_decap_8 FILLER_62_1034 ();
 sg13g2_decap_8 FILLER_62_1041 ();
 sg13g2_decap_8 FILLER_62_1048 ();
 sg13g2_decap_8 FILLER_62_1055 ();
 sg13g2_decap_8 FILLER_62_1062 ();
 sg13g2_decap_8 FILLER_62_1090 ();
 sg13g2_decap_8 FILLER_62_1097 ();
 sg13g2_decap_4 FILLER_62_1104 ();
 sg13g2_fill_2 FILLER_62_1108 ();
 sg13g2_decap_8 FILLER_62_1114 ();
 sg13g2_decap_8 FILLER_62_1121 ();
 sg13g2_decap_8 FILLER_62_1128 ();
 sg13g2_decap_8 FILLER_62_1135 ();
 sg13g2_decap_8 FILLER_62_1142 ();
 sg13g2_decap_8 FILLER_62_1149 ();
 sg13g2_decap_4 FILLER_62_1156 ();
 sg13g2_fill_1 FILLER_62_1160 ();
 sg13g2_decap_8 FILLER_62_1169 ();
 sg13g2_decap_8 FILLER_62_1176 ();
 sg13g2_decap_8 FILLER_62_1183 ();
 sg13g2_decap_4 FILLER_62_1190 ();
 sg13g2_decap_8 FILLER_62_1202 ();
 sg13g2_decap_8 FILLER_62_1209 ();
 sg13g2_decap_8 FILLER_62_1216 ();
 sg13g2_decap_8 FILLER_62_1223 ();
 sg13g2_decap_8 FILLER_62_1230 ();
 sg13g2_decap_8 FILLER_62_1237 ();
 sg13g2_fill_2 FILLER_62_1244 ();
 sg13g2_fill_1 FILLER_62_1246 ();
 sg13g2_decap_8 FILLER_62_1270 ();
 sg13g2_decap_8 FILLER_62_1277 ();
 sg13g2_decap_8 FILLER_62_1284 ();
 sg13g2_decap_8 FILLER_62_1291 ();
 sg13g2_decap_8 FILLER_62_1298 ();
 sg13g2_decap_4 FILLER_62_1305 ();
 sg13g2_fill_2 FILLER_62_1309 ();
 sg13g2_decap_8 FILLER_62_1322 ();
 sg13g2_decap_8 FILLER_62_1329 ();
 sg13g2_fill_2 FILLER_62_1344 ();
 sg13g2_decap_8 FILLER_62_1351 ();
 sg13g2_decap_8 FILLER_62_1358 ();
 sg13g2_decap_8 FILLER_62_1365 ();
 sg13g2_decap_8 FILLER_62_1372 ();
 sg13g2_decap_8 FILLER_62_1379 ();
 sg13g2_decap_8 FILLER_62_1386 ();
 sg13g2_fill_1 FILLER_62_1393 ();
 sg13g2_decap_8 FILLER_62_1403 ();
 sg13g2_decap_8 FILLER_62_1410 ();
 sg13g2_decap_8 FILLER_62_1417 ();
 sg13g2_decap_8 FILLER_62_1424 ();
 sg13g2_decap_4 FILLER_62_1431 ();
 sg13g2_fill_2 FILLER_62_1435 ();
 sg13g2_fill_1 FILLER_62_1461 ();
 sg13g2_fill_1 FILLER_62_1478 ();
 sg13g2_decap_8 FILLER_62_1503 ();
 sg13g2_decap_8 FILLER_62_1510 ();
 sg13g2_decap_8 FILLER_62_1517 ();
 sg13g2_fill_2 FILLER_62_1524 ();
 sg13g2_decap_8 FILLER_62_1538 ();
 sg13g2_decap_4 FILLER_62_1545 ();
 sg13g2_decap_8 FILLER_62_1558 ();
 sg13g2_fill_2 FILLER_62_1565 ();
 sg13g2_fill_1 FILLER_62_1567 ();
 sg13g2_decap_8 FILLER_62_1584 ();
 sg13g2_decap_8 FILLER_62_1591 ();
 sg13g2_decap_8 FILLER_62_1598 ();
 sg13g2_decap_8 FILLER_62_1605 ();
 sg13g2_decap_4 FILLER_62_1612 ();
 sg13g2_fill_2 FILLER_62_1616 ();
 sg13g2_decap_8 FILLER_62_1669 ();
 sg13g2_decap_8 FILLER_62_1676 ();
 sg13g2_decap_8 FILLER_62_1683 ();
 sg13g2_decap_8 FILLER_62_1690 ();
 sg13g2_decap_8 FILLER_62_1697 ();
 sg13g2_decap_8 FILLER_62_1704 ();
 sg13g2_decap_8 FILLER_62_1711 ();
 sg13g2_decap_8 FILLER_62_1718 ();
 sg13g2_decap_8 FILLER_62_1725 ();
 sg13g2_decap_8 FILLER_62_1732 ();
 sg13g2_decap_8 FILLER_62_1739 ();
 sg13g2_decap_8 FILLER_62_1746 ();
 sg13g2_decap_8 FILLER_62_1753 ();
 sg13g2_decap_8 FILLER_62_1760 ();
 sg13g2_fill_1 FILLER_62_1767 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_74 ();
 sg13g2_decap_8 FILLER_63_81 ();
 sg13g2_decap_8 FILLER_63_88 ();
 sg13g2_decap_8 FILLER_63_95 ();
 sg13g2_fill_2 FILLER_63_102 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_decap_8 FILLER_63_131 ();
 sg13g2_decap_8 FILLER_63_138 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_152 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_decap_8 FILLER_63_166 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_178 ();
 sg13g2_decap_8 FILLER_63_185 ();
 sg13g2_decap_8 FILLER_63_192 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_fill_1 FILLER_63_247 ();
 sg13g2_decap_8 FILLER_63_261 ();
 sg13g2_decap_4 FILLER_63_268 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_decap_4 FILLER_63_297 ();
 sg13g2_fill_2 FILLER_63_301 ();
 sg13g2_fill_1 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_335 ();
 sg13g2_decap_8 FILLER_63_342 ();
 sg13g2_decap_8 FILLER_63_349 ();
 sg13g2_decap_8 FILLER_63_356 ();
 sg13g2_decap_8 FILLER_63_363 ();
 sg13g2_decap_8 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_8 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_decap_8 FILLER_63_405 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_decap_8 FILLER_63_421 ();
 sg13g2_decap_8 FILLER_63_428 ();
 sg13g2_decap_4 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_439 ();
 sg13g2_decap_8 FILLER_63_454 ();
 sg13g2_decap_8 FILLER_63_461 ();
 sg13g2_decap_8 FILLER_63_468 ();
 sg13g2_decap_8 FILLER_63_475 ();
 sg13g2_decap_8 FILLER_63_482 ();
 sg13g2_decap_8 FILLER_63_489 ();
 sg13g2_decap_8 FILLER_63_521 ();
 sg13g2_decap_8 FILLER_63_528 ();
 sg13g2_decap_8 FILLER_63_535 ();
 sg13g2_fill_2 FILLER_63_542 ();
 sg13g2_fill_1 FILLER_63_544 ();
 sg13g2_decap_8 FILLER_63_580 ();
 sg13g2_decap_8 FILLER_63_587 ();
 sg13g2_decap_4 FILLER_63_594 ();
 sg13g2_fill_2 FILLER_63_602 ();
 sg13g2_fill_1 FILLER_63_623 ();
 sg13g2_fill_1 FILLER_63_632 ();
 sg13g2_decap_8 FILLER_63_640 ();
 sg13g2_decap_8 FILLER_63_647 ();
 sg13g2_decap_8 FILLER_63_654 ();
 sg13g2_fill_1 FILLER_63_661 ();
 sg13g2_decap_8 FILLER_63_688 ();
 sg13g2_fill_1 FILLER_63_695 ();
 sg13g2_decap_8 FILLER_63_713 ();
 sg13g2_decap_8 FILLER_63_720 ();
 sg13g2_fill_2 FILLER_63_727 ();
 sg13g2_fill_1 FILLER_63_729 ();
 sg13g2_fill_1 FILLER_63_743 ();
 sg13g2_decap_4 FILLER_63_750 ();
 sg13g2_fill_2 FILLER_63_754 ();
 sg13g2_decap_8 FILLER_63_771 ();
 sg13g2_decap_8 FILLER_63_778 ();
 sg13g2_decap_8 FILLER_63_785 ();
 sg13g2_decap_8 FILLER_63_792 ();
 sg13g2_decap_8 FILLER_63_799 ();
 sg13g2_decap_8 FILLER_63_822 ();
 sg13g2_decap_4 FILLER_63_829 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_decap_8 FILLER_63_859 ();
 sg13g2_decap_8 FILLER_63_866 ();
 sg13g2_decap_8 FILLER_63_873 ();
 sg13g2_decap_4 FILLER_63_880 ();
 sg13g2_fill_2 FILLER_63_884 ();
 sg13g2_decap_8 FILLER_63_891 ();
 sg13g2_decap_4 FILLER_63_898 ();
 sg13g2_fill_1 FILLER_63_902 ();
 sg13g2_decap_8 FILLER_63_912 ();
 sg13g2_decap_8 FILLER_63_919 ();
 sg13g2_decap_8 FILLER_63_926 ();
 sg13g2_decap_8 FILLER_63_933 ();
 sg13g2_decap_8 FILLER_63_940 ();
 sg13g2_decap_4 FILLER_63_947 ();
 sg13g2_fill_1 FILLER_63_951 ();
 sg13g2_fill_2 FILLER_63_976 ();
 sg13g2_fill_1 FILLER_63_978 ();
 sg13g2_decap_8 FILLER_63_987 ();
 sg13g2_decap_4 FILLER_63_994 ();
 sg13g2_fill_2 FILLER_63_998 ();
 sg13g2_decap_4 FILLER_63_1008 ();
 sg13g2_decap_8 FILLER_63_1024 ();
 sg13g2_decap_8 FILLER_63_1031 ();
 sg13g2_decap_8 FILLER_63_1038 ();
 sg13g2_decap_8 FILLER_63_1045 ();
 sg13g2_decap_8 FILLER_63_1052 ();
 sg13g2_decap_8 FILLER_63_1059 ();
 sg13g2_decap_8 FILLER_63_1066 ();
 sg13g2_decap_8 FILLER_63_1073 ();
 sg13g2_fill_2 FILLER_63_1080 ();
 sg13g2_fill_1 FILLER_63_1082 ();
 sg13g2_decap_8 FILLER_63_1091 ();
 sg13g2_decap_8 FILLER_63_1098 ();
 sg13g2_decap_8 FILLER_63_1105 ();
 sg13g2_decap_8 FILLER_63_1112 ();
 sg13g2_fill_2 FILLER_63_1119 ();
 sg13g2_decap_4 FILLER_63_1133 ();
 sg13g2_fill_2 FILLER_63_1137 ();
 sg13g2_fill_2 FILLER_63_1143 ();
 sg13g2_fill_1 FILLER_63_1145 ();
 sg13g2_decap_8 FILLER_63_1154 ();
 sg13g2_decap_8 FILLER_63_1166 ();
 sg13g2_decap_8 FILLER_63_1173 ();
 sg13g2_decap_8 FILLER_63_1180 ();
 sg13g2_decap_4 FILLER_63_1187 ();
 sg13g2_fill_1 FILLER_63_1194 ();
 sg13g2_decap_8 FILLER_63_1212 ();
 sg13g2_decap_8 FILLER_63_1219 ();
 sg13g2_decap_8 FILLER_63_1226 ();
 sg13g2_decap_8 FILLER_63_1233 ();
 sg13g2_fill_2 FILLER_63_1240 ();
 sg13g2_decap_4 FILLER_63_1246 ();
 sg13g2_fill_1 FILLER_63_1250 ();
 sg13g2_decap_8 FILLER_63_1264 ();
 sg13g2_decap_8 FILLER_63_1271 ();
 sg13g2_decap_8 FILLER_63_1278 ();
 sg13g2_decap_8 FILLER_63_1285 ();
 sg13g2_fill_2 FILLER_63_1292 ();
 sg13g2_fill_1 FILLER_63_1294 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_4 FILLER_63_1310 ();
 sg13g2_fill_1 FILLER_63_1318 ();
 sg13g2_decap_4 FILLER_63_1327 ();
 sg13g2_decap_4 FILLER_63_1335 ();
 sg13g2_fill_1 FILLER_63_1339 ();
 sg13g2_decap_8 FILLER_63_1356 ();
 sg13g2_decap_8 FILLER_63_1363 ();
 sg13g2_fill_1 FILLER_63_1370 ();
 sg13g2_decap_8 FILLER_63_1379 ();
 sg13g2_fill_2 FILLER_63_1386 ();
 sg13g2_decap_8 FILLER_63_1396 ();
 sg13g2_decap_8 FILLER_63_1403 ();
 sg13g2_decap_8 FILLER_63_1410 ();
 sg13g2_decap_8 FILLER_63_1417 ();
 sg13g2_decap_8 FILLER_63_1424 ();
 sg13g2_decap_8 FILLER_63_1431 ();
 sg13g2_decap_8 FILLER_63_1438 ();
 sg13g2_decap_8 FILLER_63_1445 ();
 sg13g2_decap_8 FILLER_63_1452 ();
 sg13g2_decap_4 FILLER_63_1459 ();
 sg13g2_decap_8 FILLER_63_1468 ();
 sg13g2_decap_8 FILLER_63_1475 ();
 sg13g2_decap_8 FILLER_63_1482 ();
 sg13g2_decap_8 FILLER_63_1489 ();
 sg13g2_decap_8 FILLER_63_1496 ();
 sg13g2_decap_8 FILLER_63_1503 ();
 sg13g2_decap_8 FILLER_63_1510 ();
 sg13g2_fill_1 FILLER_63_1517 ();
 sg13g2_decap_8 FILLER_63_1535 ();
 sg13g2_decap_8 FILLER_63_1542 ();
 sg13g2_decap_8 FILLER_63_1549 ();
 sg13g2_decap_8 FILLER_63_1556 ();
 sg13g2_decap_8 FILLER_63_1563 ();
 sg13g2_decap_8 FILLER_63_1570 ();
 sg13g2_decap_8 FILLER_63_1577 ();
 sg13g2_decap_8 FILLER_63_1584 ();
 sg13g2_decap_8 FILLER_63_1591 ();
 sg13g2_decap_8 FILLER_63_1598 ();
 sg13g2_fill_2 FILLER_63_1605 ();
 sg13g2_decap_8 FILLER_63_1619 ();
 sg13g2_fill_2 FILLER_63_1626 ();
 sg13g2_fill_1 FILLER_63_1628 ();
 sg13g2_decap_8 FILLER_63_1633 ();
 sg13g2_decap_8 FILLER_63_1640 ();
 sg13g2_fill_1 FILLER_63_1647 ();
 sg13g2_decap_8 FILLER_63_1654 ();
 sg13g2_decap_8 FILLER_63_1661 ();
 sg13g2_decap_8 FILLER_63_1668 ();
 sg13g2_decap_8 FILLER_63_1675 ();
 sg13g2_decap_8 FILLER_63_1682 ();
 sg13g2_decap_8 FILLER_63_1689 ();
 sg13g2_decap_8 FILLER_63_1696 ();
 sg13g2_decap_8 FILLER_63_1703 ();
 sg13g2_decap_8 FILLER_63_1710 ();
 sg13g2_decap_8 FILLER_63_1717 ();
 sg13g2_decap_8 FILLER_63_1724 ();
 sg13g2_decap_8 FILLER_63_1731 ();
 sg13g2_decap_8 FILLER_63_1738 ();
 sg13g2_decap_8 FILLER_63_1745 ();
 sg13g2_decap_8 FILLER_63_1752 ();
 sg13g2_decap_8 FILLER_63_1759 ();
 sg13g2_fill_2 FILLER_63_1766 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_4 FILLER_64_112 ();
 sg13g2_fill_2 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_136 ();
 sg13g2_decap_8 FILLER_64_143 ();
 sg13g2_decap_8 FILLER_64_150 ();
 sg13g2_decap_4 FILLER_64_157 ();
 sg13g2_fill_2 FILLER_64_161 ();
 sg13g2_fill_2 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_decap_8 FILLER_64_205 ();
 sg13g2_decap_4 FILLER_64_212 ();
 sg13g2_fill_2 FILLER_64_216 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_243 ();
 sg13g2_fill_2 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_fill_2 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_297 ();
 sg13g2_fill_2 FILLER_64_307 ();
 sg13g2_fill_1 FILLER_64_309 ();
 sg13g2_decap_4 FILLER_64_318 ();
 sg13g2_decap_8 FILLER_64_326 ();
 sg13g2_decap_8 FILLER_64_333 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_347 ();
 sg13g2_decap_4 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_8 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_395 ();
 sg13g2_fill_1 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_64_432 ();
 sg13g2_fill_2 FILLER_64_439 ();
 sg13g2_fill_1 FILLER_64_441 ();
 sg13g2_decap_4 FILLER_64_454 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_decap_8 FILLER_64_473 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_decap_8 FILLER_64_487 ();
 sg13g2_decap_4 FILLER_64_494 ();
 sg13g2_fill_1 FILLER_64_498 ();
 sg13g2_decap_4 FILLER_64_510 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_532 ();
 sg13g2_decap_8 FILLER_64_539 ();
 sg13g2_fill_1 FILLER_64_546 ();
 sg13g2_decap_8 FILLER_64_574 ();
 sg13g2_decap_8 FILLER_64_581 ();
 sg13g2_decap_8 FILLER_64_588 ();
 sg13g2_decap_8 FILLER_64_595 ();
 sg13g2_decap_8 FILLER_64_602 ();
 sg13g2_fill_1 FILLER_64_609 ();
 sg13g2_fill_1 FILLER_64_623 ();
 sg13g2_decap_8 FILLER_64_634 ();
 sg13g2_decap_8 FILLER_64_641 ();
 sg13g2_decap_8 FILLER_64_648 ();
 sg13g2_decap_4 FILLER_64_655 ();
 sg13g2_fill_1 FILLER_64_659 ();
 sg13g2_decap_8 FILLER_64_695 ();
 sg13g2_decap_8 FILLER_64_702 ();
 sg13g2_fill_2 FILLER_64_709 ();
 sg13g2_fill_1 FILLER_64_711 ();
 sg13g2_fill_1 FILLER_64_740 ();
 sg13g2_decap_8 FILLER_64_768 ();
 sg13g2_fill_1 FILLER_64_775 ();
 sg13g2_decap_8 FILLER_64_784 ();
 sg13g2_decap_8 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_798 ();
 sg13g2_decap_4 FILLER_64_805 ();
 sg13g2_fill_2 FILLER_64_809 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_fill_2 FILLER_64_843 ();
 sg13g2_fill_1 FILLER_64_845 ();
 sg13g2_decap_8 FILLER_64_854 ();
 sg13g2_decap_8 FILLER_64_861 ();
 sg13g2_decap_8 FILLER_64_868 ();
 sg13g2_decap_4 FILLER_64_875 ();
 sg13g2_fill_2 FILLER_64_879 ();
 sg13g2_decap_8 FILLER_64_896 ();
 sg13g2_decap_8 FILLER_64_903 ();
 sg13g2_decap_8 FILLER_64_910 ();
 sg13g2_decap_8 FILLER_64_917 ();
 sg13g2_decap_8 FILLER_64_924 ();
 sg13g2_decap_8 FILLER_64_931 ();
 sg13g2_decap_8 FILLER_64_938 ();
 sg13g2_decap_8 FILLER_64_945 ();
 sg13g2_decap_4 FILLER_64_952 ();
 sg13g2_fill_1 FILLER_64_956 ();
 sg13g2_fill_1 FILLER_64_962 ();
 sg13g2_decap_8 FILLER_64_977 ();
 sg13g2_decap_8 FILLER_64_984 ();
 sg13g2_decap_8 FILLER_64_991 ();
 sg13g2_decap_8 FILLER_64_998 ();
 sg13g2_decap_8 FILLER_64_1005 ();
 sg13g2_fill_2 FILLER_64_1012 ();
 sg13g2_decap_8 FILLER_64_1027 ();
 sg13g2_decap_8 FILLER_64_1034 ();
 sg13g2_decap_4 FILLER_64_1041 ();
 sg13g2_fill_1 FILLER_64_1045 ();
 sg13g2_decap_8 FILLER_64_1054 ();
 sg13g2_decap_8 FILLER_64_1061 ();
 sg13g2_decap_4 FILLER_64_1068 ();
 sg13g2_fill_2 FILLER_64_1072 ();
 sg13g2_decap_8 FILLER_64_1082 ();
 sg13g2_decap_8 FILLER_64_1089 ();
 sg13g2_decap_8 FILLER_64_1096 ();
 sg13g2_decap_8 FILLER_64_1103 ();
 sg13g2_decap_8 FILLER_64_1110 ();
 sg13g2_decap_4 FILLER_64_1117 ();
 sg13g2_fill_1 FILLER_64_1121 ();
 sg13g2_decap_8 FILLER_64_1154 ();
 sg13g2_decap_8 FILLER_64_1161 ();
 sg13g2_decap_8 FILLER_64_1168 ();
 sg13g2_decap_8 FILLER_64_1175 ();
 sg13g2_fill_1 FILLER_64_1182 ();
 sg13g2_fill_2 FILLER_64_1188 ();
 sg13g2_fill_1 FILLER_64_1190 ();
 sg13g2_decap_8 FILLER_64_1196 ();
 sg13g2_decap_8 FILLER_64_1203 ();
 sg13g2_decap_8 FILLER_64_1210 ();
 sg13g2_fill_2 FILLER_64_1217 ();
 sg13g2_decap_4 FILLER_64_1232 ();
 sg13g2_fill_2 FILLER_64_1236 ();
 sg13g2_decap_8 FILLER_64_1244 ();
 sg13g2_decap_8 FILLER_64_1251 ();
 sg13g2_decap_8 FILLER_64_1258 ();
 sg13g2_decap_8 FILLER_64_1265 ();
 sg13g2_decap_8 FILLER_64_1272 ();
 sg13g2_decap_8 FILLER_64_1279 ();
 sg13g2_decap_8 FILLER_64_1286 ();
 sg13g2_fill_2 FILLER_64_1293 ();
 sg13g2_fill_1 FILLER_64_1298 ();
 sg13g2_decap_8 FILLER_64_1307 ();
 sg13g2_decap_8 FILLER_64_1314 ();
 sg13g2_decap_8 FILLER_64_1321 ();
 sg13g2_fill_1 FILLER_64_1328 ();
 sg13g2_decap_8 FILLER_64_1337 ();
 sg13g2_decap_8 FILLER_64_1344 ();
 sg13g2_decap_8 FILLER_64_1351 ();
 sg13g2_decap_8 FILLER_64_1358 ();
 sg13g2_decap_8 FILLER_64_1365 ();
 sg13g2_decap_8 FILLER_64_1388 ();
 sg13g2_decap_8 FILLER_64_1395 ();
 sg13g2_decap_8 FILLER_64_1402 ();
 sg13g2_decap_4 FILLER_64_1409 ();
 sg13g2_fill_2 FILLER_64_1413 ();
 sg13g2_fill_2 FILLER_64_1423 ();
 sg13g2_fill_1 FILLER_64_1425 ();
 sg13g2_decap_8 FILLER_64_1452 ();
 sg13g2_decap_8 FILLER_64_1459 ();
 sg13g2_decap_8 FILLER_64_1466 ();
 sg13g2_decap_8 FILLER_64_1473 ();
 sg13g2_decap_8 FILLER_64_1480 ();
 sg13g2_fill_2 FILLER_64_1487 ();
 sg13g2_fill_1 FILLER_64_1489 ();
 sg13g2_decap_8 FILLER_64_1498 ();
 sg13g2_fill_1 FILLER_64_1505 ();
 sg13g2_fill_2 FILLER_64_1516 ();
 sg13g2_fill_1 FILLER_64_1518 ();
 sg13g2_decap_8 FILLER_64_1530 ();
 sg13g2_decap_8 FILLER_64_1537 ();
 sg13g2_decap_8 FILLER_64_1544 ();
 sg13g2_fill_1 FILLER_64_1551 ();
 sg13g2_fill_2 FILLER_64_1560 ();
 sg13g2_decap_8 FILLER_64_1580 ();
 sg13g2_decap_8 FILLER_64_1587 ();
 sg13g2_fill_2 FILLER_64_1594 ();
 sg13g2_fill_1 FILLER_64_1596 ();
 sg13g2_decap_8 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1633 ();
 sg13g2_decap_4 FILLER_64_1640 ();
 sg13g2_fill_1 FILLER_64_1644 ();
 sg13g2_decap_8 FILLER_64_1661 ();
 sg13g2_decap_8 FILLER_64_1668 ();
 sg13g2_decap_8 FILLER_64_1675 ();
 sg13g2_decap_8 FILLER_64_1682 ();
 sg13g2_decap_8 FILLER_64_1689 ();
 sg13g2_decap_8 FILLER_64_1696 ();
 sg13g2_decap_8 FILLER_64_1703 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1717 ();
 sg13g2_decap_8 FILLER_64_1724 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_decap_8 FILLER_64_1738 ();
 sg13g2_decap_8 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_8 FILLER_64_1759 ();
 sg13g2_fill_2 FILLER_64_1766 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_4 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_46 ();
 sg13g2_decap_8 FILLER_65_62 ();
 sg13g2_decap_8 FILLER_65_69 ();
 sg13g2_decap_8 FILLER_65_76 ();
 sg13g2_decap_8 FILLER_65_83 ();
 sg13g2_decap_8 FILLER_65_90 ();
 sg13g2_decap_8 FILLER_65_97 ();
 sg13g2_decap_8 FILLER_65_104 ();
 sg13g2_decap_4 FILLER_65_111 ();
 sg13g2_fill_1 FILLER_65_115 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_fill_2 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_166 ();
 sg13g2_decap_8 FILLER_65_173 ();
 sg13g2_decap_8 FILLER_65_180 ();
 sg13g2_decap_8 FILLER_65_187 ();
 sg13g2_decap_8 FILLER_65_194 ();
 sg13g2_decap_8 FILLER_65_201 ();
 sg13g2_decap_8 FILLER_65_208 ();
 sg13g2_decap_8 FILLER_65_215 ();
 sg13g2_decap_8 FILLER_65_222 ();
 sg13g2_decap_8 FILLER_65_229 ();
 sg13g2_decap_8 FILLER_65_236 ();
 sg13g2_decap_8 FILLER_65_243 ();
 sg13g2_decap_8 FILLER_65_250 ();
 sg13g2_decap_8 FILLER_65_257 ();
 sg13g2_decap_8 FILLER_65_264 ();
 sg13g2_decap_8 FILLER_65_271 ();
 sg13g2_decap_8 FILLER_65_278 ();
 sg13g2_fill_2 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_297 ();
 sg13g2_decap_8 FILLER_65_304 ();
 sg13g2_decap_8 FILLER_65_311 ();
 sg13g2_decap_4 FILLER_65_318 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_decap_8 FILLER_65_341 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_fill_2 FILLER_65_389 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_402 ();
 sg13g2_decap_8 FILLER_65_416 ();
 sg13g2_decap_8 FILLER_65_423 ();
 sg13g2_decap_8 FILLER_65_430 ();
 sg13g2_decap_8 FILLER_65_437 ();
 sg13g2_decap_8 FILLER_65_444 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_8 FILLER_65_490 ();
 sg13g2_decap_8 FILLER_65_497 ();
 sg13g2_decap_8 FILLER_65_504 ();
 sg13g2_decap_8 FILLER_65_511 ();
 sg13g2_decap_8 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_fill_2 FILLER_65_546 ();
 sg13g2_decap_8 FILLER_65_572 ();
 sg13g2_decap_8 FILLER_65_579 ();
 sg13g2_decap_8 FILLER_65_586 ();
 sg13g2_decap_8 FILLER_65_593 ();
 sg13g2_decap_8 FILLER_65_600 ();
 sg13g2_decap_8 FILLER_65_639 ();
 sg13g2_decap_8 FILLER_65_646 ();
 sg13g2_decap_8 FILLER_65_653 ();
 sg13g2_decap_8 FILLER_65_660 ();
 sg13g2_fill_2 FILLER_65_667 ();
 sg13g2_fill_1 FILLER_65_669 ();
 sg13g2_decap_4 FILLER_65_679 ();
 sg13g2_decap_8 FILLER_65_691 ();
 sg13g2_decap_8 FILLER_65_698 ();
 sg13g2_decap_8 FILLER_65_705 ();
 sg13g2_decap_8 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_719 ();
 sg13g2_fill_2 FILLER_65_726 ();
 sg13g2_fill_1 FILLER_65_728 ();
 sg13g2_fill_1 FILLER_65_737 ();
 sg13g2_decap_8 FILLER_65_752 ();
 sg13g2_decap_4 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_773 ();
 sg13g2_decap_8 FILLER_65_780 ();
 sg13g2_decap_8 FILLER_65_787 ();
 sg13g2_decap_8 FILLER_65_794 ();
 sg13g2_decap_8 FILLER_65_801 ();
 sg13g2_fill_2 FILLER_65_808 ();
 sg13g2_fill_1 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_4 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_834 ();
 sg13g2_decap_8 FILLER_65_841 ();
 sg13g2_decap_4 FILLER_65_848 ();
 sg13g2_fill_2 FILLER_65_852 ();
 sg13g2_decap_8 FILLER_65_859 ();
 sg13g2_decap_8 FILLER_65_866 ();
 sg13g2_decap_8 FILLER_65_873 ();
 sg13g2_decap_8 FILLER_65_880 ();
 sg13g2_fill_2 FILLER_65_887 ();
 sg13g2_fill_1 FILLER_65_889 ();
 sg13g2_decap_8 FILLER_65_898 ();
 sg13g2_decap_8 FILLER_65_905 ();
 sg13g2_decap_8 FILLER_65_912 ();
 sg13g2_fill_1 FILLER_65_919 ();
 sg13g2_decap_8 FILLER_65_933 ();
 sg13g2_decap_8 FILLER_65_940 ();
 sg13g2_decap_8 FILLER_65_947 ();
 sg13g2_decap_8 FILLER_65_954 ();
 sg13g2_fill_2 FILLER_65_961 ();
 sg13g2_decap_8 FILLER_65_973 ();
 sg13g2_decap_8 FILLER_65_980 ();
 sg13g2_decap_8 FILLER_65_987 ();
 sg13g2_decap_8 FILLER_65_994 ();
 sg13g2_decap_8 FILLER_65_1001 ();
 sg13g2_decap_8 FILLER_65_1008 ();
 sg13g2_decap_8 FILLER_65_1015 ();
 sg13g2_decap_8 FILLER_65_1022 ();
 sg13g2_decap_4 FILLER_65_1042 ();
 sg13g2_fill_2 FILLER_65_1046 ();
 sg13g2_decap_8 FILLER_65_1056 ();
 sg13g2_decap_8 FILLER_65_1063 ();
 sg13g2_fill_2 FILLER_65_1070 ();
 sg13g2_fill_1 FILLER_65_1072 ();
 sg13g2_decap_8 FILLER_65_1085 ();
 sg13g2_decap_8 FILLER_65_1092 ();
 sg13g2_decap_8 FILLER_65_1099 ();
 sg13g2_decap_8 FILLER_65_1106 ();
 sg13g2_decap_8 FILLER_65_1113 ();
 sg13g2_decap_8 FILLER_65_1120 ();
 sg13g2_decap_8 FILLER_65_1127 ();
 sg13g2_decap_8 FILLER_65_1134 ();
 sg13g2_decap_8 FILLER_65_1141 ();
 sg13g2_fill_1 FILLER_65_1163 ();
 sg13g2_decap_8 FILLER_65_1172 ();
 sg13g2_decap_8 FILLER_65_1197 ();
 sg13g2_decap_8 FILLER_65_1204 ();
 sg13g2_decap_8 FILLER_65_1211 ();
 sg13g2_decap_8 FILLER_65_1218 ();
 sg13g2_decap_8 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1240 ();
 sg13g2_decap_8 FILLER_65_1247 ();
 sg13g2_fill_2 FILLER_65_1254 ();
 sg13g2_fill_1 FILLER_65_1256 ();
 sg13g2_decap_8 FILLER_65_1271 ();
 sg13g2_decap_8 FILLER_65_1278 ();
 sg13g2_decap_8 FILLER_65_1285 ();
 sg13g2_fill_2 FILLER_65_1292 ();
 sg13g2_fill_1 FILLER_65_1294 ();
 sg13g2_fill_2 FILLER_65_1300 ();
 sg13g2_fill_1 FILLER_65_1302 ();
 sg13g2_decap_8 FILLER_65_1331 ();
 sg13g2_decap_8 FILLER_65_1338 ();
 sg13g2_decap_8 FILLER_65_1345 ();
 sg13g2_decap_8 FILLER_65_1352 ();
 sg13g2_fill_2 FILLER_65_1359 ();
 sg13g2_fill_2 FILLER_65_1375 ();
 sg13g2_decap_8 FILLER_65_1384 ();
 sg13g2_decap_8 FILLER_65_1391 ();
 sg13g2_decap_8 FILLER_65_1398 ();
 sg13g2_fill_2 FILLER_65_1405 ();
 sg13g2_fill_1 FILLER_65_1407 ();
 sg13g2_decap_4 FILLER_65_1416 ();
 sg13g2_decap_8 FILLER_65_1430 ();
 sg13g2_fill_2 FILLER_65_1437 ();
 sg13g2_decap_8 FILLER_65_1448 ();
 sg13g2_decap_8 FILLER_65_1455 ();
 sg13g2_decap_8 FILLER_65_1462 ();
 sg13g2_decap_8 FILLER_65_1469 ();
 sg13g2_fill_1 FILLER_65_1476 ();
 sg13g2_decap_8 FILLER_65_1481 ();
 sg13g2_fill_1 FILLER_65_1488 ();
 sg13g2_decap_8 FILLER_65_1509 ();
 sg13g2_decap_8 FILLER_65_1516 ();
 sg13g2_decap_8 FILLER_65_1523 ();
 sg13g2_decap_8 FILLER_65_1530 ();
 sg13g2_fill_2 FILLER_65_1537 ();
 sg13g2_decap_4 FILLER_65_1547 ();
 sg13g2_fill_2 FILLER_65_1558 ();
 sg13g2_decap_8 FILLER_65_1575 ();
 sg13g2_decap_8 FILLER_65_1582 ();
 sg13g2_decap_8 FILLER_65_1589 ();
 sg13g2_decap_8 FILLER_65_1596 ();
 sg13g2_decap_8 FILLER_65_1603 ();
 sg13g2_decap_8 FILLER_65_1616 ();
 sg13g2_decap_8 FILLER_65_1623 ();
 sg13g2_decap_8 FILLER_65_1630 ();
 sg13g2_decap_8 FILLER_65_1637 ();
 sg13g2_decap_4 FILLER_65_1644 ();
 sg13g2_decap_8 FILLER_65_1651 ();
 sg13g2_decap_8 FILLER_65_1658 ();
 sg13g2_decap_8 FILLER_65_1665 ();
 sg13g2_decap_8 FILLER_65_1672 ();
 sg13g2_decap_8 FILLER_65_1679 ();
 sg13g2_decap_8 FILLER_65_1686 ();
 sg13g2_decap_8 FILLER_65_1693 ();
 sg13g2_decap_8 FILLER_65_1700 ();
 sg13g2_decap_8 FILLER_65_1707 ();
 sg13g2_decap_8 FILLER_65_1714 ();
 sg13g2_decap_8 FILLER_65_1721 ();
 sg13g2_decap_8 FILLER_65_1728 ();
 sg13g2_decap_8 FILLER_65_1735 ();
 sg13g2_decap_8 FILLER_65_1742 ();
 sg13g2_decap_8 FILLER_65_1749 ();
 sg13g2_decap_8 FILLER_65_1756 ();
 sg13g2_decap_4 FILLER_65_1763 ();
 sg13g2_fill_1 FILLER_65_1767 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_4 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_46 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_4 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_132 ();
 sg13g2_decap_8 FILLER_66_139 ();
 sg13g2_decap_4 FILLER_66_146 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_decap_8 FILLER_66_164 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_decap_8 FILLER_66_178 ();
 sg13g2_decap_8 FILLER_66_185 ();
 sg13g2_fill_2 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_194 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_fill_1 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_decap_4 FILLER_66_349 ();
 sg13g2_fill_1 FILLER_66_353 ();
 sg13g2_decap_8 FILLER_66_372 ();
 sg13g2_decap_8 FILLER_66_379 ();
 sg13g2_decap_4 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_4 FILLER_66_420 ();
 sg13g2_fill_2 FILLER_66_424 ();
 sg13g2_decap_8 FILLER_66_434 ();
 sg13g2_decap_8 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_448 ();
 sg13g2_decap_4 FILLER_66_455 ();
 sg13g2_fill_2 FILLER_66_459 ();
 sg13g2_decap_8 FILLER_66_471 ();
 sg13g2_decap_8 FILLER_66_484 ();
 sg13g2_decap_8 FILLER_66_491 ();
 sg13g2_decap_8 FILLER_66_498 ();
 sg13g2_decap_4 FILLER_66_505 ();
 sg13g2_fill_1 FILLER_66_509 ();
 sg13g2_decap_8 FILLER_66_534 ();
 sg13g2_decap_8 FILLER_66_541 ();
 sg13g2_decap_8 FILLER_66_548 ();
 sg13g2_fill_2 FILLER_66_555 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_decap_8 FILLER_66_570 ();
 sg13g2_decap_8 FILLER_66_577 ();
 sg13g2_decap_8 FILLER_66_584 ();
 sg13g2_decap_8 FILLER_66_591 ();
 sg13g2_decap_8 FILLER_66_598 ();
 sg13g2_decap_4 FILLER_66_605 ();
 sg13g2_fill_1 FILLER_66_609 ();
 sg13g2_fill_2 FILLER_66_618 ();
 sg13g2_fill_2 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_638 ();
 sg13g2_decap_8 FILLER_66_645 ();
 sg13g2_decap_8 FILLER_66_652 ();
 sg13g2_decap_8 FILLER_66_659 ();
 sg13g2_decap_8 FILLER_66_666 ();
 sg13g2_decap_8 FILLER_66_673 ();
 sg13g2_decap_8 FILLER_66_680 ();
 sg13g2_decap_8 FILLER_66_690 ();
 sg13g2_decap_8 FILLER_66_697 ();
 sg13g2_decap_8 FILLER_66_704 ();
 sg13g2_decap_8 FILLER_66_711 ();
 sg13g2_decap_4 FILLER_66_718 ();
 sg13g2_fill_1 FILLER_66_722 ();
 sg13g2_decap_4 FILLER_66_731 ();
 sg13g2_fill_1 FILLER_66_735 ();
 sg13g2_fill_2 FILLER_66_747 ();
 sg13g2_decap_8 FILLER_66_757 ();
 sg13g2_decap_8 FILLER_66_764 ();
 sg13g2_decap_8 FILLER_66_771 ();
 sg13g2_decap_8 FILLER_66_778 ();
 sg13g2_decap_8 FILLER_66_785 ();
 sg13g2_decap_4 FILLER_66_792 ();
 sg13g2_fill_1 FILLER_66_796 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_8 FILLER_66_856 ();
 sg13g2_decap_4 FILLER_66_863 ();
 sg13g2_fill_1 FILLER_66_867 ();
 sg13g2_decap_8 FILLER_66_900 ();
 sg13g2_decap_8 FILLER_66_907 ();
 sg13g2_decap_8 FILLER_66_914 ();
 sg13g2_decap_8 FILLER_66_921 ();
 sg13g2_fill_2 FILLER_66_928 ();
 sg13g2_fill_2 FILLER_66_936 ();
 sg13g2_fill_1 FILLER_66_938 ();
 sg13g2_fill_2 FILLER_66_947 ();
 sg13g2_decap_4 FILLER_66_957 ();
 sg13g2_fill_2 FILLER_66_961 ();
 sg13g2_decap_8 FILLER_66_985 ();
 sg13g2_decap_4 FILLER_66_992 ();
 sg13g2_decap_8 FILLER_66_1004 ();
 sg13g2_decap_8 FILLER_66_1011 ();
 sg13g2_decap_8 FILLER_66_1018 ();
 sg13g2_decap_8 FILLER_66_1025 ();
 sg13g2_decap_8 FILLER_66_1032 ();
 sg13g2_decap_4 FILLER_66_1039 ();
 sg13g2_fill_1 FILLER_66_1043 ();
 sg13g2_decap_8 FILLER_66_1060 ();
 sg13g2_decap_8 FILLER_66_1067 ();
 sg13g2_decap_8 FILLER_66_1074 ();
 sg13g2_decap_8 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1102 ();
 sg13g2_fill_2 FILLER_66_1109 ();
 sg13g2_decap_8 FILLER_66_1119 ();
 sg13g2_fill_2 FILLER_66_1126 ();
 sg13g2_fill_1 FILLER_66_1128 ();
 sg13g2_decap_8 FILLER_66_1137 ();
 sg13g2_decap_8 FILLER_66_1144 ();
 sg13g2_decap_4 FILLER_66_1151 ();
 sg13g2_fill_2 FILLER_66_1155 ();
 sg13g2_decap_4 FILLER_66_1162 ();
 sg13g2_fill_2 FILLER_66_1166 ();
 sg13g2_decap_8 FILLER_66_1176 ();
 sg13g2_decap_8 FILLER_66_1183 ();
 sg13g2_decap_8 FILLER_66_1190 ();
 sg13g2_decap_8 FILLER_66_1197 ();
 sg13g2_decap_4 FILLER_66_1204 ();
 sg13g2_fill_2 FILLER_66_1208 ();
 sg13g2_decap_8 FILLER_66_1231 ();
 sg13g2_decap_8 FILLER_66_1238 ();
 sg13g2_decap_8 FILLER_66_1245 ();
 sg13g2_fill_2 FILLER_66_1256 ();
 sg13g2_fill_1 FILLER_66_1258 ();
 sg13g2_decap_8 FILLER_66_1271 ();
 sg13g2_decap_4 FILLER_66_1278 ();
 sg13g2_fill_2 FILLER_66_1282 ();
 sg13g2_fill_2 FILLER_66_1289 ();
 sg13g2_decap_8 FILLER_66_1299 ();
 sg13g2_decap_8 FILLER_66_1306 ();
 sg13g2_decap_8 FILLER_66_1313 ();
 sg13g2_decap_8 FILLER_66_1320 ();
 sg13g2_decap_8 FILLER_66_1327 ();
 sg13g2_fill_2 FILLER_66_1334 ();
 sg13g2_fill_1 FILLER_66_1336 ();
 sg13g2_decap_8 FILLER_66_1342 ();
 sg13g2_decap_4 FILLER_66_1349 ();
 sg13g2_decap_8 FILLER_66_1361 ();
 sg13g2_fill_1 FILLER_66_1368 ();
 sg13g2_decap_8 FILLER_66_1385 ();
 sg13g2_decap_8 FILLER_66_1392 ();
 sg13g2_decap_4 FILLER_66_1399 ();
 sg13g2_fill_2 FILLER_66_1403 ();
 sg13g2_fill_2 FILLER_66_1413 ();
 sg13g2_decap_8 FILLER_66_1420 ();
 sg13g2_decap_8 FILLER_66_1427 ();
 sg13g2_decap_8 FILLER_66_1434 ();
 sg13g2_decap_8 FILLER_66_1441 ();
 sg13g2_decap_8 FILLER_66_1448 ();
 sg13g2_decap_8 FILLER_66_1460 ();
 sg13g2_decap_8 FILLER_66_1467 ();
 sg13g2_decap_8 FILLER_66_1474 ();
 sg13g2_decap_8 FILLER_66_1481 ();
 sg13g2_fill_2 FILLER_66_1488 ();
 sg13g2_fill_1 FILLER_66_1490 ();
 sg13g2_decap_8 FILLER_66_1502 ();
 sg13g2_decap_8 FILLER_66_1509 ();
 sg13g2_decap_8 FILLER_66_1516 ();
 sg13g2_decap_8 FILLER_66_1523 ();
 sg13g2_decap_8 FILLER_66_1530 ();
 sg13g2_decap_8 FILLER_66_1537 ();
 sg13g2_decap_8 FILLER_66_1544 ();
 sg13g2_fill_1 FILLER_66_1551 ();
 sg13g2_decap_4 FILLER_66_1557 ();
 sg13g2_decap_8 FILLER_66_1574 ();
 sg13g2_decap_8 FILLER_66_1581 ();
 sg13g2_decap_8 FILLER_66_1588 ();
 sg13g2_decap_8 FILLER_66_1595 ();
 sg13g2_decap_8 FILLER_66_1602 ();
 sg13g2_decap_8 FILLER_66_1609 ();
 sg13g2_decap_4 FILLER_66_1616 ();
 sg13g2_decap_8 FILLER_66_1646 ();
 sg13g2_decap_8 FILLER_66_1653 ();
 sg13g2_decap_8 FILLER_66_1660 ();
 sg13g2_decap_4 FILLER_66_1671 ();
 sg13g2_decap_8 FILLER_66_1700 ();
 sg13g2_decap_8 FILLER_66_1707 ();
 sg13g2_decap_8 FILLER_66_1714 ();
 sg13g2_decap_8 FILLER_66_1721 ();
 sg13g2_decap_8 FILLER_66_1728 ();
 sg13g2_decap_8 FILLER_66_1735 ();
 sg13g2_decap_8 FILLER_66_1742 ();
 sg13g2_decap_8 FILLER_66_1749 ();
 sg13g2_decap_8 FILLER_66_1756 ();
 sg13g2_decap_4 FILLER_66_1763 ();
 sg13g2_fill_1 FILLER_66_1767 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_28 ();
 sg13g2_fill_1 FILLER_67_30 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_46 ();
 sg13g2_decap_8 FILLER_67_53 ();
 sg13g2_decap_8 FILLER_67_60 ();
 sg13g2_decap_4 FILLER_67_67 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_fill_2 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_4 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_decap_8 FILLER_67_170 ();
 sg13g2_decap_4 FILLER_67_177 ();
 sg13g2_fill_1 FILLER_67_206 ();
 sg13g2_decap_8 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_219 ();
 sg13g2_decap_8 FILLER_67_226 ();
 sg13g2_decap_8 FILLER_67_233 ();
 sg13g2_decap_4 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_decap_8 FILLER_67_281 ();
 sg13g2_decap_8 FILLER_67_288 ();
 sg13g2_decap_4 FILLER_67_295 ();
 sg13g2_decap_8 FILLER_67_307 ();
 sg13g2_decap_8 FILLER_67_314 ();
 sg13g2_decap_8 FILLER_67_321 ();
 sg13g2_decap_8 FILLER_67_328 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_decap_4 FILLER_67_350 ();
 sg13g2_fill_1 FILLER_67_354 ();
 sg13g2_decap_8 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_decap_8 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_67_415 ();
 sg13g2_decap_4 FILLER_67_422 ();
 sg13g2_fill_2 FILLER_67_426 ();
 sg13g2_decap_8 FILLER_67_433 ();
 sg13g2_decap_8 FILLER_67_440 ();
 sg13g2_decap_8 FILLER_67_447 ();
 sg13g2_fill_2 FILLER_67_466 ();
 sg13g2_decap_8 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_fill_2 FILLER_67_511 ();
 sg13g2_fill_1 FILLER_67_513 ();
 sg13g2_decap_4 FILLER_67_519 ();
 sg13g2_decap_8 FILLER_67_537 ();
 sg13g2_decap_8 FILLER_67_544 ();
 sg13g2_decap_4 FILLER_67_551 ();
 sg13g2_decap_8 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_4 FILLER_67_609 ();
 sg13g2_fill_2 FILLER_67_613 ();
 sg13g2_decap_8 FILLER_67_635 ();
 sg13g2_decap_8 FILLER_67_642 ();
 sg13g2_decap_8 FILLER_67_649 ();
 sg13g2_decap_8 FILLER_67_656 ();
 sg13g2_decap_8 FILLER_67_663 ();
 sg13g2_decap_4 FILLER_67_670 ();
 sg13g2_fill_2 FILLER_67_674 ();
 sg13g2_fill_1 FILLER_67_680 ();
 sg13g2_decap_8 FILLER_67_694 ();
 sg13g2_decap_8 FILLER_67_701 ();
 sg13g2_decap_8 FILLER_67_708 ();
 sg13g2_decap_8 FILLER_67_715 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_fill_2 FILLER_67_770 ();
 sg13g2_fill_1 FILLER_67_772 ();
 sg13g2_decap_8 FILLER_67_786 ();
 sg13g2_decap_8 FILLER_67_793 ();
 sg13g2_decap_8 FILLER_67_800 ();
 sg13g2_decap_4 FILLER_67_807 ();
 sg13g2_fill_1 FILLER_67_811 ();
 sg13g2_decap_8 FILLER_67_816 ();
 sg13g2_decap_8 FILLER_67_823 ();
 sg13g2_decap_8 FILLER_67_830 ();
 sg13g2_decap_8 FILLER_67_837 ();
 sg13g2_decap_8 FILLER_67_844 ();
 sg13g2_decap_8 FILLER_67_851 ();
 sg13g2_decap_8 FILLER_67_858 ();
 sg13g2_decap_8 FILLER_67_865 ();
 sg13g2_fill_2 FILLER_67_872 ();
 sg13g2_decap_8 FILLER_67_885 ();
 sg13g2_decap_8 FILLER_67_892 ();
 sg13g2_decap_8 FILLER_67_899 ();
 sg13g2_decap_8 FILLER_67_906 ();
 sg13g2_decap_8 FILLER_67_913 ();
 sg13g2_decap_8 FILLER_67_920 ();
 sg13g2_fill_2 FILLER_67_927 ();
 sg13g2_fill_1 FILLER_67_929 ();
 sg13g2_fill_2 FILLER_67_947 ();
 sg13g2_decap_8 FILLER_67_965 ();
 sg13g2_decap_8 FILLER_67_972 ();
 sg13g2_decap_8 FILLER_67_979 ();
 sg13g2_fill_2 FILLER_67_986 ();
 sg13g2_decap_8 FILLER_67_994 ();
 sg13g2_decap_8 FILLER_67_1001 ();
 sg13g2_fill_2 FILLER_67_1008 ();
 sg13g2_fill_1 FILLER_67_1010 ();
 sg13g2_decap_8 FILLER_67_1019 ();
 sg13g2_decap_8 FILLER_67_1026 ();
 sg13g2_decap_8 FILLER_67_1033 ();
 sg13g2_fill_2 FILLER_67_1040 ();
 sg13g2_decap_8 FILLER_67_1050 ();
 sg13g2_decap_4 FILLER_67_1057 ();
 sg13g2_fill_1 FILLER_67_1061 ();
 sg13g2_decap_4 FILLER_67_1070 ();
 sg13g2_fill_2 FILLER_67_1074 ();
 sg13g2_decap_8 FILLER_67_1092 ();
 sg13g2_decap_8 FILLER_67_1099 ();
 sg13g2_decap_8 FILLER_67_1106 ();
 sg13g2_fill_2 FILLER_67_1113 ();
 sg13g2_decap_8 FILLER_67_1127 ();
 sg13g2_decap_8 FILLER_67_1134 ();
 sg13g2_decap_8 FILLER_67_1141 ();
 sg13g2_decap_8 FILLER_67_1148 ();
 sg13g2_decap_8 FILLER_67_1155 ();
 sg13g2_decap_8 FILLER_67_1162 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1176 ();
 sg13g2_fill_1 FILLER_67_1183 ();
 sg13g2_decap_8 FILLER_67_1188 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_fill_1 FILLER_67_1209 ();
 sg13g2_fill_1 FILLER_67_1220 ();
 sg13g2_fill_2 FILLER_67_1229 ();
 sg13g2_decap_8 FILLER_67_1240 ();
 sg13g2_decap_8 FILLER_67_1247 ();
 sg13g2_decap_4 FILLER_67_1254 ();
 sg13g2_fill_1 FILLER_67_1258 ();
 sg13g2_decap_8 FILLER_67_1268 ();
 sg13g2_decap_4 FILLER_67_1275 ();
 sg13g2_fill_1 FILLER_67_1279 ();
 sg13g2_decap_8 FILLER_67_1296 ();
 sg13g2_decap_4 FILLER_67_1303 ();
 sg13g2_decap_8 FILLER_67_1315 ();
 sg13g2_decap_4 FILLER_67_1322 ();
 sg13g2_fill_1 FILLER_67_1326 ();
 sg13g2_decap_8 FILLER_67_1341 ();
 sg13g2_decap_8 FILLER_67_1348 ();
 sg13g2_decap_8 FILLER_67_1355 ();
 sg13g2_decap_8 FILLER_67_1362 ();
 sg13g2_decap_8 FILLER_67_1369 ();
 sg13g2_decap_8 FILLER_67_1376 ();
 sg13g2_decap_4 FILLER_67_1383 ();
 sg13g2_decap_8 FILLER_67_1392 ();
 sg13g2_decap_8 FILLER_67_1399 ();
 sg13g2_decap_8 FILLER_67_1406 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_decap_8 FILLER_67_1420 ();
 sg13g2_decap_8 FILLER_67_1427 ();
 sg13g2_decap_8 FILLER_67_1434 ();
 sg13g2_decap_8 FILLER_67_1441 ();
 sg13g2_decap_4 FILLER_67_1448 ();
 sg13g2_decap_8 FILLER_67_1475 ();
 sg13g2_decap_4 FILLER_67_1482 ();
 sg13g2_fill_2 FILLER_67_1486 ();
 sg13g2_decap_8 FILLER_67_1500 ();
 sg13g2_decap_8 FILLER_67_1507 ();
 sg13g2_decap_8 FILLER_67_1514 ();
 sg13g2_decap_8 FILLER_67_1521 ();
 sg13g2_fill_1 FILLER_67_1528 ();
 sg13g2_decap_8 FILLER_67_1537 ();
 sg13g2_decap_8 FILLER_67_1544 ();
 sg13g2_decap_8 FILLER_67_1551 ();
 sg13g2_decap_8 FILLER_67_1558 ();
 sg13g2_decap_8 FILLER_67_1570 ();
 sg13g2_fill_1 FILLER_67_1577 ();
 sg13g2_decap_4 FILLER_67_1586 ();
 sg13g2_fill_1 FILLER_67_1590 ();
 sg13g2_decap_8 FILLER_67_1595 ();
 sg13g2_fill_1 FILLER_67_1602 ();
 sg13g2_decap_4 FILLER_67_1626 ();
 sg13g2_fill_1 FILLER_67_1630 ();
 sg13g2_fill_1 FILLER_67_1635 ();
 sg13g2_fill_2 FILLER_67_1654 ();
 sg13g2_decap_8 FILLER_67_1682 ();
 sg13g2_decap_8 FILLER_67_1689 ();
 sg13g2_decap_8 FILLER_67_1696 ();
 sg13g2_decap_8 FILLER_67_1703 ();
 sg13g2_decap_8 FILLER_67_1710 ();
 sg13g2_decap_8 FILLER_67_1717 ();
 sg13g2_decap_8 FILLER_67_1724 ();
 sg13g2_decap_8 FILLER_67_1731 ();
 sg13g2_decap_8 FILLER_67_1738 ();
 sg13g2_decap_8 FILLER_67_1745 ();
 sg13g2_decap_8 FILLER_67_1752 ();
 sg13g2_decap_8 FILLER_67_1759 ();
 sg13g2_fill_2 FILLER_67_1766 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_4 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_18 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_4 FILLER_68_91 ();
 sg13g2_fill_1 FILLER_68_95 ();
 sg13g2_fill_2 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_103 ();
 sg13g2_decap_8 FILLER_68_108 ();
 sg13g2_decap_8 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_122 ();
 sg13g2_fill_1 FILLER_68_124 ();
 sg13g2_decap_8 FILLER_68_138 ();
 sg13g2_decap_4 FILLER_68_145 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_4 FILLER_68_196 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_decap_8 FILLER_68_211 ();
 sg13g2_decap_8 FILLER_68_254 ();
 sg13g2_decap_4 FILLER_68_261 ();
 sg13g2_fill_1 FILLER_68_265 ();
 sg13g2_decap_8 FILLER_68_270 ();
 sg13g2_decap_8 FILLER_68_277 ();
 sg13g2_decap_4 FILLER_68_284 ();
 sg13g2_fill_1 FILLER_68_288 ();
 sg13g2_decap_8 FILLER_68_302 ();
 sg13g2_decap_8 FILLER_68_309 ();
 sg13g2_decap_8 FILLER_68_321 ();
 sg13g2_fill_2 FILLER_68_328 ();
 sg13g2_fill_2 FILLER_68_338 ();
 sg13g2_fill_1 FILLER_68_340 ();
 sg13g2_decap_8 FILLER_68_349 ();
 sg13g2_decap_4 FILLER_68_356 ();
 sg13g2_fill_2 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_4 FILLER_68_391 ();
 sg13g2_fill_2 FILLER_68_395 ();
 sg13g2_decap_8 FILLER_68_401 ();
 sg13g2_decap_8 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_68_415 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_decap_4 FILLER_68_439 ();
 sg13g2_fill_1 FILLER_68_443 ();
 sg13g2_decap_8 FILLER_68_452 ();
 sg13g2_decap_8 FILLER_68_459 ();
 sg13g2_decap_8 FILLER_68_478 ();
 sg13g2_decap_8 FILLER_68_485 ();
 sg13g2_decap_8 FILLER_68_492 ();
 sg13g2_decap_8 FILLER_68_499 ();
 sg13g2_decap_8 FILLER_68_506 ();
 sg13g2_decap_8 FILLER_68_513 ();
 sg13g2_decap_4 FILLER_68_520 ();
 sg13g2_fill_2 FILLER_68_524 ();
 sg13g2_decap_8 FILLER_68_545 ();
 sg13g2_decap_8 FILLER_68_552 ();
 sg13g2_decap_4 FILLER_68_559 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_decap_8 FILLER_68_577 ();
 sg13g2_decap_8 FILLER_68_584 ();
 sg13g2_decap_4 FILLER_68_591 ();
 sg13g2_fill_2 FILLER_68_595 ();
 sg13g2_decap_8 FILLER_68_605 ();
 sg13g2_decap_8 FILLER_68_612 ();
 sg13g2_fill_1 FILLER_68_619 ();
 sg13g2_decap_8 FILLER_68_631 ();
 sg13g2_decap_8 FILLER_68_638 ();
 sg13g2_decap_8 FILLER_68_645 ();
 sg13g2_decap_8 FILLER_68_652 ();
 sg13g2_decap_4 FILLER_68_659 ();
 sg13g2_fill_2 FILLER_68_663 ();
 sg13g2_fill_2 FILLER_68_691 ();
 sg13g2_decap_8 FILLER_68_706 ();
 sg13g2_decap_8 FILLER_68_713 ();
 sg13g2_decap_8 FILLER_68_720 ();
 sg13g2_decap_8 FILLER_68_727 ();
 sg13g2_decap_8 FILLER_68_734 ();
 sg13g2_decap_8 FILLER_68_741 ();
 sg13g2_decap_8 FILLER_68_748 ();
 sg13g2_decap_8 FILLER_68_755 ();
 sg13g2_decap_4 FILLER_68_762 ();
 sg13g2_fill_2 FILLER_68_766 ();
 sg13g2_fill_2 FILLER_68_781 ();
 sg13g2_fill_1 FILLER_68_783 ();
 sg13g2_decap_4 FILLER_68_795 ();
 sg13g2_fill_2 FILLER_68_799 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_4 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_849 ();
 sg13g2_decap_4 FILLER_68_856 ();
 sg13g2_decap_4 FILLER_68_873 ();
 sg13g2_fill_2 FILLER_68_877 ();
 sg13g2_decap_8 FILLER_68_891 ();
 sg13g2_decap_8 FILLER_68_898 ();
 sg13g2_decap_8 FILLER_68_905 ();
 sg13g2_decap_8 FILLER_68_912 ();
 sg13g2_decap_8 FILLER_68_919 ();
 sg13g2_decap_8 FILLER_68_926 ();
 sg13g2_decap_8 FILLER_68_933 ();
 sg13g2_decap_4 FILLER_68_940 ();
 sg13g2_fill_1 FILLER_68_944 ();
 sg13g2_fill_1 FILLER_68_950 ();
 sg13g2_fill_2 FILLER_68_963 ();
 sg13g2_fill_1 FILLER_68_965 ();
 sg13g2_decap_8 FILLER_68_972 ();
 sg13g2_decap_8 FILLER_68_979 ();
 sg13g2_fill_2 FILLER_68_986 ();
 sg13g2_decap_8 FILLER_68_1000 ();
 sg13g2_decap_4 FILLER_68_1007 ();
 sg13g2_fill_1 FILLER_68_1011 ();
 sg13g2_decap_8 FILLER_68_1016 ();
 sg13g2_fill_1 FILLER_68_1023 ();
 sg13g2_decap_8 FILLER_68_1032 ();
 sg13g2_decap_8 FILLER_68_1039 ();
 sg13g2_decap_8 FILLER_68_1046 ();
 sg13g2_decap_8 FILLER_68_1053 ();
 sg13g2_decap_8 FILLER_68_1060 ();
 sg13g2_fill_1 FILLER_68_1067 ();
 sg13g2_decap_8 FILLER_68_1073 ();
 sg13g2_decap_4 FILLER_68_1080 ();
 sg13g2_decap_8 FILLER_68_1087 ();
 sg13g2_decap_8 FILLER_68_1094 ();
 sg13g2_decap_8 FILLER_68_1101 ();
 sg13g2_fill_2 FILLER_68_1108 ();
 sg13g2_fill_1 FILLER_68_1110 ();
 sg13g2_decap_8 FILLER_68_1117 ();
 sg13g2_decap_8 FILLER_68_1124 ();
 sg13g2_decap_8 FILLER_68_1131 ();
 sg13g2_decap_8 FILLER_68_1138 ();
 sg13g2_decap_4 FILLER_68_1145 ();
 sg13g2_fill_2 FILLER_68_1149 ();
 sg13g2_decap_8 FILLER_68_1177 ();
 sg13g2_decap_8 FILLER_68_1184 ();
 sg13g2_decap_8 FILLER_68_1191 ();
 sg13g2_decap_8 FILLER_68_1198 ();
 sg13g2_decap_8 FILLER_68_1205 ();
 sg13g2_decap_8 FILLER_68_1212 ();
 sg13g2_decap_8 FILLER_68_1219 ();
 sg13g2_decap_8 FILLER_68_1226 ();
 sg13g2_decap_8 FILLER_68_1233 ();
 sg13g2_decap_8 FILLER_68_1240 ();
 sg13g2_decap_4 FILLER_68_1247 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_decap_8 FILLER_68_1258 ();
 sg13g2_decap_8 FILLER_68_1265 ();
 sg13g2_decap_8 FILLER_68_1272 ();
 sg13g2_decap_4 FILLER_68_1279 ();
 sg13g2_fill_2 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1318 ();
 sg13g2_decap_4 FILLER_68_1325 ();
 sg13g2_fill_2 FILLER_68_1329 ();
 sg13g2_decap_8 FILLER_68_1334 ();
 sg13g2_decap_8 FILLER_68_1341 ();
 sg13g2_decap_8 FILLER_68_1348 ();
 sg13g2_decap_8 FILLER_68_1355 ();
 sg13g2_fill_1 FILLER_68_1362 ();
 sg13g2_decap_8 FILLER_68_1403 ();
 sg13g2_decap_8 FILLER_68_1410 ();
 sg13g2_fill_1 FILLER_68_1417 ();
 sg13g2_decap_8 FILLER_68_1426 ();
 sg13g2_decap_8 FILLER_68_1433 ();
 sg13g2_decap_8 FILLER_68_1440 ();
 sg13g2_decap_8 FILLER_68_1447 ();
 sg13g2_fill_2 FILLER_68_1454 ();
 sg13g2_decap_8 FILLER_68_1461 ();
 sg13g2_decap_8 FILLER_68_1468 ();
 sg13g2_decap_8 FILLER_68_1475 ();
 sg13g2_decap_4 FILLER_68_1482 ();
 sg13g2_fill_2 FILLER_68_1486 ();
 sg13g2_decap_8 FILLER_68_1492 ();
 sg13g2_decap_8 FILLER_68_1499 ();
 sg13g2_fill_2 FILLER_68_1506 ();
 sg13g2_fill_1 FILLER_68_1512 ();
 sg13g2_decap_8 FILLER_68_1526 ();
 sg13g2_decap_8 FILLER_68_1533 ();
 sg13g2_decap_8 FILLER_68_1540 ();
 sg13g2_decap_8 FILLER_68_1547 ();
 sg13g2_decap_8 FILLER_68_1554 ();
 sg13g2_decap_8 FILLER_68_1561 ();
 sg13g2_decap_8 FILLER_68_1568 ();
 sg13g2_decap_8 FILLER_68_1579 ();
 sg13g2_decap_8 FILLER_68_1603 ();
 sg13g2_decap_8 FILLER_68_1610 ();
 sg13g2_decap_8 FILLER_68_1617 ();
 sg13g2_decap_8 FILLER_68_1624 ();
 sg13g2_decap_8 FILLER_68_1631 ();
 sg13g2_fill_1 FILLER_68_1638 ();
 sg13g2_decap_8 FILLER_68_1643 ();
 sg13g2_decap_4 FILLER_68_1650 ();
 sg13g2_fill_1 FILLER_68_1654 ();
 sg13g2_decap_8 FILLER_68_1668 ();
 sg13g2_decap_8 FILLER_68_1675 ();
 sg13g2_decap_8 FILLER_68_1682 ();
 sg13g2_decap_8 FILLER_68_1689 ();
 sg13g2_decap_8 FILLER_68_1696 ();
 sg13g2_decap_8 FILLER_68_1703 ();
 sg13g2_decap_8 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1717 ();
 sg13g2_decap_8 FILLER_68_1724 ();
 sg13g2_decap_8 FILLER_68_1731 ();
 sg13g2_decap_8 FILLER_68_1738 ();
 sg13g2_decap_8 FILLER_68_1745 ();
 sg13g2_decap_8 FILLER_68_1752 ();
 sg13g2_decap_8 FILLER_68_1759 ();
 sg13g2_fill_2 FILLER_68_1766 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_47 ();
 sg13g2_decap_8 FILLER_69_54 ();
 sg13g2_decap_8 FILLER_69_61 ();
 sg13g2_decap_8 FILLER_69_68 ();
 sg13g2_decap_4 FILLER_69_75 ();
 sg13g2_fill_2 FILLER_69_79 ();
 sg13g2_decap_8 FILLER_69_85 ();
 sg13g2_decap_8 FILLER_69_92 ();
 sg13g2_decap_8 FILLER_69_99 ();
 sg13g2_decap_8 FILLER_69_106 ();
 sg13g2_decap_8 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_decap_8 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_139 ();
 sg13g2_decap_8 FILLER_69_151 ();
 sg13g2_decap_8 FILLER_69_158 ();
 sg13g2_decap_8 FILLER_69_165 ();
 sg13g2_decap_8 FILLER_69_172 ();
 sg13g2_decap_8 FILLER_69_179 ();
 sg13g2_decap_8 FILLER_69_186 ();
 sg13g2_decap_8 FILLER_69_193 ();
 sg13g2_decap_4 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_209 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_243 ();
 sg13g2_decap_8 FILLER_69_250 ();
 sg13g2_decap_4 FILLER_69_257 ();
 sg13g2_decap_8 FILLER_69_274 ();
 sg13g2_decap_8 FILLER_69_281 ();
 sg13g2_fill_1 FILLER_69_288 ();
 sg13g2_decap_4 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_312 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_fill_1 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_328 ();
 sg13g2_fill_2 FILLER_69_335 ();
 sg13g2_fill_1 FILLER_69_337 ();
 sg13g2_decap_8 FILLER_69_346 ();
 sg13g2_decap_8 FILLER_69_353 ();
 sg13g2_decap_8 FILLER_69_360 ();
 sg13g2_decap_8 FILLER_69_367 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_4 FILLER_69_409 ();
 sg13g2_fill_1 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_fill_2 FILLER_69_430 ();
 sg13g2_decap_8 FILLER_69_440 ();
 sg13g2_decap_8 FILLER_69_447 ();
 sg13g2_decap_8 FILLER_69_454 ();
 sg13g2_decap_8 FILLER_69_461 ();
 sg13g2_fill_2 FILLER_69_468 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_decap_8 FILLER_69_485 ();
 sg13g2_decap_8 FILLER_69_492 ();
 sg13g2_decap_8 FILLER_69_499 ();
 sg13g2_decap_8 FILLER_69_506 ();
 sg13g2_fill_1 FILLER_69_513 ();
 sg13g2_decap_8 FILLER_69_531 ();
 sg13g2_decap_8 FILLER_69_538 ();
 sg13g2_decap_8 FILLER_69_545 ();
 sg13g2_decap_8 FILLER_69_552 ();
 sg13g2_decap_8 FILLER_69_559 ();
 sg13g2_decap_8 FILLER_69_566 ();
 sg13g2_decap_8 FILLER_69_573 ();
 sg13g2_decap_8 FILLER_69_580 ();
 sg13g2_fill_1 FILLER_69_593 ();
 sg13g2_fill_1 FILLER_69_597 ();
 sg13g2_decap_8 FILLER_69_618 ();
 sg13g2_decap_8 FILLER_69_625 ();
 sg13g2_decap_8 FILLER_69_632 ();
 sg13g2_fill_2 FILLER_69_639 ();
 sg13g2_fill_1 FILLER_69_641 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_decap_8 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_682 ();
 sg13g2_fill_2 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_691 ();
 sg13g2_decap_8 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_708 ();
 sg13g2_fill_1 FILLER_69_710 ();
 sg13g2_decap_4 FILLER_69_716 ();
 sg13g2_fill_2 FILLER_69_720 ();
 sg13g2_fill_1 FILLER_69_730 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_decap_8 FILLER_69_756 ();
 sg13g2_decap_8 FILLER_69_763 ();
 sg13g2_decap_8 FILLER_69_770 ();
 sg13g2_decap_4 FILLER_69_777 ();
 sg13g2_decap_8 FILLER_69_798 ();
 sg13g2_decap_8 FILLER_69_805 ();
 sg13g2_decap_8 FILLER_69_812 ();
 sg13g2_decap_8 FILLER_69_819 ();
 sg13g2_fill_2 FILLER_69_851 ();
 sg13g2_fill_1 FILLER_69_853 ();
 sg13g2_decap_8 FILLER_69_865 ();
 sg13g2_decap_4 FILLER_69_872 ();
 sg13g2_fill_2 FILLER_69_876 ();
 sg13g2_decap_4 FILLER_69_886 ();
 sg13g2_fill_2 FILLER_69_890 ();
 sg13g2_decap_8 FILLER_69_895 ();
 sg13g2_decap_8 FILLER_69_902 ();
 sg13g2_fill_2 FILLER_69_909 ();
 sg13g2_decap_8 FILLER_69_924 ();
 sg13g2_decap_8 FILLER_69_931 ();
 sg13g2_decap_8 FILLER_69_938 ();
 sg13g2_decap_8 FILLER_69_945 ();
 sg13g2_decap_8 FILLER_69_952 ();
 sg13g2_fill_1 FILLER_69_959 ();
 sg13g2_decap_8 FILLER_69_974 ();
 sg13g2_decap_8 FILLER_69_981 ();
 sg13g2_fill_1 FILLER_69_991 ();
 sg13g2_fill_2 FILLER_69_996 ();
 sg13g2_fill_1 FILLER_69_998 ();
 sg13g2_decap_8 FILLER_69_1037 ();
 sg13g2_decap_8 FILLER_69_1044 ();
 sg13g2_decap_8 FILLER_69_1051 ();
 sg13g2_decap_4 FILLER_69_1058 ();
 sg13g2_fill_1 FILLER_69_1062 ();
 sg13g2_decap_8 FILLER_69_1079 ();
 sg13g2_decap_8 FILLER_69_1086 ();
 sg13g2_decap_8 FILLER_69_1093 ();
 sg13g2_decap_4 FILLER_69_1100 ();
 sg13g2_decap_8 FILLER_69_1120 ();
 sg13g2_decap_8 FILLER_69_1127 ();
 sg13g2_decap_8 FILLER_69_1134 ();
 sg13g2_decap_8 FILLER_69_1141 ();
 sg13g2_decap_8 FILLER_69_1148 ();
 sg13g2_decap_8 FILLER_69_1155 ();
 sg13g2_decap_8 FILLER_69_1166 ();
 sg13g2_decap_8 FILLER_69_1173 ();
 sg13g2_decap_8 FILLER_69_1180 ();
 sg13g2_fill_2 FILLER_69_1187 ();
 sg13g2_fill_1 FILLER_69_1189 ();
 sg13g2_decap_8 FILLER_69_1203 ();
 sg13g2_decap_8 FILLER_69_1210 ();
 sg13g2_decap_8 FILLER_69_1217 ();
 sg13g2_decap_8 FILLER_69_1224 ();
 sg13g2_decap_8 FILLER_69_1231 ();
 sg13g2_decap_8 FILLER_69_1238 ();
 sg13g2_decap_8 FILLER_69_1245 ();
 sg13g2_decap_8 FILLER_69_1252 ();
 sg13g2_decap_4 FILLER_69_1259 ();
 sg13g2_fill_2 FILLER_69_1263 ();
 sg13g2_fill_1 FILLER_69_1277 ();
 sg13g2_decap_8 FILLER_69_1292 ();
 sg13g2_decap_4 FILLER_69_1299 ();
 sg13g2_decap_8 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_69_1318 ();
 sg13g2_fill_2 FILLER_69_1325 ();
 sg13g2_fill_1 FILLER_69_1327 ();
 sg13g2_decap_8 FILLER_69_1344 ();
 sg13g2_decap_8 FILLER_69_1351 ();
 sg13g2_decap_8 FILLER_69_1358 ();
 sg13g2_decap_8 FILLER_69_1365 ();
 sg13g2_decap_8 FILLER_69_1372 ();
 sg13g2_fill_2 FILLER_69_1379 ();
 sg13g2_decap_8 FILLER_69_1391 ();
 sg13g2_decap_8 FILLER_69_1398 ();
 sg13g2_fill_2 FILLER_69_1405 ();
 sg13g2_fill_1 FILLER_69_1407 ();
 sg13g2_fill_1 FILLER_69_1431 ();
 sg13g2_decap_8 FILLER_69_1440 ();
 sg13g2_decap_8 FILLER_69_1447 ();
 sg13g2_fill_1 FILLER_69_1454 ();
 sg13g2_decap_8 FILLER_69_1472 ();
 sg13g2_decap_8 FILLER_69_1479 ();
 sg13g2_decap_8 FILLER_69_1486 ();
 sg13g2_decap_8 FILLER_69_1493 ();
 sg13g2_fill_1 FILLER_69_1500 ();
 sg13g2_fill_2 FILLER_69_1514 ();
 sg13g2_fill_1 FILLER_69_1516 ();
 sg13g2_fill_2 FILLER_69_1523 ();
 sg13g2_fill_1 FILLER_69_1525 ();
 sg13g2_decap_8 FILLER_69_1542 ();
 sg13g2_decap_8 FILLER_69_1549 ();
 sg13g2_decap_8 FILLER_69_1556 ();
 sg13g2_fill_2 FILLER_69_1571 ();
 sg13g2_fill_1 FILLER_69_1573 ();
 sg13g2_decap_8 FILLER_69_1593 ();
 sg13g2_decap_8 FILLER_69_1600 ();
 sg13g2_decap_8 FILLER_69_1607 ();
 sg13g2_decap_8 FILLER_69_1614 ();
 sg13g2_decap_8 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1635 ();
 sg13g2_decap_8 FILLER_69_1642 ();
 sg13g2_decap_8 FILLER_69_1649 ();
 sg13g2_decap_8 FILLER_69_1681 ();
 sg13g2_decap_8 FILLER_69_1688 ();
 sg13g2_decap_8 FILLER_69_1695 ();
 sg13g2_decap_8 FILLER_69_1702 ();
 sg13g2_decap_8 FILLER_69_1709 ();
 sg13g2_decap_8 FILLER_69_1716 ();
 sg13g2_decap_8 FILLER_69_1723 ();
 sg13g2_decap_8 FILLER_69_1730 ();
 sg13g2_decap_8 FILLER_69_1737 ();
 sg13g2_decap_8 FILLER_69_1744 ();
 sg13g2_decap_8 FILLER_69_1751 ();
 sg13g2_decap_8 FILLER_69_1758 ();
 sg13g2_fill_2 FILLER_69_1765 ();
 sg13g2_fill_1 FILLER_69_1767 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_9 ();
 sg13g2_decap_8 FILLER_70_36 ();
 sg13g2_decap_8 FILLER_70_43 ();
 sg13g2_decap_8 FILLER_70_50 ();
 sg13g2_decap_8 FILLER_70_57 ();
 sg13g2_decap_4 FILLER_70_64 ();
 sg13g2_fill_2 FILLER_70_68 ();
 sg13g2_decap_4 FILLER_70_96 ();
 sg13g2_decap_4 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_187 ();
 sg13g2_decap_8 FILLER_70_194 ();
 sg13g2_decap_8 FILLER_70_201 ();
 sg13g2_decap_8 FILLER_70_208 ();
 sg13g2_decap_8 FILLER_70_215 ();
 sg13g2_decap_8 FILLER_70_222 ();
 sg13g2_decap_8 FILLER_70_229 ();
 sg13g2_decap_8 FILLER_70_236 ();
 sg13g2_decap_8 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_8 FILLER_70_264 ();
 sg13g2_decap_8 FILLER_70_271 ();
 sg13g2_decap_8 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_285 ();
 sg13g2_decap_8 FILLER_70_295 ();
 sg13g2_decap_8 FILLER_70_302 ();
 sg13g2_decap_8 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_316 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_2 FILLER_70_335 ();
 sg13g2_decap_8 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_354 ();
 sg13g2_fill_1 FILLER_70_361 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_376 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_fill_1 FILLER_70_390 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_4 FILLER_70_420 ();
 sg13g2_fill_2 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_446 ();
 sg13g2_fill_1 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_457 ();
 sg13g2_fill_2 FILLER_70_464 ();
 sg13g2_fill_1 FILLER_70_466 ();
 sg13g2_fill_2 FILLER_70_475 ();
 sg13g2_decap_8 FILLER_70_490 ();
 sg13g2_decap_8 FILLER_70_497 ();
 sg13g2_decap_8 FILLER_70_504 ();
 sg13g2_decap_4 FILLER_70_511 ();
 sg13g2_decap_8 FILLER_70_534 ();
 sg13g2_decap_8 FILLER_70_541 ();
 sg13g2_decap_8 FILLER_70_548 ();
 sg13g2_decap_8 FILLER_70_555 ();
 sg13g2_fill_2 FILLER_70_562 ();
 sg13g2_fill_1 FILLER_70_564 ();
 sg13g2_decap_4 FILLER_70_569 ();
 sg13g2_fill_2 FILLER_70_573 ();
 sg13g2_fill_2 FILLER_70_591 ();
 sg13g2_fill_1 FILLER_70_593 ();
 sg13g2_decap_4 FILLER_70_602 ();
 sg13g2_decap_4 FILLER_70_619 ();
 sg13g2_fill_2 FILLER_70_623 ();
 sg13g2_decap_8 FILLER_70_639 ();
 sg13g2_fill_2 FILLER_70_646 ();
 sg13g2_fill_1 FILLER_70_648 ();
 sg13g2_decap_8 FILLER_70_654 ();
 sg13g2_decap_4 FILLER_70_661 ();
 sg13g2_fill_2 FILLER_70_677 ();
 sg13g2_decap_8 FILLER_70_700 ();
 sg13g2_fill_1 FILLER_70_707 ();
 sg13g2_decap_8 FILLER_70_730 ();
 sg13g2_decap_8 FILLER_70_737 ();
 sg13g2_decap_8 FILLER_70_744 ();
 sg13g2_decap_8 FILLER_70_751 ();
 sg13g2_decap_8 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_765 ();
 sg13g2_fill_2 FILLER_70_772 ();
 sg13g2_decap_8 FILLER_70_789 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_817 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_fill_2 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_8 FILLER_70_856 ();
 sg13g2_decap_8 FILLER_70_863 ();
 sg13g2_decap_8 FILLER_70_870 ();
 sg13g2_fill_2 FILLER_70_877 ();
 sg13g2_fill_1 FILLER_70_895 ();
 sg13g2_decap_8 FILLER_70_914 ();
 sg13g2_decap_8 FILLER_70_921 ();
 sg13g2_decap_4 FILLER_70_928 ();
 sg13g2_fill_1 FILLER_70_932 ();
 sg13g2_fill_2 FILLER_70_941 ();
 sg13g2_decap_8 FILLER_70_949 ();
 sg13g2_decap_8 FILLER_70_956 ();
 sg13g2_fill_2 FILLER_70_963 ();
 sg13g2_fill_1 FILLER_70_965 ();
 sg13g2_decap_8 FILLER_70_972 ();
 sg13g2_decap_8 FILLER_70_979 ();
 sg13g2_decap_8 FILLER_70_986 ();
 sg13g2_decap_8 FILLER_70_993 ();
 sg13g2_decap_8 FILLER_70_1000 ();
 sg13g2_fill_2 FILLER_70_1007 ();
 sg13g2_fill_1 FILLER_70_1009 ();
 sg13g2_decap_8 FILLER_70_1028 ();
 sg13g2_decap_8 FILLER_70_1035 ();
 sg13g2_decap_8 FILLER_70_1042 ();
 sg13g2_decap_8 FILLER_70_1049 ();
 sg13g2_decap_8 FILLER_70_1056 ();
 sg13g2_decap_4 FILLER_70_1063 ();
 sg13g2_fill_2 FILLER_70_1072 ();
 sg13g2_fill_1 FILLER_70_1074 ();
 sg13g2_decap_8 FILLER_70_1083 ();
 sg13g2_decap_8 FILLER_70_1090 ();
 sg13g2_decap_4 FILLER_70_1097 ();
 sg13g2_fill_1 FILLER_70_1101 ();
 sg13g2_decap_8 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_decap_8 FILLER_70_1137 ();
 sg13g2_decap_4 FILLER_70_1152 ();
 sg13g2_fill_1 FILLER_70_1156 ();
 sg13g2_fill_1 FILLER_70_1162 ();
 sg13g2_fill_1 FILLER_70_1173 ();
 sg13g2_decap_8 FILLER_70_1203 ();
 sg13g2_decap_8 FILLER_70_1210 ();
 sg13g2_decap_8 FILLER_70_1217 ();
 sg13g2_decap_8 FILLER_70_1224 ();
 sg13g2_decap_8 FILLER_70_1231 ();
 sg13g2_decap_8 FILLER_70_1238 ();
 sg13g2_decap_8 FILLER_70_1245 ();
 sg13g2_fill_1 FILLER_70_1252 ();
 sg13g2_fill_1 FILLER_70_1263 ();
 sg13g2_decap_4 FILLER_70_1274 ();
 sg13g2_fill_1 FILLER_70_1278 ();
 sg13g2_decap_4 FILLER_70_1290 ();
 sg13g2_fill_1 FILLER_70_1307 ();
 sg13g2_decap_8 FILLER_70_1316 ();
 sg13g2_decap_8 FILLER_70_1323 ();
 sg13g2_decap_4 FILLER_70_1330 ();
 sg13g2_fill_1 FILLER_70_1334 ();
 sg13g2_decap_8 FILLER_70_1340 ();
 sg13g2_decap_8 FILLER_70_1347 ();
 sg13g2_decap_8 FILLER_70_1354 ();
 sg13g2_decap_8 FILLER_70_1361 ();
 sg13g2_decap_4 FILLER_70_1368 ();
 sg13g2_fill_1 FILLER_70_1372 ();
 sg13g2_decap_8 FILLER_70_1377 ();
 sg13g2_decap_8 FILLER_70_1384 ();
 sg13g2_decap_8 FILLER_70_1391 ();
 sg13g2_decap_4 FILLER_70_1398 ();
 sg13g2_fill_2 FILLER_70_1402 ();
 sg13g2_decap_8 FILLER_70_1412 ();
 sg13g2_decap_4 FILLER_70_1419 ();
 sg13g2_fill_2 FILLER_70_1423 ();
 sg13g2_decap_8 FILLER_70_1439 ();
 sg13g2_decap_8 FILLER_70_1446 ();
 sg13g2_fill_2 FILLER_70_1453 ();
 sg13g2_fill_1 FILLER_70_1455 ();
 sg13g2_decap_8 FILLER_70_1486 ();
 sg13g2_decap_8 FILLER_70_1493 ();
 sg13g2_decap_8 FILLER_70_1500 ();
 sg13g2_fill_1 FILLER_70_1507 ();
 sg13g2_fill_1 FILLER_70_1520 ();
 sg13g2_decap_8 FILLER_70_1525 ();
 sg13g2_decap_8 FILLER_70_1532 ();
 sg13g2_decap_8 FILLER_70_1539 ();
 sg13g2_decap_8 FILLER_70_1546 ();
 sg13g2_decap_8 FILLER_70_1553 ();
 sg13g2_decap_8 FILLER_70_1560 ();
 sg13g2_decap_8 FILLER_70_1567 ();
 sg13g2_decap_8 FILLER_70_1582 ();
 sg13g2_decap_8 FILLER_70_1589 ();
 sg13g2_fill_2 FILLER_70_1596 ();
 sg13g2_decap_8 FILLER_70_1606 ();
 sg13g2_decap_8 FILLER_70_1613 ();
 sg13g2_decap_8 FILLER_70_1620 ();
 sg13g2_decap_8 FILLER_70_1627 ();
 sg13g2_decap_8 FILLER_70_1634 ();
 sg13g2_decap_8 FILLER_70_1667 ();
 sg13g2_decap_8 FILLER_70_1674 ();
 sg13g2_decap_8 FILLER_70_1681 ();
 sg13g2_decap_8 FILLER_70_1688 ();
 sg13g2_fill_1 FILLER_70_1695 ();
 sg13g2_decap_8 FILLER_70_1700 ();
 sg13g2_decap_8 FILLER_70_1707 ();
 sg13g2_decap_8 FILLER_70_1714 ();
 sg13g2_decap_8 FILLER_70_1721 ();
 sg13g2_decap_8 FILLER_70_1728 ();
 sg13g2_decap_8 FILLER_70_1735 ();
 sg13g2_decap_8 FILLER_70_1742 ();
 sg13g2_decap_8 FILLER_70_1749 ();
 sg13g2_decap_8 FILLER_70_1756 ();
 sg13g2_decap_4 FILLER_70_1763 ();
 sg13g2_fill_1 FILLER_70_1767 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_25 ();
 sg13g2_decap_8 FILLER_71_32 ();
 sg13g2_decap_8 FILLER_71_39 ();
 sg13g2_decap_8 FILLER_71_46 ();
 sg13g2_decap_8 FILLER_71_53 ();
 sg13g2_decap_8 FILLER_71_60 ();
 sg13g2_decap_8 FILLER_71_67 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_decap_8 FILLER_71_81 ();
 sg13g2_decap_8 FILLER_71_88 ();
 sg13g2_decap_8 FILLER_71_95 ();
 sg13g2_decap_4 FILLER_71_102 ();
 sg13g2_fill_1 FILLER_71_106 ();
 sg13g2_decap_8 FILLER_71_136 ();
 sg13g2_decap_8 FILLER_71_143 ();
 sg13g2_decap_4 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_154 ();
 sg13g2_decap_4 FILLER_71_166 ();
 sg13g2_fill_2 FILLER_71_170 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_4 FILLER_71_183 ();
 sg13g2_fill_1 FILLER_71_187 ();
 sg13g2_decap_8 FILLER_71_201 ();
 sg13g2_decap_8 FILLER_71_208 ();
 sg13g2_decap_8 FILLER_71_215 ();
 sg13g2_decap_8 FILLER_71_222 ();
 sg13g2_fill_2 FILLER_71_229 ();
 sg13g2_decap_8 FILLER_71_244 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_decap_8 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_281 ();
 sg13g2_fill_1 FILLER_71_288 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_4 FILLER_71_299 ();
 sg13g2_fill_1 FILLER_71_303 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_fill_2 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_352 ();
 sg13g2_fill_1 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_387 ();
 sg13g2_fill_2 FILLER_71_394 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_decap_8 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_424 ();
 sg13g2_decap_8 FILLER_71_437 ();
 sg13g2_decap_8 FILLER_71_444 ();
 sg13g2_decap_8 FILLER_71_451 ();
 sg13g2_decap_4 FILLER_71_458 ();
 sg13g2_fill_2 FILLER_71_475 ();
 sg13g2_fill_2 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_495 ();
 sg13g2_fill_2 FILLER_71_502 ();
 sg13g2_fill_1 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_537 ();
 sg13g2_decap_8 FILLER_71_544 ();
 sg13g2_decap_8 FILLER_71_551 ();
 sg13g2_fill_2 FILLER_71_558 ();
 sg13g2_fill_1 FILLER_71_560 ();
 sg13g2_fill_1 FILLER_71_573 ();
 sg13g2_decap_8 FILLER_71_584 ();
 sg13g2_decap_8 FILLER_71_591 ();
 sg13g2_decap_4 FILLER_71_598 ();
 sg13g2_fill_2 FILLER_71_602 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_decap_8 FILLER_71_624 ();
 sg13g2_decap_8 FILLER_71_631 ();
 sg13g2_decap_8 FILLER_71_638 ();
 sg13g2_decap_8 FILLER_71_645 ();
 sg13g2_decap_8 FILLER_71_652 ();
 sg13g2_fill_2 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_661 ();
 sg13g2_decap_8 FILLER_71_666 ();
 sg13g2_decap_8 FILLER_71_673 ();
 sg13g2_fill_2 FILLER_71_680 ();
 sg13g2_fill_1 FILLER_71_682 ();
 sg13g2_decap_8 FILLER_71_696 ();
 sg13g2_decap_8 FILLER_71_703 ();
 sg13g2_decap_8 FILLER_71_710 ();
 sg13g2_decap_8 FILLER_71_717 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_8 FILLER_71_748 ();
 sg13g2_decap_4 FILLER_71_755 ();
 sg13g2_fill_1 FILLER_71_759 ();
 sg13g2_decap_8 FILLER_71_766 ();
 sg13g2_decap_8 FILLER_71_773 ();
 sg13g2_decap_4 FILLER_71_780 ();
 sg13g2_fill_1 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_decap_8 FILLER_71_807 ();
 sg13g2_decap_8 FILLER_71_822 ();
 sg13g2_decap_4 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_fill_1 FILLER_71_878 ();
 sg13g2_decap_8 FILLER_71_900 ();
 sg13g2_decap_8 FILLER_71_907 ();
 sg13g2_decap_8 FILLER_71_914 ();
 sg13g2_decap_8 FILLER_71_921 ();
 sg13g2_decap_8 FILLER_71_928 ();
 sg13g2_decap_8 FILLER_71_959 ();
 sg13g2_fill_2 FILLER_71_966 ();
 sg13g2_decap_8 FILLER_71_976 ();
 sg13g2_decap_8 FILLER_71_983 ();
 sg13g2_decap_8 FILLER_71_990 ();
 sg13g2_decap_8 FILLER_71_997 ();
 sg13g2_decap_8 FILLER_71_1028 ();
 sg13g2_decap_8 FILLER_71_1035 ();
 sg13g2_decap_8 FILLER_71_1042 ();
 sg13g2_decap_8 FILLER_71_1049 ();
 sg13g2_decap_8 FILLER_71_1056 ();
 sg13g2_decap_4 FILLER_71_1063 ();
 sg13g2_decap_4 FILLER_71_1085 ();
 sg13g2_fill_1 FILLER_71_1089 ();
 sg13g2_decap_8 FILLER_71_1100 ();
 sg13g2_decap_8 FILLER_71_1124 ();
 sg13g2_decap_8 FILLER_71_1131 ();
 sg13g2_decap_8 FILLER_71_1138 ();
 sg13g2_decap_4 FILLER_71_1145 ();
 sg13g2_fill_1 FILLER_71_1149 ();
 sg13g2_decap_8 FILLER_71_1154 ();
 sg13g2_decap_8 FILLER_71_1161 ();
 sg13g2_decap_8 FILLER_71_1168 ();
 sg13g2_decap_8 FILLER_71_1175 ();
 sg13g2_decap_4 FILLER_71_1182 ();
 sg13g2_fill_1 FILLER_71_1186 ();
 sg13g2_decap_4 FILLER_71_1196 ();
 sg13g2_fill_1 FILLER_71_1200 ();
 sg13g2_decap_8 FILLER_71_1219 ();
 sg13g2_decap_4 FILLER_71_1226 ();
 sg13g2_fill_1 FILLER_71_1230 ();
 sg13g2_fill_2 FILLER_71_1244 ();
 sg13g2_fill_1 FILLER_71_1246 ();
 sg13g2_decap_8 FILLER_71_1261 ();
 sg13g2_fill_2 FILLER_71_1268 ();
 sg13g2_fill_1 FILLER_71_1270 ();
 sg13g2_fill_2 FILLER_71_1279 ();
 sg13g2_fill_1 FILLER_71_1281 ();
 sg13g2_decap_8 FILLER_71_1288 ();
 sg13g2_decap_8 FILLER_71_1295 ();
 sg13g2_fill_1 FILLER_71_1302 ();
 sg13g2_decap_8 FILLER_71_1313 ();
 sg13g2_decap_8 FILLER_71_1320 ();
 sg13g2_decap_8 FILLER_71_1327 ();
 sg13g2_decap_8 FILLER_71_1334 ();
 sg13g2_decap_8 FILLER_71_1341 ();
 sg13g2_fill_1 FILLER_71_1348 ();
 sg13g2_decap_8 FILLER_71_1357 ();
 sg13g2_decap_8 FILLER_71_1364 ();
 sg13g2_fill_2 FILLER_71_1371 ();
 sg13g2_fill_1 FILLER_71_1373 ();
 sg13g2_fill_2 FILLER_71_1377 ();
 sg13g2_fill_1 FILLER_71_1379 ();
 sg13g2_decap_8 FILLER_71_1385 ();
 sg13g2_decap_8 FILLER_71_1392 ();
 sg13g2_decap_4 FILLER_71_1399 ();
 sg13g2_fill_2 FILLER_71_1403 ();
 sg13g2_decap_8 FILLER_71_1416 ();
 sg13g2_decap_8 FILLER_71_1423 ();
 sg13g2_decap_4 FILLER_71_1430 ();
 sg13g2_fill_2 FILLER_71_1462 ();
 sg13g2_decap_8 FILLER_71_1472 ();
 sg13g2_decap_8 FILLER_71_1479 ();
 sg13g2_decap_8 FILLER_71_1486 ();
 sg13g2_decap_8 FILLER_71_1493 ();
 sg13g2_decap_8 FILLER_71_1512 ();
 sg13g2_decap_4 FILLER_71_1519 ();
 sg13g2_fill_2 FILLER_71_1523 ();
 sg13g2_decap_8 FILLER_71_1533 ();
 sg13g2_decap_8 FILLER_71_1540 ();
 sg13g2_decap_8 FILLER_71_1547 ();
 sg13g2_decap_4 FILLER_71_1554 ();
 sg13g2_fill_1 FILLER_71_1558 ();
 sg13g2_decap_8 FILLER_71_1571 ();
 sg13g2_decap_8 FILLER_71_1578 ();
 sg13g2_decap_8 FILLER_71_1585 ();
 sg13g2_fill_2 FILLER_71_1592 ();
 sg13g2_fill_1 FILLER_71_1594 ();
 sg13g2_decap_8 FILLER_71_1611 ();
 sg13g2_decap_8 FILLER_71_1618 ();
 sg13g2_decap_8 FILLER_71_1625 ();
 sg13g2_decap_8 FILLER_71_1632 ();
 sg13g2_decap_8 FILLER_71_1639 ();
 sg13g2_decap_4 FILLER_71_1646 ();
 sg13g2_fill_2 FILLER_71_1650 ();
 sg13g2_decap_8 FILLER_71_1656 ();
 sg13g2_decap_8 FILLER_71_1663 ();
 sg13g2_decap_8 FILLER_71_1670 ();
 sg13g2_decap_8 FILLER_71_1677 ();
 sg13g2_fill_1 FILLER_71_1684 ();
 sg13g2_decap_8 FILLER_71_1724 ();
 sg13g2_decap_8 FILLER_71_1731 ();
 sg13g2_decap_8 FILLER_71_1738 ();
 sg13g2_decap_8 FILLER_71_1745 ();
 sg13g2_decap_8 FILLER_71_1752 ();
 sg13g2_decap_8 FILLER_71_1759 ();
 sg13g2_fill_2 FILLER_71_1766 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_fill_1 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_54 ();
 sg13g2_decap_8 FILLER_72_61 ();
 sg13g2_decap_8 FILLER_72_68 ();
 sg13g2_decap_8 FILLER_72_75 ();
 sg13g2_decap_8 FILLER_72_82 ();
 sg13g2_decap_8 FILLER_72_89 ();
 sg13g2_decap_8 FILLER_72_96 ();
 sg13g2_decap_8 FILLER_72_103 ();
 sg13g2_decap_8 FILLER_72_110 ();
 sg13g2_decap_8 FILLER_72_117 ();
 sg13g2_decap_8 FILLER_72_124 ();
 sg13g2_decap_8 FILLER_72_131 ();
 sg13g2_decap_8 FILLER_72_138 ();
 sg13g2_decap_8 FILLER_72_145 ();
 sg13g2_decap_8 FILLER_72_152 ();
 sg13g2_decap_8 FILLER_72_159 ();
 sg13g2_decap_8 FILLER_72_166 ();
 sg13g2_decap_8 FILLER_72_173 ();
 sg13g2_decap_8 FILLER_72_180 ();
 sg13g2_decap_8 FILLER_72_187 ();
 sg13g2_decap_8 FILLER_72_194 ();
 sg13g2_decap_8 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_208 ();
 sg13g2_decap_8 FILLER_72_221 ();
 sg13g2_decap_4 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_232 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_261 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_299 ();
 sg13g2_decap_8 FILLER_72_306 ();
 sg13g2_decap_8 FILLER_72_313 ();
 sg13g2_decap_4 FILLER_72_320 ();
 sg13g2_decap_8 FILLER_72_333 ();
 sg13g2_decap_4 FILLER_72_340 ();
 sg13g2_decap_8 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_4 FILLER_72_377 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_fill_1 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_436 ();
 sg13g2_decap_8 FILLER_72_443 ();
 sg13g2_decap_8 FILLER_72_450 ();
 sg13g2_fill_1 FILLER_72_457 ();
 sg13g2_fill_2 FILLER_72_480 ();
 sg13g2_fill_1 FILLER_72_482 ();
 sg13g2_decap_8 FILLER_72_489 ();
 sg13g2_decap_4 FILLER_72_496 ();
 sg13g2_fill_2 FILLER_72_500 ();
 sg13g2_decap_8 FILLER_72_510 ();
 sg13g2_decap_8 FILLER_72_517 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_538 ();
 sg13g2_decap_8 FILLER_72_545 ();
 sg13g2_decap_8 FILLER_72_552 ();
 sg13g2_decap_4 FILLER_72_559 ();
 sg13g2_fill_2 FILLER_72_563 ();
 sg13g2_decap_4 FILLER_72_568 ();
 sg13g2_fill_1 FILLER_72_572 ();
 sg13g2_fill_1 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_588 ();
 sg13g2_decap_8 FILLER_72_595 ();
 sg13g2_decap_8 FILLER_72_602 ();
 sg13g2_decap_4 FILLER_72_609 ();
 sg13g2_decap_8 FILLER_72_628 ();
 sg13g2_decap_8 FILLER_72_635 ();
 sg13g2_decap_8 FILLER_72_642 ();
 sg13g2_decap_8 FILLER_72_649 ();
 sg13g2_decap_4 FILLER_72_656 ();
 sg13g2_fill_1 FILLER_72_660 ();
 sg13g2_decap_8 FILLER_72_667 ();
 sg13g2_fill_2 FILLER_72_674 ();
 sg13g2_fill_1 FILLER_72_684 ();
 sg13g2_decap_8 FILLER_72_690 ();
 sg13g2_decap_8 FILLER_72_697 ();
 sg13g2_decap_8 FILLER_72_704 ();
 sg13g2_decap_8 FILLER_72_711 ();
 sg13g2_decap_8 FILLER_72_718 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_decap_8 FILLER_72_732 ();
 sg13g2_fill_2 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_814 ();
 sg13g2_fill_2 FILLER_72_821 ();
 sg13g2_fill_1 FILLER_72_823 ();
 sg13g2_decap_8 FILLER_72_835 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_8 FILLER_72_856 ();
 sg13g2_decap_8 FILLER_72_863 ();
 sg13g2_fill_1 FILLER_72_870 ();
 sg13g2_decap_8 FILLER_72_879 ();
 sg13g2_decap_8 FILLER_72_886 ();
 sg13g2_decap_8 FILLER_72_893 ();
 sg13g2_decap_8 FILLER_72_900 ();
 sg13g2_decap_8 FILLER_72_907 ();
 sg13g2_decap_8 FILLER_72_914 ();
 sg13g2_decap_8 FILLER_72_921 ();
 sg13g2_decap_8 FILLER_72_928 ();
 sg13g2_decap_8 FILLER_72_935 ();
 sg13g2_fill_1 FILLER_72_942 ();
 sg13g2_fill_2 FILLER_72_949 ();
 sg13g2_fill_1 FILLER_72_951 ();
 sg13g2_decap_8 FILLER_72_965 ();
 sg13g2_fill_1 FILLER_72_972 ();
 sg13g2_decap_8 FILLER_72_982 ();
 sg13g2_decap_8 FILLER_72_994 ();
 sg13g2_decap_4 FILLER_72_1001 ();
 sg13g2_fill_1 FILLER_72_1005 ();
 sg13g2_decap_8 FILLER_72_1014 ();
 sg13g2_decap_8 FILLER_72_1021 ();
 sg13g2_decap_8 FILLER_72_1028 ();
 sg13g2_decap_8 FILLER_72_1035 ();
 sg13g2_fill_2 FILLER_72_1042 ();
 sg13g2_fill_1 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1053 ();
 sg13g2_decap_8 FILLER_72_1060 ();
 sg13g2_decap_8 FILLER_72_1067 ();
 sg13g2_decap_8 FILLER_72_1080 ();
 sg13g2_fill_2 FILLER_72_1087 ();
 sg13g2_decap_8 FILLER_72_1093 ();
 sg13g2_decap_8 FILLER_72_1100 ();
 sg13g2_decap_4 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1119 ();
 sg13g2_decap_8 FILLER_72_1126 ();
 sg13g2_decap_8 FILLER_72_1133 ();
 sg13g2_decap_8 FILLER_72_1140 ();
 sg13g2_decap_8 FILLER_72_1147 ();
 sg13g2_decap_8 FILLER_72_1154 ();
 sg13g2_decap_8 FILLER_72_1187 ();
 sg13g2_decap_8 FILLER_72_1194 ();
 sg13g2_decap_8 FILLER_72_1201 ();
 sg13g2_decap_8 FILLER_72_1208 ();
 sg13g2_decap_4 FILLER_72_1215 ();
 sg13g2_decap_8 FILLER_72_1224 ();
 sg13g2_decap_8 FILLER_72_1231 ();
 sg13g2_decap_8 FILLER_72_1238 ();
 sg13g2_fill_2 FILLER_72_1245 ();
 sg13g2_fill_2 FILLER_72_1257 ();
 sg13g2_fill_1 FILLER_72_1259 ();
 sg13g2_decap_8 FILLER_72_1281 ();
 sg13g2_decap_4 FILLER_72_1288 ();
 sg13g2_fill_1 FILLER_72_1292 ();
 sg13g2_decap_8 FILLER_72_1301 ();
 sg13g2_decap_8 FILLER_72_1308 ();
 sg13g2_decap_8 FILLER_72_1315 ();
 sg13g2_decap_8 FILLER_72_1322 ();
 sg13g2_decap_8 FILLER_72_1329 ();
 sg13g2_decap_4 FILLER_72_1336 ();
 sg13g2_fill_1 FILLER_72_1340 ();
 sg13g2_decap_8 FILLER_72_1354 ();
 sg13g2_decap_8 FILLER_72_1361 ();
 sg13g2_decap_4 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1372 ();
 sg13g2_decap_8 FILLER_72_1392 ();
 sg13g2_decap_8 FILLER_72_1399 ();
 sg13g2_decap_8 FILLER_72_1406 ();
 sg13g2_decap_8 FILLER_72_1413 ();
 sg13g2_decap_8 FILLER_72_1420 ();
 sg13g2_decap_8 FILLER_72_1427 ();
 sg13g2_decap_8 FILLER_72_1434 ();
 sg13g2_decap_8 FILLER_72_1441 ();
 sg13g2_decap_8 FILLER_72_1448 ();
 sg13g2_decap_8 FILLER_72_1455 ();
 sg13g2_decap_8 FILLER_72_1462 ();
 sg13g2_decap_8 FILLER_72_1469 ();
 sg13g2_decap_4 FILLER_72_1476 ();
 sg13g2_decap_8 FILLER_72_1488 ();
 sg13g2_decap_8 FILLER_72_1495 ();
 sg13g2_decap_8 FILLER_72_1502 ();
 sg13g2_decap_8 FILLER_72_1509 ();
 sg13g2_decap_8 FILLER_72_1516 ();
 sg13g2_decap_8 FILLER_72_1523 ();
 sg13g2_decap_8 FILLER_72_1530 ();
 sg13g2_decap_8 FILLER_72_1537 ();
 sg13g2_decap_4 FILLER_72_1544 ();
 sg13g2_fill_2 FILLER_72_1548 ();
 sg13g2_decap_8 FILLER_72_1575 ();
 sg13g2_decap_8 FILLER_72_1582 ();
 sg13g2_decap_8 FILLER_72_1589 ();
 sg13g2_decap_4 FILLER_72_1596 ();
 sg13g2_fill_2 FILLER_72_1600 ();
 sg13g2_decap_8 FILLER_72_1615 ();
 sg13g2_decap_8 FILLER_72_1622 ();
 sg13g2_decap_8 FILLER_72_1629 ();
 sg13g2_decap_8 FILLER_72_1636 ();
 sg13g2_fill_2 FILLER_72_1643 ();
 sg13g2_fill_1 FILLER_72_1645 ();
 sg13g2_fill_2 FILLER_72_1671 ();
 sg13g2_decap_8 FILLER_72_1683 ();
 sg13g2_decap_8 FILLER_72_1690 ();
 sg13g2_decap_8 FILLER_72_1697 ();
 sg13g2_decap_8 FILLER_72_1704 ();
 sg13g2_decap_8 FILLER_72_1720 ();
 sg13g2_decap_8 FILLER_72_1727 ();
 sg13g2_decap_8 FILLER_72_1734 ();
 sg13g2_decap_8 FILLER_72_1741 ();
 sg13g2_decap_8 FILLER_72_1748 ();
 sg13g2_decap_8 FILLER_72_1755 ();
 sg13g2_decap_4 FILLER_72_1762 ();
 sg13g2_fill_2 FILLER_72_1766 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_41 ();
 sg13g2_fill_2 FILLER_73_54 ();
 sg13g2_decap_8 FILLER_73_60 ();
 sg13g2_decap_8 FILLER_73_67 ();
 sg13g2_decap_4 FILLER_73_74 ();
 sg13g2_fill_1 FILLER_73_78 ();
 sg13g2_decap_8 FILLER_73_95 ();
 sg13g2_decap_8 FILLER_73_102 ();
 sg13g2_decap_8 FILLER_73_109 ();
 sg13g2_decap_8 FILLER_73_116 ();
 sg13g2_decap_8 FILLER_73_136 ();
 sg13g2_decap_8 FILLER_73_143 ();
 sg13g2_fill_1 FILLER_73_150 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_fill_2 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_194 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_fill_1 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_215 ();
 sg13g2_decap_8 FILLER_73_222 ();
 sg13g2_decap_4 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_243 ();
 sg13g2_decap_8 FILLER_73_248 ();
 sg13g2_fill_2 FILLER_73_282 ();
 sg13g2_fill_1 FILLER_73_284 ();
 sg13g2_decap_8 FILLER_73_300 ();
 sg13g2_decap_8 FILLER_73_307 ();
 sg13g2_fill_2 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_335 ();
 sg13g2_decap_8 FILLER_73_361 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_fill_2 FILLER_73_403 ();
 sg13g2_fill_1 FILLER_73_405 ();
 sg13g2_fill_1 FILLER_73_422 ();
 sg13g2_decap_8 FILLER_73_433 ();
 sg13g2_decap_8 FILLER_73_440 ();
 sg13g2_decap_8 FILLER_73_447 ();
 sg13g2_decap_8 FILLER_73_454 ();
 sg13g2_decap_4 FILLER_73_461 ();
 sg13g2_fill_1 FILLER_73_465 ();
 sg13g2_fill_2 FILLER_73_475 ();
 sg13g2_decap_8 FILLER_73_487 ();
 sg13g2_decap_8 FILLER_73_494 ();
 sg13g2_decap_8 FILLER_73_501 ();
 sg13g2_decap_4 FILLER_73_508 ();
 sg13g2_fill_1 FILLER_73_512 ();
 sg13g2_decap_8 FILLER_73_521 ();
 sg13g2_decap_8 FILLER_73_528 ();
 sg13g2_decap_8 FILLER_73_535 ();
 sg13g2_decap_4 FILLER_73_542 ();
 sg13g2_decap_8 FILLER_73_558 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_decap_8 FILLER_73_599 ();
 sg13g2_decap_8 FILLER_73_606 ();
 sg13g2_decap_8 FILLER_73_613 ();
 sg13g2_decap_8 FILLER_73_620 ();
 sg13g2_decap_8 FILLER_73_627 ();
 sg13g2_decap_8 FILLER_73_634 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_decap_8 FILLER_73_648 ();
 sg13g2_decap_8 FILLER_73_655 ();
 sg13g2_fill_1 FILLER_73_662 ();
 sg13g2_decap_8 FILLER_73_677 ();
 sg13g2_decap_8 FILLER_73_684 ();
 sg13g2_decap_4 FILLER_73_704 ();
 sg13g2_fill_2 FILLER_73_708 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_fill_1 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_742 ();
 sg13g2_decap_8 FILLER_73_749 ();
 sg13g2_decap_8 FILLER_73_756 ();
 sg13g2_decap_8 FILLER_73_763 ();
 sg13g2_decap_4 FILLER_73_770 ();
 sg13g2_decap_8 FILLER_73_778 ();
 sg13g2_decap_8 FILLER_73_785 ();
 sg13g2_decap_8 FILLER_73_792 ();
 sg13g2_decap_8 FILLER_73_799 ();
 sg13g2_fill_2 FILLER_73_806 ();
 sg13g2_fill_1 FILLER_73_808 ();
 sg13g2_fill_2 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_decap_8 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_73_868 ();
 sg13g2_decap_8 FILLER_73_875 ();
 sg13g2_decap_8 FILLER_73_882 ();
 sg13g2_decap_8 FILLER_73_915 ();
 sg13g2_decap_8 FILLER_73_922 ();
 sg13g2_decap_8 FILLER_73_929 ();
 sg13g2_fill_1 FILLER_73_936 ();
 sg13g2_decap_8 FILLER_73_942 ();
 sg13g2_decap_4 FILLER_73_949 ();
 sg13g2_fill_2 FILLER_73_961 ();
 sg13g2_fill_1 FILLER_73_963 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_decap_8 FILLER_73_1002 ();
 sg13g2_decap_8 FILLER_73_1009 ();
 sg13g2_decap_8 FILLER_73_1016 ();
 sg13g2_decap_8 FILLER_73_1023 ();
 sg13g2_decap_8 FILLER_73_1030 ();
 sg13g2_decap_8 FILLER_73_1037 ();
 sg13g2_decap_8 FILLER_73_1044 ();
 sg13g2_decap_8 FILLER_73_1051 ();
 sg13g2_decap_8 FILLER_73_1058 ();
 sg13g2_decap_8 FILLER_73_1065 ();
 sg13g2_decap_8 FILLER_73_1072 ();
 sg13g2_decap_8 FILLER_73_1079 ();
 sg13g2_decap_8 FILLER_73_1086 ();
 sg13g2_fill_2 FILLER_73_1093 ();
 sg13g2_fill_1 FILLER_73_1095 ();
 sg13g2_fill_1 FILLER_73_1121 ();
 sg13g2_decap_8 FILLER_73_1127 ();
 sg13g2_decap_4 FILLER_73_1134 ();
 sg13g2_fill_2 FILLER_73_1138 ();
 sg13g2_decap_8 FILLER_73_1175 ();
 sg13g2_decap_8 FILLER_73_1182 ();
 sg13g2_decap_8 FILLER_73_1189 ();
 sg13g2_decap_8 FILLER_73_1196 ();
 sg13g2_decap_8 FILLER_73_1203 ();
 sg13g2_fill_2 FILLER_73_1210 ();
 sg13g2_decap_8 FILLER_73_1255 ();
 sg13g2_decap_8 FILLER_73_1262 ();
 sg13g2_fill_1 FILLER_73_1269 ();
 sg13g2_decap_8 FILLER_73_1274 ();
 sg13g2_decap_8 FILLER_73_1281 ();
 sg13g2_decap_8 FILLER_73_1288 ();
 sg13g2_decap_8 FILLER_73_1295 ();
 sg13g2_decap_8 FILLER_73_1302 ();
 sg13g2_decap_4 FILLER_73_1309 ();
 sg13g2_fill_2 FILLER_73_1313 ();
 sg13g2_fill_1 FILLER_73_1319 ();
 sg13g2_fill_2 FILLER_73_1325 ();
 sg13g2_fill_1 FILLER_73_1327 ();
 sg13g2_decap_8 FILLER_73_1354 ();
 sg13g2_decap_8 FILLER_73_1374 ();
 sg13g2_decap_8 FILLER_73_1381 ();
 sg13g2_decap_8 FILLER_73_1388 ();
 sg13g2_fill_2 FILLER_73_1395 ();
 sg13g2_fill_1 FILLER_73_1397 ();
 sg13g2_fill_1 FILLER_73_1402 ();
 sg13g2_decap_8 FILLER_73_1411 ();
 sg13g2_decap_8 FILLER_73_1418 ();
 sg13g2_decap_8 FILLER_73_1425 ();
 sg13g2_decap_8 FILLER_73_1432 ();
 sg13g2_decap_8 FILLER_73_1439 ();
 sg13g2_decap_8 FILLER_73_1446 ();
 sg13g2_decap_8 FILLER_73_1453 ();
 sg13g2_decap_8 FILLER_73_1460 ();
 sg13g2_decap_8 FILLER_73_1467 ();
 sg13g2_decap_8 FILLER_73_1474 ();
 sg13g2_decap_8 FILLER_73_1481 ();
 sg13g2_decap_8 FILLER_73_1488 ();
 sg13g2_decap_8 FILLER_73_1495 ();
 sg13g2_decap_4 FILLER_73_1502 ();
 sg13g2_fill_1 FILLER_73_1506 ();
 sg13g2_decap_8 FILLER_73_1515 ();
 sg13g2_decap_8 FILLER_73_1522 ();
 sg13g2_decap_8 FILLER_73_1529 ();
 sg13g2_decap_8 FILLER_73_1536 ();
 sg13g2_decap_8 FILLER_73_1543 ();
 sg13g2_fill_2 FILLER_73_1550 ();
 sg13g2_fill_1 FILLER_73_1552 ();
 sg13g2_fill_1 FILLER_73_1562 ();
 sg13g2_decap_8 FILLER_73_1571 ();
 sg13g2_decap_8 FILLER_73_1578 ();
 sg13g2_decap_4 FILLER_73_1585 ();
 sg13g2_decap_8 FILLER_73_1597 ();
 sg13g2_fill_2 FILLER_73_1604 ();
 sg13g2_decap_8 FILLER_73_1624 ();
 sg13g2_decap_8 FILLER_73_1631 ();
 sg13g2_decap_8 FILLER_73_1638 ();
 sg13g2_decap_8 FILLER_73_1655 ();
 sg13g2_decap_8 FILLER_73_1662 ();
 sg13g2_decap_8 FILLER_73_1669 ();
 sg13g2_decap_8 FILLER_73_1676 ();
 sg13g2_decap_8 FILLER_73_1683 ();
 sg13g2_decap_8 FILLER_73_1690 ();
 sg13g2_decap_4 FILLER_73_1697 ();
 sg13g2_fill_2 FILLER_73_1701 ();
 sg13g2_fill_2 FILLER_73_1728 ();
 sg13g2_decap_8 FILLER_73_1743 ();
 sg13g2_decap_8 FILLER_73_1750 ();
 sg13g2_decap_8 FILLER_73_1757 ();
 sg13g2_decap_4 FILLER_73_1764 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_28 ();
 sg13g2_fill_2 FILLER_74_32 ();
 sg13g2_fill_2 FILLER_74_47 ();
 sg13g2_fill_2 FILLER_74_59 ();
 sg13g2_fill_1 FILLER_74_61 ();
 sg13g2_fill_2 FILLER_74_80 ();
 sg13g2_fill_1 FILLER_74_90 ();
 sg13g2_decap_8 FILLER_74_107 ();
 sg13g2_decap_8 FILLER_74_114 ();
 sg13g2_decap_8 FILLER_74_121 ();
 sg13g2_decap_8 FILLER_74_128 ();
 sg13g2_decap_8 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_142 ();
 sg13g2_decap_8 FILLER_74_149 ();
 sg13g2_decap_8 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_163 ();
 sg13g2_fill_1 FILLER_74_165 ();
 sg13g2_decap_4 FILLER_74_170 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_fill_1 FILLER_74_213 ();
 sg13g2_decap_8 FILLER_74_225 ();
 sg13g2_decap_8 FILLER_74_232 ();
 sg13g2_decap_8 FILLER_74_239 ();
 sg13g2_decap_8 FILLER_74_246 ();
 sg13g2_decap_8 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_260 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_2 FILLER_74_294 ();
 sg13g2_fill_1 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_4 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_360 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_decap_8 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_381 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_fill_2 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_406 ();
 sg13g2_decap_4 FILLER_74_412 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_4 FILLER_74_455 ();
 sg13g2_fill_2 FILLER_74_459 ();
 sg13g2_fill_2 FILLER_74_469 ();
 sg13g2_fill_1 FILLER_74_471 ();
 sg13g2_decap_8 FILLER_74_488 ();
 sg13g2_decap_8 FILLER_74_495 ();
 sg13g2_fill_2 FILLER_74_502 ();
 sg13g2_decap_8 FILLER_74_508 ();
 sg13g2_decap_8 FILLER_74_515 ();
 sg13g2_decap_8 FILLER_74_522 ();
 sg13g2_decap_8 FILLER_74_529 ();
 sg13g2_decap_8 FILLER_74_536 ();
 sg13g2_decap_8 FILLER_74_543 ();
 sg13g2_decap_8 FILLER_74_550 ();
 sg13g2_decap_4 FILLER_74_557 ();
 sg13g2_fill_1 FILLER_74_561 ();
 sg13g2_decap_8 FILLER_74_570 ();
 sg13g2_decap_8 FILLER_74_577 ();
 sg13g2_decap_8 FILLER_74_584 ();
 sg13g2_decap_8 FILLER_74_591 ();
 sg13g2_decap_8 FILLER_74_598 ();
 sg13g2_decap_4 FILLER_74_605 ();
 sg13g2_fill_2 FILLER_74_609 ();
 sg13g2_fill_1 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_625 ();
 sg13g2_decap_8 FILLER_74_632 ();
 sg13g2_decap_8 FILLER_74_639 ();
 sg13g2_decap_8 FILLER_74_646 ();
 sg13g2_decap_8 FILLER_74_653 ();
 sg13g2_decap_8 FILLER_74_660 ();
 sg13g2_decap_8 FILLER_74_667 ();
 sg13g2_decap_8 FILLER_74_674 ();
 sg13g2_decap_8 FILLER_74_681 ();
 sg13g2_decap_8 FILLER_74_688 ();
 sg13g2_decap_8 FILLER_74_695 ();
 sg13g2_decap_8 FILLER_74_702 ();
 sg13g2_decap_8 FILLER_74_709 ();
 sg13g2_decap_8 FILLER_74_716 ();
 sg13g2_decap_8 FILLER_74_723 ();
 sg13g2_decap_8 FILLER_74_730 ();
 sg13g2_decap_8 FILLER_74_737 ();
 sg13g2_decap_4 FILLER_74_744 ();
 sg13g2_fill_2 FILLER_74_748 ();
 sg13g2_fill_1 FILLER_74_765 ();
 sg13g2_fill_2 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_819 ();
 sg13g2_decap_4 FILLER_74_826 ();
 sg13g2_fill_2 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_fill_2 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_857 ();
 sg13g2_decap_8 FILLER_74_864 ();
 sg13g2_decap_8 FILLER_74_871 ();
 sg13g2_fill_2 FILLER_74_878 ();
 sg13g2_decap_4 FILLER_74_896 ();
 sg13g2_decap_8 FILLER_74_904 ();
 sg13g2_decap_8 FILLER_74_911 ();
 sg13g2_decap_8 FILLER_74_918 ();
 sg13g2_decap_4 FILLER_74_925 ();
 sg13g2_decap_4 FILLER_74_942 ();
 sg13g2_decap_4 FILLER_74_965 ();
 sg13g2_fill_1 FILLER_74_969 ();
 sg13g2_decap_8 FILLER_74_983 ();
 sg13g2_decap_8 FILLER_74_990 ();
 sg13g2_decap_8 FILLER_74_997 ();
 sg13g2_decap_8 FILLER_74_1004 ();
 sg13g2_decap_8 FILLER_74_1011 ();
 sg13g2_decap_4 FILLER_74_1018 ();
 sg13g2_fill_1 FILLER_74_1022 ();
 sg13g2_decap_4 FILLER_74_1046 ();
 sg13g2_decap_4 FILLER_74_1062 ();
 sg13g2_fill_2 FILLER_74_1066 ();
 sg13g2_decap_4 FILLER_74_1076 ();
 sg13g2_fill_1 FILLER_74_1080 ();
 sg13g2_decap_8 FILLER_74_1086 ();
 sg13g2_decap_8 FILLER_74_1093 ();
 sg13g2_decap_8 FILLER_74_1100 ();
 sg13g2_decap_4 FILLER_74_1107 ();
 sg13g2_decap_8 FILLER_74_1134 ();
 sg13g2_decap_8 FILLER_74_1141 ();
 sg13g2_fill_2 FILLER_74_1148 ();
 sg13g2_fill_1 FILLER_74_1150 ();
 sg13g2_decap_8 FILLER_74_1155 ();
 sg13g2_decap_8 FILLER_74_1172 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_decap_8 FILLER_74_1186 ();
 sg13g2_decap_8 FILLER_74_1193 ();
 sg13g2_decap_8 FILLER_74_1200 ();
 sg13g2_fill_1 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1218 ();
 sg13g2_decap_4 FILLER_74_1225 ();
 sg13g2_fill_2 FILLER_74_1229 ();
 sg13g2_decap_8 FILLER_74_1235 ();
 sg13g2_decap_8 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1249 ();
 sg13g2_decap_8 FILLER_74_1256 ();
 sg13g2_decap_8 FILLER_74_1263 ();
 sg13g2_decap_4 FILLER_74_1270 ();
 sg13g2_fill_2 FILLER_74_1274 ();
 sg13g2_decap_8 FILLER_74_1284 ();
 sg13g2_decap_8 FILLER_74_1291 ();
 sg13g2_fill_2 FILLER_74_1298 ();
 sg13g2_fill_1 FILLER_74_1300 ();
 sg13g2_decap_4 FILLER_74_1304 ();
 sg13g2_fill_2 FILLER_74_1308 ();
 sg13g2_fill_2 FILLER_74_1318 ();
 sg13g2_decap_8 FILLER_74_1338 ();
 sg13g2_decap_8 FILLER_74_1345 ();
 sg13g2_fill_2 FILLER_74_1352 ();
 sg13g2_decap_8 FILLER_74_1365 ();
 sg13g2_decap_8 FILLER_74_1372 ();
 sg13g2_decap_8 FILLER_74_1379 ();
 sg13g2_decap_4 FILLER_74_1386 ();
 sg13g2_fill_2 FILLER_74_1390 ();
 sg13g2_decap_8 FILLER_74_1418 ();
 sg13g2_decap_8 FILLER_74_1425 ();
 sg13g2_decap_8 FILLER_74_1432 ();
 sg13g2_fill_2 FILLER_74_1439 ();
 sg13g2_decap_8 FILLER_74_1454 ();
 sg13g2_fill_2 FILLER_74_1461 ();
 sg13g2_fill_1 FILLER_74_1463 ();
 sg13g2_decap_8 FILLER_74_1484 ();
 sg13g2_decap_4 FILLER_74_1491 ();
 sg13g2_fill_2 FILLER_74_1495 ();
 sg13g2_fill_2 FILLER_74_1510 ();
 sg13g2_decap_8 FILLER_74_1525 ();
 sg13g2_decap_8 FILLER_74_1532 ();
 sg13g2_decap_8 FILLER_74_1539 ();
 sg13g2_fill_1 FILLER_74_1546 ();
 sg13g2_fill_2 FILLER_74_1556 ();
 sg13g2_fill_1 FILLER_74_1558 ();
 sg13g2_decap_8 FILLER_74_1562 ();
 sg13g2_decap_8 FILLER_74_1569 ();
 sg13g2_decap_8 FILLER_74_1576 ();
 sg13g2_decap_8 FILLER_74_1583 ();
 sg13g2_decap_8 FILLER_74_1590 ();
 sg13g2_decap_8 FILLER_74_1597 ();
 sg13g2_decap_4 FILLER_74_1604 ();
 sg13g2_fill_2 FILLER_74_1608 ();
 sg13g2_decap_8 FILLER_74_1618 ();
 sg13g2_decap_8 FILLER_74_1625 ();
 sg13g2_decap_8 FILLER_74_1632 ();
 sg13g2_decap_8 FILLER_74_1639 ();
 sg13g2_fill_1 FILLER_74_1646 ();
 sg13g2_decap_8 FILLER_74_1673 ();
 sg13g2_decap_8 FILLER_74_1680 ();
 sg13g2_decap_8 FILLER_74_1687 ();
 sg13g2_decap_8 FILLER_74_1694 ();
 sg13g2_decap_8 FILLER_74_1701 ();
 sg13g2_fill_1 FILLER_74_1708 ();
 sg13g2_fill_2 FILLER_74_1719 ();
 sg13g2_fill_1 FILLER_74_1721 ();
 sg13g2_decap_8 FILLER_74_1748 ();
 sg13g2_decap_8 FILLER_74_1755 ();
 sg13g2_decap_4 FILLER_74_1762 ();
 sg13g2_fill_2 FILLER_74_1766 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_fill_2 FILLER_75_23 ();
 sg13g2_decap_4 FILLER_75_38 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_4 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_81 ();
 sg13g2_fill_1 FILLER_75_86 ();
 sg13g2_decap_8 FILLER_75_93 ();
 sg13g2_decap_8 FILLER_75_100 ();
 sg13g2_decap_8 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_decap_8 FILLER_75_121 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_135 ();
 sg13g2_decap_8 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_192 ();
 sg13g2_decap_8 FILLER_75_199 ();
 sg13g2_decap_8 FILLER_75_206 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_227 ();
 sg13g2_decap_8 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_241 ();
 sg13g2_decap_8 FILLER_75_248 ();
 sg13g2_decap_8 FILLER_75_255 ();
 sg13g2_decap_8 FILLER_75_262 ();
 sg13g2_decap_8 FILLER_75_269 ();
 sg13g2_decap_8 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_decap_8 FILLER_75_290 ();
 sg13g2_decap_8 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_316 ();
 sg13g2_fill_1 FILLER_75_318 ();
 sg13g2_fill_1 FILLER_75_330 ();
 sg13g2_decap_4 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_decap_8 FILLER_75_363 ();
 sg13g2_decap_8 FILLER_75_370 ();
 sg13g2_decap_4 FILLER_75_377 ();
 sg13g2_fill_1 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_414 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_8 FILLER_75_428 ();
 sg13g2_decap_8 FILLER_75_435 ();
 sg13g2_decap_8 FILLER_75_442 ();
 sg13g2_decap_8 FILLER_75_449 ();
 sg13g2_decap_8 FILLER_75_456 ();
 sg13g2_decap_8 FILLER_75_463 ();
 sg13g2_fill_2 FILLER_75_475 ();
 sg13g2_fill_1 FILLER_75_477 ();
 sg13g2_decap_8 FILLER_75_482 ();
 sg13g2_decap_8 FILLER_75_489 ();
 sg13g2_decap_8 FILLER_75_496 ();
 sg13g2_decap_8 FILLER_75_515 ();
 sg13g2_decap_8 FILLER_75_522 ();
 sg13g2_decap_4 FILLER_75_529 ();
 sg13g2_fill_2 FILLER_75_533 ();
 sg13g2_decap_8 FILLER_75_547 ();
 sg13g2_decap_4 FILLER_75_554 ();
 sg13g2_fill_2 FILLER_75_558 ();
 sg13g2_fill_2 FILLER_75_564 ();
 sg13g2_fill_1 FILLER_75_566 ();
 sg13g2_decap_4 FILLER_75_570 ();
 sg13g2_fill_2 FILLER_75_574 ();
 sg13g2_decap_8 FILLER_75_589 ();
 sg13g2_decap_4 FILLER_75_596 ();
 sg13g2_fill_2 FILLER_75_600 ();
 sg13g2_decap_8 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_633 ();
 sg13g2_decap_8 FILLER_75_640 ();
 sg13g2_decap_8 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_654 ();
 sg13g2_decap_8 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_668 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_decap_4 FILLER_75_682 ();
 sg13g2_fill_2 FILLER_75_686 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_fill_1 FILLER_75_760 ();
 sg13g2_fill_2 FILLER_75_764 ();
 sg13g2_fill_2 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_785 ();
 sg13g2_decap_8 FILLER_75_792 ();
 sg13g2_decap_4 FILLER_75_799 ();
 sg13g2_fill_1 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_809 ();
 sg13g2_decap_8 FILLER_75_816 ();
 sg13g2_decap_8 FILLER_75_823 ();
 sg13g2_decap_4 FILLER_75_838 ();
 sg13g2_fill_2 FILLER_75_842 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_decap_8 FILLER_75_855 ();
 sg13g2_decap_4 FILLER_75_862 ();
 sg13g2_decap_8 FILLER_75_892 ();
 sg13g2_decap_8 FILLER_75_899 ();
 sg13g2_decap_8 FILLER_75_906 ();
 sg13g2_fill_1 FILLER_75_913 ();
 sg13g2_fill_2 FILLER_75_922 ();
 sg13g2_fill_1 FILLER_75_924 ();
 sg13g2_decap_8 FILLER_75_930 ();
 sg13g2_decap_8 FILLER_75_937 ();
 sg13g2_decap_8 FILLER_75_944 ();
 sg13g2_decap_8 FILLER_75_951 ();
 sg13g2_decap_8 FILLER_75_958 ();
 sg13g2_decap_8 FILLER_75_965 ();
 sg13g2_decap_8 FILLER_75_972 ();
 sg13g2_decap_8 FILLER_75_979 ();
 sg13g2_decap_8 FILLER_75_986 ();
 sg13g2_decap_8 FILLER_75_993 ();
 sg13g2_decap_8 FILLER_75_1000 ();
 sg13g2_decap_8 FILLER_75_1007 ();
 sg13g2_fill_1 FILLER_75_1014 ();
 sg13g2_fill_2 FILLER_75_1028 ();
 sg13g2_decap_8 FILLER_75_1034 ();
 sg13g2_fill_2 FILLER_75_1041 ();
 sg13g2_fill_1 FILLER_75_1043 ();
 sg13g2_fill_1 FILLER_75_1049 ();
 sg13g2_decap_8 FILLER_75_1064 ();
 sg13g2_decap_8 FILLER_75_1071 ();
 sg13g2_decap_8 FILLER_75_1078 ();
 sg13g2_decap_8 FILLER_75_1085 ();
 sg13g2_decap_8 FILLER_75_1092 ();
 sg13g2_decap_8 FILLER_75_1099 ();
 sg13g2_decap_8 FILLER_75_1106 ();
 sg13g2_decap_8 FILLER_75_1113 ();
 sg13g2_decap_8 FILLER_75_1128 ();
 sg13g2_decap_8 FILLER_75_1135 ();
 sg13g2_decap_8 FILLER_75_1142 ();
 sg13g2_decap_8 FILLER_75_1149 ();
 sg13g2_fill_1 FILLER_75_1164 ();
 sg13g2_decap_8 FILLER_75_1171 ();
 sg13g2_decap_8 FILLER_75_1178 ();
 sg13g2_fill_1 FILLER_75_1185 ();
 sg13g2_decap_8 FILLER_75_1194 ();
 sg13g2_decap_8 FILLER_75_1201 ();
 sg13g2_fill_2 FILLER_75_1208 ();
 sg13g2_fill_1 FILLER_75_1210 ();
 sg13g2_decap_8 FILLER_75_1232 ();
 sg13g2_decap_8 FILLER_75_1239 ();
 sg13g2_decap_8 FILLER_75_1246 ();
 sg13g2_decap_8 FILLER_75_1253 ();
 sg13g2_decap_8 FILLER_75_1260 ();
 sg13g2_decap_8 FILLER_75_1267 ();
 sg13g2_fill_1 FILLER_75_1274 ();
 sg13g2_decap_8 FILLER_75_1278 ();
 sg13g2_decap_4 FILLER_75_1285 ();
 sg13g2_fill_2 FILLER_75_1292 ();
 sg13g2_fill_1 FILLER_75_1294 ();
 sg13g2_fill_1 FILLER_75_1300 ();
 sg13g2_decap_8 FILLER_75_1309 ();
 sg13g2_decap_8 FILLER_75_1316 ();
 sg13g2_decap_8 FILLER_75_1323 ();
 sg13g2_decap_4 FILLER_75_1330 ();
 sg13g2_fill_1 FILLER_75_1334 ();
 sg13g2_decap_8 FILLER_75_1348 ();
 sg13g2_decap_8 FILLER_75_1355 ();
 sg13g2_fill_2 FILLER_75_1362 ();
 sg13g2_fill_1 FILLER_75_1364 ();
 sg13g2_decap_8 FILLER_75_1370 ();
 sg13g2_decap_8 FILLER_75_1377 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_fill_1 FILLER_75_1413 ();
 sg13g2_decap_8 FILLER_75_1422 ();
 sg13g2_decap_8 FILLER_75_1429 ();
 sg13g2_decap_4 FILLER_75_1436 ();
 sg13g2_fill_2 FILLER_75_1440 ();
 sg13g2_decap_4 FILLER_75_1452 ();
 sg13g2_decap_8 FILLER_75_1468 ();
 sg13g2_decap_8 FILLER_75_1475 ();
 sg13g2_decap_4 FILLER_75_1482 ();
 sg13g2_fill_2 FILLER_75_1486 ();
 sg13g2_fill_1 FILLER_75_1499 ();
 sg13g2_decap_8 FILLER_75_1530 ();
 sg13g2_decap_8 FILLER_75_1537 ();
 sg13g2_decap_8 FILLER_75_1544 ();
 sg13g2_decap_4 FILLER_75_1551 ();
 sg13g2_decap_4 FILLER_75_1563 ();
 sg13g2_fill_1 FILLER_75_1567 ();
 sg13g2_decap_8 FILLER_75_1573 ();
 sg13g2_decap_8 FILLER_75_1580 ();
 sg13g2_decap_8 FILLER_75_1587 ();
 sg13g2_decap_8 FILLER_75_1594 ();
 sg13g2_decap_8 FILLER_75_1601 ();
 sg13g2_decap_8 FILLER_75_1608 ();
 sg13g2_decap_8 FILLER_75_1615 ();
 sg13g2_decap_8 FILLER_75_1622 ();
 sg13g2_decap_8 FILLER_75_1629 ();
 sg13g2_fill_1 FILLER_75_1636 ();
 sg13g2_fill_1 FILLER_75_1642 ();
 sg13g2_decap_4 FILLER_75_1652 ();
 sg13g2_fill_2 FILLER_75_1656 ();
 sg13g2_decap_8 FILLER_75_1662 ();
 sg13g2_decap_8 FILLER_75_1669 ();
 sg13g2_decap_8 FILLER_75_1676 ();
 sg13g2_decap_8 FILLER_75_1683 ();
 sg13g2_fill_1 FILLER_75_1690 ();
 sg13g2_decap_8 FILLER_75_1736 ();
 sg13g2_decap_8 FILLER_75_1743 ();
 sg13g2_decap_8 FILLER_75_1750 ();
 sg13g2_decap_8 FILLER_75_1757 ();
 sg13g2_decap_4 FILLER_75_1764 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_fill_2 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_31 ();
 sg13g2_fill_2 FILLER_76_38 ();
 sg13g2_fill_1 FILLER_76_40 ();
 sg13g2_fill_2 FILLER_76_57 ();
 sg13g2_decap_8 FILLER_76_69 ();
 sg13g2_decap_8 FILLER_76_76 ();
 sg13g2_decap_8 FILLER_76_83 ();
 sg13g2_decap_8 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_97 ();
 sg13g2_decap_8 FILLER_76_104 ();
 sg13g2_decap_8 FILLER_76_111 ();
 sg13g2_decap_8 FILLER_76_118 ();
 sg13g2_decap_8 FILLER_76_125 ();
 sg13g2_decap_8 FILLER_76_132 ();
 sg13g2_fill_2 FILLER_76_139 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_decap_8 FILLER_76_155 ();
 sg13g2_decap_8 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_169 ();
 sg13g2_decap_8 FILLER_76_176 ();
 sg13g2_decap_8 FILLER_76_183 ();
 sg13g2_decap_8 FILLER_76_190 ();
 sg13g2_decap_8 FILLER_76_197 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_8 FILLER_76_211 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_decap_8 FILLER_76_225 ();
 sg13g2_decap_8 FILLER_76_232 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_decap_4 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_257 ();
 sg13g2_decap_8 FILLER_76_267 ();
 sg13g2_decap_8 FILLER_76_274 ();
 sg13g2_decap_4 FILLER_76_281 ();
 sg13g2_fill_2 FILLER_76_285 ();
 sg13g2_decap_8 FILLER_76_291 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_decap_8 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_312 ();
 sg13g2_decap_4 FILLER_76_319 ();
 sg13g2_fill_1 FILLER_76_323 ();
 sg13g2_decap_8 FILLER_76_327 ();
 sg13g2_decap_8 FILLER_76_334 ();
 sg13g2_decap_8 FILLER_76_341 ();
 sg13g2_decap_8 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_76_355 ();
 sg13g2_decap_8 FILLER_76_362 ();
 sg13g2_fill_1 FILLER_76_369 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_389 ();
 sg13g2_fill_1 FILLER_76_391 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_decap_8 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_76_436 ();
 sg13g2_decap_8 FILLER_76_443 ();
 sg13g2_decap_8 FILLER_76_450 ();
 sg13g2_decap_8 FILLER_76_457 ();
 sg13g2_decap_4 FILLER_76_464 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_fill_2 FILLER_76_497 ();
 sg13g2_fill_1 FILLER_76_499 ();
 sg13g2_decap_8 FILLER_76_506 ();
 sg13g2_decap_8 FILLER_76_513 ();
 sg13g2_decap_8 FILLER_76_529 ();
 sg13g2_decap_8 FILLER_76_544 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_decap_8 FILLER_76_577 ();
 sg13g2_decap_8 FILLER_76_584 ();
 sg13g2_decap_8 FILLER_76_591 ();
 sg13g2_decap_4 FILLER_76_598 ();
 sg13g2_fill_1 FILLER_76_602 ();
 sg13g2_decap_8 FILLER_76_625 ();
 sg13g2_decap_4 FILLER_76_632 ();
 sg13g2_fill_2 FILLER_76_636 ();
 sg13g2_decap_4 FILLER_76_683 ();
 sg13g2_fill_1 FILLER_76_687 ();
 sg13g2_fill_2 FILLER_76_693 ();
 sg13g2_decap_4 FILLER_76_703 ();
 sg13g2_fill_2 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_741 ();
 sg13g2_fill_1 FILLER_76_743 ();
 sg13g2_fill_2 FILLER_76_759 ();
 sg13g2_fill_2 FILLER_76_764 ();
 sg13g2_fill_2 FILLER_76_769 ();
 sg13g2_decap_8 FILLER_76_790 ();
 sg13g2_decap_8 FILLER_76_797 ();
 sg13g2_decap_4 FILLER_76_819 ();
 sg13g2_fill_1 FILLER_76_823 ();
 sg13g2_fill_1 FILLER_76_850 ();
 sg13g2_decap_8 FILLER_76_859 ();
 sg13g2_decap_8 FILLER_76_866 ();
 sg13g2_decap_8 FILLER_76_873 ();
 sg13g2_decap_8 FILLER_76_880 ();
 sg13g2_decap_8 FILLER_76_887 ();
 sg13g2_decap_8 FILLER_76_894 ();
 sg13g2_decap_4 FILLER_76_901 ();
 sg13g2_fill_2 FILLER_76_905 ();
 sg13g2_fill_1 FILLER_76_931 ();
 sg13g2_decap_8 FILLER_76_940 ();
 sg13g2_decap_8 FILLER_76_947 ();
 sg13g2_decap_8 FILLER_76_967 ();
 sg13g2_decap_8 FILLER_76_974 ();
 sg13g2_decap_8 FILLER_76_981 ();
 sg13g2_decap_8 FILLER_76_988 ();
 sg13g2_decap_8 FILLER_76_995 ();
 sg13g2_decap_8 FILLER_76_1002 ();
 sg13g2_decap_4 FILLER_76_1030 ();
 sg13g2_fill_1 FILLER_76_1034 ();
 sg13g2_decap_8 FILLER_76_1039 ();
 sg13g2_decap_8 FILLER_76_1046 ();
 sg13g2_decap_8 FILLER_76_1053 ();
 sg13g2_fill_2 FILLER_76_1060 ();
 sg13g2_decap_8 FILLER_76_1067 ();
 sg13g2_decap_4 FILLER_76_1074 ();
 sg13g2_fill_1 FILLER_76_1078 ();
 sg13g2_decap_8 FILLER_76_1092 ();
 sg13g2_decap_8 FILLER_76_1099 ();
 sg13g2_decap_8 FILLER_76_1106 ();
 sg13g2_decap_8 FILLER_76_1113 ();
 sg13g2_decap_8 FILLER_76_1120 ();
 sg13g2_decap_8 FILLER_76_1127 ();
 sg13g2_decap_8 FILLER_76_1134 ();
 sg13g2_decap_8 FILLER_76_1141 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_fill_2 FILLER_76_1155 ();
 sg13g2_fill_1 FILLER_76_1157 ();
 sg13g2_decap_8 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1184 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_4 FILLER_76_1198 ();
 sg13g2_fill_2 FILLER_76_1210 ();
 sg13g2_fill_2 FILLER_76_1218 ();
 sg13g2_fill_1 FILLER_76_1220 ();
 sg13g2_decap_8 FILLER_76_1225 ();
 sg13g2_decap_8 FILLER_76_1232 ();
 sg13g2_decap_8 FILLER_76_1239 ();
 sg13g2_decap_8 FILLER_76_1246 ();
 sg13g2_decap_8 FILLER_76_1253 ();
 sg13g2_fill_2 FILLER_76_1260 ();
 sg13g2_fill_1 FILLER_76_1271 ();
 sg13g2_fill_1 FILLER_76_1275 ();
 sg13g2_decap_8 FILLER_76_1297 ();
 sg13g2_decap_8 FILLER_76_1304 ();
 sg13g2_decap_8 FILLER_76_1311 ();
 sg13g2_decap_8 FILLER_76_1318 ();
 sg13g2_decap_8 FILLER_76_1325 ();
 sg13g2_decap_8 FILLER_76_1332 ();
 sg13g2_fill_1 FILLER_76_1339 ();
 sg13g2_decap_8 FILLER_76_1345 ();
 sg13g2_decap_8 FILLER_76_1352 ();
 sg13g2_decap_8 FILLER_76_1359 ();
 sg13g2_decap_8 FILLER_76_1366 ();
 sg13g2_decap_8 FILLER_76_1373 ();
 sg13g2_decap_4 FILLER_76_1380 ();
 sg13g2_fill_2 FILLER_76_1384 ();
 sg13g2_decap_8 FILLER_76_1391 ();
 sg13g2_decap_8 FILLER_76_1418 ();
 sg13g2_decap_8 FILLER_76_1425 ();
 sg13g2_decap_8 FILLER_76_1432 ();
 sg13g2_decap_4 FILLER_76_1439 ();
 sg13g2_fill_1 FILLER_76_1443 ();
 sg13g2_decap_8 FILLER_76_1464 ();
 sg13g2_fill_2 FILLER_76_1471 ();
 sg13g2_fill_1 FILLER_76_1473 ();
 sg13g2_fill_1 FILLER_76_1487 ();
 sg13g2_decap_8 FILLER_76_1510 ();
 sg13g2_fill_1 FILLER_76_1517 ();
 sg13g2_decap_8 FILLER_76_1530 ();
 sg13g2_decap_8 FILLER_76_1537 ();
 sg13g2_decap_8 FILLER_76_1544 ();
 sg13g2_decap_8 FILLER_76_1551 ();
 sg13g2_decap_8 FILLER_76_1558 ();
 sg13g2_decap_8 FILLER_76_1565 ();
 sg13g2_decap_4 FILLER_76_1572 ();
 sg13g2_fill_2 FILLER_76_1576 ();
 sg13g2_decap_8 FILLER_76_1591 ();
 sg13g2_fill_1 FILLER_76_1598 ();
 sg13g2_decap_8 FILLER_76_1607 ();
 sg13g2_fill_1 FILLER_76_1614 ();
 sg13g2_decap_8 FILLER_76_1655 ();
 sg13g2_decap_8 FILLER_76_1662 ();
 sg13g2_decap_8 FILLER_76_1669 ();
 sg13g2_decap_8 FILLER_76_1676 ();
 sg13g2_decap_8 FILLER_76_1683 ();
 sg13g2_decap_8 FILLER_76_1690 ();
 sg13g2_decap_8 FILLER_76_1697 ();
 sg13g2_fill_2 FILLER_76_1704 ();
 sg13g2_decap_8 FILLER_76_1724 ();
 sg13g2_decap_8 FILLER_76_1731 ();
 sg13g2_decap_8 FILLER_76_1738 ();
 sg13g2_decap_8 FILLER_76_1745 ();
 sg13g2_decap_8 FILLER_76_1752 ();
 sg13g2_decap_8 FILLER_76_1759 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_fill_1 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_41 ();
 sg13g2_decap_8 FILLER_77_48 ();
 sg13g2_decap_8 FILLER_77_55 ();
 sg13g2_decap_8 FILLER_77_62 ();
 sg13g2_decap_8 FILLER_77_69 ();
 sg13g2_decap_8 FILLER_77_76 ();
 sg13g2_decap_8 FILLER_77_83 ();
 sg13g2_decap_8 FILLER_77_90 ();
 sg13g2_decap_8 FILLER_77_97 ();
 sg13g2_decap_8 FILLER_77_104 ();
 sg13g2_decap_8 FILLER_77_111 ();
 sg13g2_decap_8 FILLER_77_118 ();
 sg13g2_decap_8 FILLER_77_125 ();
 sg13g2_decap_4 FILLER_77_132 ();
 sg13g2_decap_8 FILLER_77_146 ();
 sg13g2_decap_8 FILLER_77_153 ();
 sg13g2_decap_8 FILLER_77_160 ();
 sg13g2_decap_8 FILLER_77_167 ();
 sg13g2_decap_8 FILLER_77_174 ();
 sg13g2_decap_8 FILLER_77_181 ();
 sg13g2_decap_8 FILLER_77_188 ();
 sg13g2_fill_2 FILLER_77_195 ();
 sg13g2_fill_1 FILLER_77_197 ();
 sg13g2_decap_4 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_decap_8 FILLER_77_251 ();
 sg13g2_decap_8 FILLER_77_258 ();
 sg13g2_decap_8 FILLER_77_265 ();
 sg13g2_decap_8 FILLER_77_272 ();
 sg13g2_decap_8 FILLER_77_279 ();
 sg13g2_decap_8 FILLER_77_286 ();
 sg13g2_decap_8 FILLER_77_293 ();
 sg13g2_decap_8 FILLER_77_300 ();
 sg13g2_decap_4 FILLER_77_307 ();
 sg13g2_fill_1 FILLER_77_311 ();
 sg13g2_decap_8 FILLER_77_320 ();
 sg13g2_decap_8 FILLER_77_327 ();
 sg13g2_decap_8 FILLER_77_334 ();
 sg13g2_decap_4 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_365 ();
 sg13g2_fill_2 FILLER_77_372 ();
 sg13g2_fill_1 FILLER_77_374 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_461 ();
 sg13g2_fill_2 FILLER_77_468 ();
 sg13g2_fill_1 FILLER_77_470 ();
 sg13g2_decap_8 FILLER_77_479 ();
 sg13g2_decap_4 FILLER_77_486 ();
 sg13g2_decap_8 FILLER_77_516 ();
 sg13g2_decap_8 FILLER_77_523 ();
 sg13g2_decap_8 FILLER_77_530 ();
 sg13g2_decap_8 FILLER_77_537 ();
 sg13g2_decap_8 FILLER_77_544 ();
 sg13g2_decap_4 FILLER_77_551 ();
 sg13g2_fill_1 FILLER_77_555 ();
 sg13g2_fill_2 FILLER_77_564 ();
 sg13g2_fill_1 FILLER_77_566 ();
 sg13g2_decap_8 FILLER_77_572 ();
 sg13g2_decap_8 FILLER_77_579 ();
 sg13g2_decap_8 FILLER_77_586 ();
 sg13g2_decap_8 FILLER_77_593 ();
 sg13g2_decap_8 FILLER_77_600 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_fill_2 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_8 FILLER_77_639 ();
 sg13g2_decap_8 FILLER_77_646 ();
 sg13g2_decap_4 FILLER_77_653 ();
 sg13g2_fill_2 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_663 ();
 sg13g2_decap_4 FILLER_77_670 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_4 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_decap_4 FILLER_77_739 ();
 sg13g2_fill_1 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_794 ();
 sg13g2_decap_4 FILLER_77_801 ();
 sg13g2_fill_2 FILLER_77_805 ();
 sg13g2_fill_1 FILLER_77_853 ();
 sg13g2_decap_8 FILLER_77_862 ();
 sg13g2_decap_8 FILLER_77_869 ();
 sg13g2_decap_8 FILLER_77_876 ();
 sg13g2_decap_8 FILLER_77_883 ();
 sg13g2_decap_8 FILLER_77_890 ();
 sg13g2_decap_8 FILLER_77_897 ();
 sg13g2_fill_2 FILLER_77_904 ();
 sg13g2_decap_8 FILLER_77_919 ();
 sg13g2_fill_1 FILLER_77_926 ();
 sg13g2_decap_8 FILLER_77_940 ();
 sg13g2_decap_4 FILLER_77_947 ();
 sg13g2_fill_1 FILLER_77_951 ();
 sg13g2_decap_8 FILLER_77_978 ();
 sg13g2_decap_8 FILLER_77_985 ();
 sg13g2_decap_8 FILLER_77_992 ();
 sg13g2_fill_1 FILLER_77_999 ();
 sg13g2_decap_8 FILLER_77_1033 ();
 sg13g2_decap_8 FILLER_77_1040 ();
 sg13g2_decap_4 FILLER_77_1047 ();
 sg13g2_fill_2 FILLER_77_1051 ();
 sg13g2_fill_2 FILLER_77_1079 ();
 sg13g2_fill_1 FILLER_77_1087 ();
 sg13g2_decap_4 FILLER_77_1091 ();
 sg13g2_decap_4 FILLER_77_1101 ();
 sg13g2_fill_2 FILLER_77_1105 ();
 sg13g2_fill_2 FILLER_77_1112 ();
 sg13g2_decap_8 FILLER_77_1122 ();
 sg13g2_decap_8 FILLER_77_1137 ();
 sg13g2_decap_8 FILLER_77_1144 ();
 sg13g2_decap_8 FILLER_77_1177 ();
 sg13g2_decap_8 FILLER_77_1184 ();
 sg13g2_decap_8 FILLER_77_1191 ();
 sg13g2_decap_8 FILLER_77_1198 ();
 sg13g2_decap_4 FILLER_77_1205 ();
 sg13g2_fill_2 FILLER_77_1209 ();
 sg13g2_decap_8 FILLER_77_1220 ();
 sg13g2_decap_8 FILLER_77_1227 ();
 sg13g2_fill_1 FILLER_77_1234 ();
 sg13g2_decap_8 FILLER_77_1245 ();
 sg13g2_decap_8 FILLER_77_1252 ();
 sg13g2_fill_1 FILLER_77_1268 ();
 sg13g2_decap_8 FILLER_77_1302 ();
 sg13g2_decap_8 FILLER_77_1309 ();
 sg13g2_decap_8 FILLER_77_1316 ();
 sg13g2_decap_8 FILLER_77_1323 ();
 sg13g2_decap_8 FILLER_77_1330 ();
 sg13g2_decap_4 FILLER_77_1337 ();
 sg13g2_fill_1 FILLER_77_1341 ();
 sg13g2_decap_8 FILLER_77_1350 ();
 sg13g2_fill_2 FILLER_77_1357 ();
 sg13g2_decap_8 FILLER_77_1365 ();
 sg13g2_decap_8 FILLER_77_1372 ();
 sg13g2_fill_2 FILLER_77_1379 ();
 sg13g2_decap_8 FILLER_77_1384 ();
 sg13g2_decap_8 FILLER_77_1391 ();
 sg13g2_decap_8 FILLER_77_1398 ();
 sg13g2_decap_8 FILLER_77_1405 ();
 sg13g2_decap_8 FILLER_77_1412 ();
 sg13g2_decap_8 FILLER_77_1419 ();
 sg13g2_decap_8 FILLER_77_1426 ();
 sg13g2_decap_4 FILLER_77_1433 ();
 sg13g2_fill_2 FILLER_77_1437 ();
 sg13g2_fill_1 FILLER_77_1447 ();
 sg13g2_fill_1 FILLER_77_1452 ();
 sg13g2_decap_8 FILLER_77_1457 ();
 sg13g2_decap_8 FILLER_77_1464 ();
 sg13g2_decap_8 FILLER_77_1471 ();
 sg13g2_decap_8 FILLER_77_1478 ();
 sg13g2_decap_8 FILLER_77_1485 ();
 sg13g2_fill_1 FILLER_77_1492 ();
 sg13g2_decap_8 FILLER_77_1496 ();
 sg13g2_fill_2 FILLER_77_1503 ();
 sg13g2_decap_8 FILLER_77_1513 ();
 sg13g2_decap_8 FILLER_77_1520 ();
 sg13g2_decap_8 FILLER_77_1527 ();
 sg13g2_decap_8 FILLER_77_1534 ();
 sg13g2_decap_8 FILLER_77_1541 ();
 sg13g2_decap_8 FILLER_77_1548 ();
 sg13g2_decap_8 FILLER_77_1555 ();
 sg13g2_fill_2 FILLER_77_1562 ();
 sg13g2_decap_8 FILLER_77_1571 ();
 sg13g2_decap_8 FILLER_77_1578 ();
 sg13g2_decap_8 FILLER_77_1585 ();
 sg13g2_decap_8 FILLER_77_1592 ();
 sg13g2_decap_8 FILLER_77_1599 ();
 sg13g2_fill_2 FILLER_77_1606 ();
 sg13g2_fill_1 FILLER_77_1608 ();
 sg13g2_decap_4 FILLER_77_1622 ();
 sg13g2_decap_8 FILLER_77_1643 ();
 sg13g2_decap_8 FILLER_77_1650 ();
 sg13g2_decap_8 FILLER_77_1657 ();
 sg13g2_decap_8 FILLER_77_1664 ();
 sg13g2_decap_8 FILLER_77_1671 ();
 sg13g2_decap_8 FILLER_77_1678 ();
 sg13g2_decap_8 FILLER_77_1685 ();
 sg13g2_decap_8 FILLER_77_1692 ();
 sg13g2_decap_8 FILLER_77_1699 ();
 sg13g2_decap_8 FILLER_77_1706 ();
 sg13g2_decap_4 FILLER_77_1713 ();
 sg13g2_fill_1 FILLER_77_1717 ();
 sg13g2_decap_8 FILLER_77_1722 ();
 sg13g2_decap_8 FILLER_77_1729 ();
 sg13g2_decap_8 FILLER_77_1736 ();
 sg13g2_decap_8 FILLER_77_1743 ();
 sg13g2_decap_8 FILLER_77_1750 ();
 sg13g2_decap_8 FILLER_77_1757 ();
 sg13g2_decap_4 FILLER_77_1764 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_4 FILLER_78_14 ();
 sg13g2_fill_1 FILLER_78_18 ();
 sg13g2_fill_1 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_50 ();
 sg13g2_decap_8 FILLER_78_57 ();
 sg13g2_decap_8 FILLER_78_64 ();
 sg13g2_decap_8 FILLER_78_71 ();
 sg13g2_decap_8 FILLER_78_78 ();
 sg13g2_fill_1 FILLER_78_85 ();
 sg13g2_decap_8 FILLER_78_103 ();
 sg13g2_decap_8 FILLER_78_114 ();
 sg13g2_fill_2 FILLER_78_121 ();
 sg13g2_fill_1 FILLER_78_123 ();
 sg13g2_decap_8 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_136 ();
 sg13g2_decap_8 FILLER_78_155 ();
 sg13g2_fill_1 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_171 ();
 sg13g2_decap_8 FILLER_78_178 ();
 sg13g2_decap_8 FILLER_78_185 ();
 sg13g2_decap_8 FILLER_78_192 ();
 sg13g2_decap_8 FILLER_78_199 ();
 sg13g2_decap_8 FILLER_78_206 ();
 sg13g2_decap_4 FILLER_78_213 ();
 sg13g2_decap_8 FILLER_78_228 ();
 sg13g2_fill_1 FILLER_78_235 ();
 sg13g2_decap_4 FILLER_78_246 ();
 sg13g2_fill_1 FILLER_78_250 ();
 sg13g2_fill_1 FILLER_78_283 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_decap_4 FILLER_78_303 ();
 sg13g2_fill_2 FILLER_78_307 ();
 sg13g2_fill_1 FILLER_78_313 ();
 sg13g2_decap_8 FILLER_78_318 ();
 sg13g2_decap_8 FILLER_78_325 ();
 sg13g2_decap_8 FILLER_78_332 ();
 sg13g2_fill_1 FILLER_78_339 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_4 FILLER_78_417 ();
 sg13g2_fill_1 FILLER_78_421 ();
 sg13g2_fill_1 FILLER_78_451 ();
 sg13g2_decap_8 FILLER_78_460 ();
 sg13g2_fill_2 FILLER_78_467 ();
 sg13g2_fill_1 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_474 ();
 sg13g2_decap_8 FILLER_78_481 ();
 sg13g2_decap_8 FILLER_78_488 ();
 sg13g2_fill_2 FILLER_78_495 ();
 sg13g2_decap_8 FILLER_78_520 ();
 sg13g2_decap_8 FILLER_78_527 ();
 sg13g2_decap_8 FILLER_78_534 ();
 sg13g2_decap_8 FILLER_78_541 ();
 sg13g2_fill_2 FILLER_78_548 ();
 sg13g2_decap_4 FILLER_78_558 ();
 sg13g2_fill_2 FILLER_78_562 ();
 sg13g2_decap_8 FILLER_78_572 ();
 sg13g2_decap_8 FILLER_78_579 ();
 sg13g2_decap_8 FILLER_78_586 ();
 sg13g2_decap_8 FILLER_78_593 ();
 sg13g2_decap_8 FILLER_78_600 ();
 sg13g2_decap_8 FILLER_78_607 ();
 sg13g2_decap_4 FILLER_78_614 ();
 sg13g2_decap_4 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_648 ();
 sg13g2_decap_8 FILLER_78_655 ();
 sg13g2_decap_8 FILLER_78_662 ();
 sg13g2_decap_8 FILLER_78_669 ();
 sg13g2_decap_4 FILLER_78_676 ();
 sg13g2_decap_4 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_702 ();
 sg13g2_fill_1 FILLER_78_709 ();
 sg13g2_decap_8 FILLER_78_723 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_decap_8 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_744 ();
 sg13g2_decap_4 FILLER_78_751 ();
 sg13g2_fill_2 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_fill_1 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_8 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_decap_8 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_78_867 ();
 sg13g2_decap_8 FILLER_78_874 ();
 sg13g2_decap_8 FILLER_78_881 ();
 sg13g2_decap_8 FILLER_78_888 ();
 sg13g2_decap_8 FILLER_78_895 ();
 sg13g2_fill_1 FILLER_78_902 ();
 sg13g2_decap_8 FILLER_78_916 ();
 sg13g2_decap_8 FILLER_78_923 ();
 sg13g2_decap_8 FILLER_78_930 ();
 sg13g2_decap_8 FILLER_78_937 ();
 sg13g2_decap_8 FILLER_78_950 ();
 sg13g2_decap_4 FILLER_78_957 ();
 sg13g2_fill_1 FILLER_78_961 ();
 sg13g2_decap_8 FILLER_78_966 ();
 sg13g2_decap_8 FILLER_78_973 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_fill_2 FILLER_78_987 ();
 sg13g2_decap_8 FILLER_78_1002 ();
 sg13g2_fill_2 FILLER_78_1009 ();
 sg13g2_decap_8 FILLER_78_1028 ();
 sg13g2_decap_8 FILLER_78_1035 ();
 sg13g2_decap_8 FILLER_78_1042 ();
 sg13g2_decap_8 FILLER_78_1049 ();
 sg13g2_decap_8 FILLER_78_1056 ();
 sg13g2_decap_8 FILLER_78_1063 ();
 sg13g2_decap_8 FILLER_78_1070 ();
 sg13g2_decap_8 FILLER_78_1077 ();
 sg13g2_decap_4 FILLER_78_1084 ();
 sg13g2_fill_1 FILLER_78_1102 ();
 sg13g2_decap_8 FILLER_78_1124 ();
 sg13g2_decap_8 FILLER_78_1131 ();
 sg13g2_decap_8 FILLER_78_1138 ();
 sg13g2_decap_8 FILLER_78_1145 ();
 sg13g2_decap_8 FILLER_78_1152 ();
 sg13g2_fill_2 FILLER_78_1159 ();
 sg13g2_fill_1 FILLER_78_1161 ();
 sg13g2_fill_2 FILLER_78_1166 ();
 sg13g2_fill_1 FILLER_78_1168 ();
 sg13g2_decap_8 FILLER_78_1174 ();
 sg13g2_decap_8 FILLER_78_1181 ();
 sg13g2_decap_8 FILLER_78_1188 ();
 sg13g2_decap_8 FILLER_78_1195 ();
 sg13g2_fill_2 FILLER_78_1202 ();
 sg13g2_fill_1 FILLER_78_1204 ();
 sg13g2_fill_2 FILLER_78_1209 ();
 sg13g2_fill_1 FILLER_78_1211 ();
 sg13g2_decap_8 FILLER_78_1225 ();
 sg13g2_decap_8 FILLER_78_1245 ();
 sg13g2_decap_8 FILLER_78_1252 ();
 sg13g2_fill_1 FILLER_78_1274 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_8 FILLER_78_1310 ();
 sg13g2_decap_8 FILLER_78_1317 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_fill_1 FILLER_78_1326 ();
 sg13g2_decap_4 FILLER_78_1330 ();
 sg13g2_fill_1 FILLER_78_1334 ();
 sg13g2_decap_8 FILLER_78_1364 ();
 sg13g2_decap_8 FILLER_78_1371 ();
 sg13g2_fill_2 FILLER_78_1385 ();
 sg13g2_decap_8 FILLER_78_1408 ();
 sg13g2_decap_8 FILLER_78_1415 ();
 sg13g2_decap_8 FILLER_78_1422 ();
 sg13g2_decap_8 FILLER_78_1429 ();
 sg13g2_decap_8 FILLER_78_1436 ();
 sg13g2_decap_8 FILLER_78_1443 ();
 sg13g2_decap_8 FILLER_78_1450 ();
 sg13g2_decap_8 FILLER_78_1457 ();
 sg13g2_decap_8 FILLER_78_1464 ();
 sg13g2_decap_8 FILLER_78_1471 ();
 sg13g2_decap_8 FILLER_78_1478 ();
 sg13g2_decap_8 FILLER_78_1485 ();
 sg13g2_fill_1 FILLER_78_1492 ();
 sg13g2_decap_8 FILLER_78_1498 ();
 sg13g2_decap_8 FILLER_78_1505 ();
 sg13g2_decap_8 FILLER_78_1512 ();
 sg13g2_decap_8 FILLER_78_1519 ();
 sg13g2_decap_8 FILLER_78_1526 ();
 sg13g2_decap_8 FILLER_78_1533 ();
 sg13g2_decap_4 FILLER_78_1540 ();
 sg13g2_fill_2 FILLER_78_1544 ();
 sg13g2_decap_8 FILLER_78_1585 ();
 sg13g2_decap_4 FILLER_78_1592 ();
 sg13g2_fill_2 FILLER_78_1596 ();
 sg13g2_decap_8 FILLER_78_1603 ();
 sg13g2_decap_8 FILLER_78_1610 ();
 sg13g2_decap_8 FILLER_78_1617 ();
 sg13g2_decap_8 FILLER_78_1624 ();
 sg13g2_decap_4 FILLER_78_1631 ();
 sg13g2_fill_1 FILLER_78_1635 ();
 sg13g2_fill_2 FILLER_78_1647 ();
 sg13g2_decap_8 FILLER_78_1674 ();
 sg13g2_decap_4 FILLER_78_1681 ();
 sg13g2_fill_1 FILLER_78_1685 ();
 sg13g2_decap_8 FILLER_78_1696 ();
 sg13g2_decap_4 FILLER_78_1703 ();
 sg13g2_decap_8 FILLER_78_1746 ();
 sg13g2_decap_8 FILLER_78_1753 ();
 sg13g2_decap_8 FILLER_78_1760 ();
 sg13g2_fill_1 FILLER_78_1767 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_47 ();
 sg13g2_decap_8 FILLER_79_54 ();
 sg13g2_decap_8 FILLER_79_61 ();
 sg13g2_decap_8 FILLER_79_68 ();
 sg13g2_decap_8 FILLER_79_75 ();
 sg13g2_decap_8 FILLER_79_82 ();
 sg13g2_decap_8 FILLER_79_89 ();
 sg13g2_decap_4 FILLER_79_96 ();
 sg13g2_fill_2 FILLER_79_114 ();
 sg13g2_fill_1 FILLER_79_116 ();
 sg13g2_decap_8 FILLER_79_130 ();
 sg13g2_decap_4 FILLER_79_137 ();
 sg13g2_fill_2 FILLER_79_141 ();
 sg13g2_fill_2 FILLER_79_151 ();
 sg13g2_fill_1 FILLER_79_153 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_fill_1 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_180 ();
 sg13g2_fill_2 FILLER_79_187 ();
 sg13g2_decap_8 FILLER_79_194 ();
 sg13g2_decap_8 FILLER_79_201 ();
 sg13g2_decap_8 FILLER_79_208 ();
 sg13g2_decap_8 FILLER_79_215 ();
 sg13g2_decap_4 FILLER_79_222 ();
 sg13g2_fill_1 FILLER_79_226 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_2 FILLER_79_258 ();
 sg13g2_fill_1 FILLER_79_260 ();
 sg13g2_fill_2 FILLER_79_265 ();
 sg13g2_decap_8 FILLER_79_271 ();
 sg13g2_fill_1 FILLER_79_278 ();
 sg13g2_decap_8 FILLER_79_300 ();
 sg13g2_decap_8 FILLER_79_307 ();
 sg13g2_decap_4 FILLER_79_314 ();
 sg13g2_fill_2 FILLER_79_318 ();
 sg13g2_decap_8 FILLER_79_328 ();
 sg13g2_decap_4 FILLER_79_335 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_4 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_8 FILLER_79_403 ();
 sg13g2_decap_8 FILLER_79_410 ();
 sg13g2_decap_4 FILLER_79_417 ();
 sg13g2_decap_4 FILLER_79_436 ();
 sg13g2_decap_8 FILLER_79_460 ();
 sg13g2_decap_8 FILLER_79_467 ();
 sg13g2_decap_8 FILLER_79_474 ();
 sg13g2_decap_4 FILLER_79_481 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_fill_2 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_514 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_535 ();
 sg13g2_fill_2 FILLER_79_542 ();
 sg13g2_decap_8 FILLER_79_554 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_8 FILLER_79_575 ();
 sg13g2_decap_8 FILLER_79_582 ();
 sg13g2_fill_2 FILLER_79_589 ();
 sg13g2_decap_8 FILLER_79_603 ();
 sg13g2_fill_1 FILLER_79_619 ();
 sg13g2_decap_4 FILLER_79_628 ();
 sg13g2_decap_8 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_8 FILLER_79_696 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_4 FILLER_79_717 ();
 sg13g2_decap_4 FILLER_79_734 ();
 sg13g2_fill_2 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_fill_2 FILLER_79_764 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_fill_2 FILLER_79_862 ();
 sg13g2_fill_1 FILLER_79_864 ();
 sg13g2_decap_4 FILLER_79_873 ();
 sg13g2_fill_2 FILLER_79_877 ();
 sg13g2_decap_8 FILLER_79_884 ();
 sg13g2_decap_8 FILLER_79_891 ();
 sg13g2_decap_8 FILLER_79_898 ();
 sg13g2_decap_8 FILLER_79_905 ();
 sg13g2_decap_8 FILLER_79_912 ();
 sg13g2_decap_8 FILLER_79_919 ();
 sg13g2_decap_8 FILLER_79_926 ();
 sg13g2_decap_8 FILLER_79_933 ();
 sg13g2_decap_8 FILLER_79_940 ();
 sg13g2_decap_8 FILLER_79_947 ();
 sg13g2_decap_8 FILLER_79_954 ();
 sg13g2_decap_8 FILLER_79_961 ();
 sg13g2_decap_8 FILLER_79_968 ();
 sg13g2_decap_8 FILLER_79_975 ();
 sg13g2_decap_8 FILLER_79_982 ();
 sg13g2_decap_8 FILLER_79_989 ();
 sg13g2_decap_8 FILLER_79_996 ();
 sg13g2_decap_8 FILLER_79_1003 ();
 sg13g2_decap_4 FILLER_79_1010 ();
 sg13g2_fill_2 FILLER_79_1014 ();
 sg13g2_decap_8 FILLER_79_1024 ();
 sg13g2_decap_8 FILLER_79_1031 ();
 sg13g2_decap_8 FILLER_79_1038 ();
 sg13g2_decap_8 FILLER_79_1045 ();
 sg13g2_decap_8 FILLER_79_1052 ();
 sg13g2_decap_8 FILLER_79_1059 ();
 sg13g2_decap_8 FILLER_79_1066 ();
 sg13g2_decap_8 FILLER_79_1073 ();
 sg13g2_decap_8 FILLER_79_1080 ();
 sg13g2_decap_8 FILLER_79_1087 ();
 sg13g2_decap_4 FILLER_79_1094 ();
 sg13g2_fill_2 FILLER_79_1098 ();
 sg13g2_decap_8 FILLER_79_1106 ();
 sg13g2_decap_8 FILLER_79_1113 ();
 sg13g2_decap_8 FILLER_79_1120 ();
 sg13g2_decap_8 FILLER_79_1127 ();
 sg13g2_decap_8 FILLER_79_1134 ();
 sg13g2_decap_8 FILLER_79_1141 ();
 sg13g2_decap_4 FILLER_79_1148 ();
 sg13g2_decap_8 FILLER_79_1165 ();
 sg13g2_decap_8 FILLER_79_1172 ();
 sg13g2_decap_8 FILLER_79_1179 ();
 sg13g2_decap_8 FILLER_79_1186 ();
 sg13g2_fill_2 FILLER_79_1197 ();
 sg13g2_fill_1 FILLER_79_1209 ();
 sg13g2_decap_8 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1225 ();
 sg13g2_decap_8 FILLER_79_1232 ();
 sg13g2_fill_2 FILLER_79_1239 ();
 sg13g2_fill_2 FILLER_79_1276 ();
 sg13g2_fill_1 FILLER_79_1287 ();
 sg13g2_decap_8 FILLER_79_1292 ();
 sg13g2_decap_8 FILLER_79_1299 ();
 sg13g2_decap_8 FILLER_79_1306 ();
 sg13g2_decap_8 FILLER_79_1313 ();
 sg13g2_decap_8 FILLER_79_1320 ();
 sg13g2_decap_8 FILLER_79_1369 ();
 sg13g2_decap_4 FILLER_79_1376 ();
 sg13g2_fill_1 FILLER_79_1380 ();
 sg13g2_fill_2 FILLER_79_1384 ();
 sg13g2_fill_1 FILLER_79_1386 ();
 sg13g2_decap_8 FILLER_79_1391 ();
 sg13g2_decap_8 FILLER_79_1398 ();
 sg13g2_decap_8 FILLER_79_1405 ();
 sg13g2_decap_8 FILLER_79_1412 ();
 sg13g2_decap_8 FILLER_79_1419 ();
 sg13g2_decap_8 FILLER_79_1426 ();
 sg13g2_decap_8 FILLER_79_1433 ();
 sg13g2_decap_8 FILLER_79_1440 ();
 sg13g2_decap_8 FILLER_79_1447 ();
 sg13g2_decap_8 FILLER_79_1454 ();
 sg13g2_decap_8 FILLER_79_1461 ();
 sg13g2_decap_8 FILLER_79_1468 ();
 sg13g2_decap_8 FILLER_79_1475 ();
 sg13g2_decap_8 FILLER_79_1482 ();
 sg13g2_decap_8 FILLER_79_1489 ();
 sg13g2_decap_8 FILLER_79_1517 ();
 sg13g2_decap_8 FILLER_79_1524 ();
 sg13g2_decap_8 FILLER_79_1531 ();
 sg13g2_decap_8 FILLER_79_1538 ();
 sg13g2_decap_8 FILLER_79_1545 ();
 sg13g2_decap_4 FILLER_79_1552 ();
 sg13g2_fill_1 FILLER_79_1556 ();
 sg13g2_decap_8 FILLER_79_1561 ();
 sg13g2_decap_8 FILLER_79_1568 ();
 sg13g2_decap_8 FILLER_79_1575 ();
 sg13g2_decap_8 FILLER_79_1582 ();
 sg13g2_decap_4 FILLER_79_1589 ();
 sg13g2_decap_4 FILLER_79_1603 ();
 sg13g2_fill_1 FILLER_79_1607 ();
 sg13g2_decap_8 FILLER_79_1621 ();
 sg13g2_decap_8 FILLER_79_1628 ();
 sg13g2_decap_8 FILLER_79_1635 ();
 sg13g2_decap_4 FILLER_79_1642 ();
 sg13g2_fill_2 FILLER_79_1646 ();
 sg13g2_decap_8 FILLER_79_1674 ();
 sg13g2_decap_8 FILLER_79_1681 ();
 sg13g2_fill_1 FILLER_79_1688 ();
 sg13g2_decap_8 FILLER_79_1702 ();
 sg13g2_decap_8 FILLER_79_1709 ();
 sg13g2_decap_8 FILLER_79_1716 ();
 sg13g2_decap_8 FILLER_79_1723 ();
 sg13g2_decap_8 FILLER_79_1730 ();
 sg13g2_decap_4 FILLER_79_1737 ();
 sg13g2_fill_2 FILLER_79_1741 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_21 ();
 sg13g2_fill_1 FILLER_80_27 ();
 sg13g2_decap_8 FILLER_80_36 ();
 sg13g2_decap_8 FILLER_80_43 ();
 sg13g2_decap_8 FILLER_80_50 ();
 sg13g2_decap_8 FILLER_80_57 ();
 sg13g2_decap_8 FILLER_80_76 ();
 sg13g2_decap_8 FILLER_80_83 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_1 FILLER_80_92 ();
 sg13g2_decap_8 FILLER_80_104 ();
 sg13g2_decap_8 FILLER_80_111 ();
 sg13g2_decap_8 FILLER_80_118 ();
 sg13g2_decap_8 FILLER_80_125 ();
 sg13g2_decap_8 FILLER_80_132 ();
 sg13g2_decap_8 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_decap_8 FILLER_80_153 ();
 sg13g2_decap_4 FILLER_80_160 ();
 sg13g2_fill_1 FILLER_80_164 ();
 sg13g2_fill_2 FILLER_80_173 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_decap_4 FILLER_80_179 ();
 sg13g2_fill_2 FILLER_80_183 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_fill_2 FILLER_80_221 ();
 sg13g2_fill_1 FILLER_80_240 ();
 sg13g2_decap_8 FILLER_80_246 ();
 sg13g2_decap_8 FILLER_80_253 ();
 sg13g2_decap_8 FILLER_80_260 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_decap_4 FILLER_80_281 ();
 sg13g2_fill_2 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_4 FILLER_80_354 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_4 FILLER_80_378 ();
 sg13g2_fill_1 FILLER_80_382 ();
 sg13g2_fill_1 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_415 ();
 sg13g2_fill_2 FILLER_80_422 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_fill_2 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_463 ();
 sg13g2_decap_8 FILLER_80_470 ();
 sg13g2_decap_8 FILLER_80_477 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_491 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_4 FILLER_80_554 ();
 sg13g2_fill_2 FILLER_80_562 ();
 sg13g2_decap_8 FILLER_80_579 ();
 sg13g2_decap_4 FILLER_80_586 ();
 sg13g2_fill_1 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_fill_1 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_4 FILLER_80_651 ();
 sg13g2_fill_2 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_fill_2 FILLER_80_669 ();
 sg13g2_fill_1 FILLER_80_671 ();
 sg13g2_fill_1 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_fill_1 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_731 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_fill_2 FILLER_80_769 ();
 sg13g2_fill_1 FILLER_80_771 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_fill_1 FILLER_80_818 ();
 sg13g2_decap_4 FILLER_80_828 ();
 sg13g2_fill_1 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_fill_2 FILLER_80_844 ();
 sg13g2_fill_1 FILLER_80_846 ();
 sg13g2_fill_1 FILLER_80_861 ();
 sg13g2_decap_4 FILLER_80_888 ();
 sg13g2_decap_8 FILLER_80_905 ();
 sg13g2_decap_8 FILLER_80_912 ();
 sg13g2_decap_8 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_4 FILLER_80_933 ();
 sg13g2_fill_2 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_4 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_fill_2 FILLER_80_1003 ();
 sg13g2_fill_1 FILLER_80_1005 ();
 sg13g2_decap_8 FILLER_80_1014 ();
 sg13g2_decap_8 FILLER_80_1021 ();
 sg13g2_decap_8 FILLER_80_1028 ();
 sg13g2_decap_8 FILLER_80_1035 ();
 sg13g2_decap_8 FILLER_80_1042 ();
 sg13g2_decap_8 FILLER_80_1049 ();
 sg13g2_decap_4 FILLER_80_1056 ();
 sg13g2_fill_1 FILLER_80_1060 ();
 sg13g2_decap_8 FILLER_80_1066 ();
 sg13g2_decap_8 FILLER_80_1073 ();
 sg13g2_fill_2 FILLER_80_1080 ();
 sg13g2_decap_8 FILLER_80_1090 ();
 sg13g2_decap_8 FILLER_80_1104 ();
 sg13g2_decap_8 FILLER_80_1111 ();
 sg13g2_decap_8 FILLER_80_1118 ();
 sg13g2_decap_4 FILLER_80_1125 ();
 sg13g2_fill_2 FILLER_80_1129 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_4 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1265 ();
 sg13g2_decap_4 FILLER_80_1272 ();
 sg13g2_fill_2 FILLER_80_1279 ();
 sg13g2_fill_2 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1298 ();
 sg13g2_fill_1 FILLER_80_1305 ();
 sg13g2_decap_4 FILLER_80_1319 ();
 sg13g2_fill_2 FILLER_80_1323 ();
 sg13g2_fill_2 FILLER_80_1334 ();
 sg13g2_fill_1 FILLER_80_1336 ();
 sg13g2_fill_2 FILLER_80_1344 ();
 sg13g2_decap_8 FILLER_80_1362 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_decap_8 FILLER_80_1376 ();
 sg13g2_fill_2 FILLER_80_1383 ();
 sg13g2_fill_1 FILLER_80_1385 ();
 sg13g2_decap_8 FILLER_80_1392 ();
 sg13g2_decap_4 FILLER_80_1399 ();
 sg13g2_fill_1 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1408 ();
 sg13g2_decap_8 FILLER_80_1415 ();
 sg13g2_decap_4 FILLER_80_1430 ();
 sg13g2_fill_2 FILLER_80_1434 ();
 sg13g2_decap_8 FILLER_80_1463 ();
 sg13g2_decap_8 FILLER_80_1470 ();
 sg13g2_decap_8 FILLER_80_1477 ();
 sg13g2_decap_8 FILLER_80_1484 ();
 sg13g2_fill_2 FILLER_80_1491 ();
 sg13g2_decap_8 FILLER_80_1519 ();
 sg13g2_decap_8 FILLER_80_1526 ();
 sg13g2_fill_2 FILLER_80_1533 ();
 sg13g2_fill_1 FILLER_80_1535 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_4 FILLER_80_1564 ();
 sg13g2_fill_1 FILLER_80_1568 ();
 sg13g2_decap_8 FILLER_80_1608 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_fill_2 FILLER_80_1657 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_4 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_decap_8 FILLER_80_1701 ();
 sg13g2_decap_8 FILLER_80_1708 ();
 sg13g2_decap_8 FILLER_80_1715 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_fill_2 FILLER_80_1732 ();
 sg13g2_fill_1 FILLER_80_1734 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 sg13g2_decap_8 FILLER_81_0 ();
 sg13g2_decap_4 FILLER_81_7 ();
 sg13g2_decap_8 FILLER_81_36 ();
 sg13g2_decap_8 FILLER_81_43 ();
 sg13g2_decap_4 FILLER_81_50 ();
 sg13g2_fill_2 FILLER_81_54 ();
 sg13g2_fill_2 FILLER_81_68 ();
 sg13g2_decap_8 FILLER_81_74 ();
 sg13g2_fill_1 FILLER_81_81 ();
 sg13g2_decap_8 FILLER_81_91 ();
 sg13g2_decap_8 FILLER_81_98 ();
 sg13g2_decap_8 FILLER_81_105 ();
 sg13g2_decap_8 FILLER_81_112 ();
 sg13g2_decap_8 FILLER_81_119 ();
 sg13g2_decap_8 FILLER_81_126 ();
 sg13g2_decap_8 FILLER_81_133 ();
 sg13g2_decap_8 FILLER_81_140 ();
 sg13g2_decap_8 FILLER_81_147 ();
 sg13g2_decap_8 FILLER_81_154 ();
 sg13g2_decap_8 FILLER_81_161 ();
 sg13g2_decap_4 FILLER_81_168 ();
 sg13g2_fill_2 FILLER_81_172 ();
 sg13g2_decap_4 FILLER_81_178 ();
 sg13g2_fill_1 FILLER_81_182 ();
 sg13g2_decap_8 FILLER_81_196 ();
 sg13g2_decap_8 FILLER_81_203 ();
 sg13g2_decap_8 FILLER_81_210 ();
 sg13g2_decap_8 FILLER_81_217 ();
 sg13g2_fill_1 FILLER_81_224 ();
 sg13g2_fill_2 FILLER_81_233 ();
 sg13g2_decap_4 FILLER_81_240 ();
 sg13g2_fill_2 FILLER_81_244 ();
 sg13g2_decap_8 FILLER_81_251 ();
 sg13g2_decap_8 FILLER_81_258 ();
 sg13g2_decap_8 FILLER_81_265 ();
 sg13g2_decap_8 FILLER_81_272 ();
 sg13g2_decap_8 FILLER_81_279 ();
 sg13g2_decap_8 FILLER_81_286 ();
 sg13g2_decap_8 FILLER_81_293 ();
 sg13g2_decap_8 FILLER_81_300 ();
 sg13g2_decap_8 FILLER_81_307 ();
 sg13g2_decap_8 FILLER_81_314 ();
 sg13g2_decap_8 FILLER_81_321 ();
 sg13g2_decap_8 FILLER_81_328 ();
 sg13g2_decap_8 FILLER_81_335 ();
 sg13g2_fill_2 FILLER_81_342 ();
 sg13g2_fill_1 FILLER_81_344 ();
 sg13g2_decap_8 FILLER_81_353 ();
 sg13g2_decap_8 FILLER_81_368 ();
 sg13g2_decap_8 FILLER_81_381 ();
 sg13g2_decap_8 FILLER_81_388 ();
 sg13g2_decap_8 FILLER_81_395 ();
 sg13g2_decap_4 FILLER_81_402 ();
 sg13g2_fill_1 FILLER_81_406 ();
 sg13g2_decap_8 FILLER_81_413 ();
 sg13g2_fill_1 FILLER_81_420 ();
 sg13g2_decap_8 FILLER_81_424 ();
 sg13g2_decap_8 FILLER_81_431 ();
 sg13g2_decap_8 FILLER_81_438 ();
 sg13g2_decap_8 FILLER_81_445 ();
 sg13g2_decap_8 FILLER_81_452 ();
 sg13g2_decap_8 FILLER_81_459 ();
 sg13g2_decap_8 FILLER_81_466 ();
 sg13g2_decap_8 FILLER_81_473 ();
 sg13g2_decap_8 FILLER_81_480 ();
 sg13g2_decap_8 FILLER_81_487 ();
 sg13g2_decap_8 FILLER_81_494 ();
 sg13g2_decap_8 FILLER_81_501 ();
 sg13g2_decap_8 FILLER_81_508 ();
 sg13g2_decap_8 FILLER_81_515 ();
 sg13g2_fill_1 FILLER_81_522 ();
 sg13g2_decap_8 FILLER_81_531 ();
 sg13g2_decap_8 FILLER_81_538 ();
 sg13g2_decap_8 FILLER_81_545 ();
 sg13g2_decap_4 FILLER_81_552 ();
 sg13g2_fill_2 FILLER_81_556 ();
 sg13g2_decap_8 FILLER_81_580 ();
 sg13g2_decap_8 FILLER_81_587 ();
 sg13g2_decap_8 FILLER_81_594 ();
 sg13g2_decap_4 FILLER_81_601 ();
 sg13g2_fill_1 FILLER_81_605 ();
 sg13g2_fill_1 FILLER_81_611 ();
 sg13g2_decap_8 FILLER_81_620 ();
 sg13g2_decap_8 FILLER_81_627 ();
 sg13g2_decap_8 FILLER_81_634 ();
 sg13g2_decap_4 FILLER_81_641 ();
 sg13g2_fill_1 FILLER_81_645 ();
 sg13g2_fill_2 FILLER_81_688 ();
 sg13g2_decap_8 FILLER_81_702 ();
 sg13g2_decap_4 FILLER_81_709 ();
 sg13g2_fill_1 FILLER_81_713 ();
 sg13g2_decap_4 FILLER_81_719 ();
 sg13g2_decap_8 FILLER_81_731 ();
 sg13g2_decap_8 FILLER_81_738 ();
 sg13g2_decap_8 FILLER_81_745 ();
 sg13g2_decap_8 FILLER_81_752 ();
 sg13g2_decap_8 FILLER_81_759 ();
 sg13g2_decap_4 FILLER_81_766 ();
 sg13g2_fill_2 FILLER_81_770 ();
 sg13g2_decap_8 FILLER_81_776 ();
 sg13g2_decap_4 FILLER_81_783 ();
 sg13g2_decap_8 FILLER_81_792 ();
 sg13g2_decap_8 FILLER_81_799 ();
 sg13g2_decap_8 FILLER_81_844 ();
 sg13g2_decap_8 FILLER_81_851 ();
 sg13g2_decap_8 FILLER_81_858 ();
 sg13g2_decap_8 FILLER_81_865 ();
 sg13g2_fill_1 FILLER_81_872 ();
 sg13g2_decap_8 FILLER_81_877 ();
 sg13g2_decap_8 FILLER_81_884 ();
 sg13g2_decap_8 FILLER_81_891 ();
 sg13g2_decap_8 FILLER_81_898 ();
 sg13g2_decap_8 FILLER_81_905 ();
 sg13g2_decap_8 FILLER_81_912 ();
 sg13g2_decap_8 FILLER_81_919 ();
 sg13g2_decap_4 FILLER_81_926 ();
 sg13g2_fill_2 FILLER_81_930 ();
 sg13g2_decap_8 FILLER_81_936 ();
 sg13g2_decap_8 FILLER_81_943 ();
 sg13g2_decap_8 FILLER_81_950 ();
 sg13g2_decap_4 FILLER_81_957 ();
 sg13g2_fill_2 FILLER_81_961 ();
 sg13g2_decap_8 FILLER_81_981 ();
 sg13g2_decap_8 FILLER_81_988 ();
 sg13g2_decap_8 FILLER_81_995 ();
 sg13g2_fill_2 FILLER_81_1002 ();
 sg13g2_decap_8 FILLER_81_1017 ();
 sg13g2_decap_4 FILLER_81_1024 ();
 sg13g2_fill_2 FILLER_81_1028 ();
 sg13g2_decap_8 FILLER_81_1043 ();
 sg13g2_decap_4 FILLER_81_1050 ();
 sg13g2_fill_1 FILLER_81_1054 ();
 sg13g2_decap_8 FILLER_81_1106 ();
 sg13g2_decap_8 FILLER_81_1113 ();
 sg13g2_decap_8 FILLER_81_1120 ();
 sg13g2_fill_2 FILLER_81_1127 ();
 sg13g2_decap_8 FILLER_81_1137 ();
 sg13g2_decap_8 FILLER_81_1144 ();
 sg13g2_decap_8 FILLER_81_1151 ();
 sg13g2_decap_8 FILLER_81_1158 ();
 sg13g2_fill_2 FILLER_81_1165 ();
 sg13g2_fill_1 FILLER_81_1167 ();
 sg13g2_decap_8 FILLER_81_1194 ();
 sg13g2_decap_8 FILLER_81_1201 ();
 sg13g2_decap_8 FILLER_81_1208 ();
 sg13g2_fill_2 FILLER_81_1215 ();
 sg13g2_decap_4 FILLER_81_1225 ();
 sg13g2_decap_8 FILLER_81_1234 ();
 sg13g2_decap_8 FILLER_81_1241 ();
 sg13g2_decap_8 FILLER_81_1248 ();
 sg13g2_decap_8 FILLER_81_1255 ();
 sg13g2_decap_8 FILLER_81_1262 ();
 sg13g2_decap_8 FILLER_81_1269 ();
 sg13g2_decap_8 FILLER_81_1276 ();
 sg13g2_decap_8 FILLER_81_1283 ();
 sg13g2_decap_4 FILLER_81_1290 ();
 sg13g2_decap_8 FILLER_81_1310 ();
 sg13g2_decap_8 FILLER_81_1317 ();
 sg13g2_decap_8 FILLER_81_1324 ();
 sg13g2_decap_8 FILLER_81_1331 ();
 sg13g2_decap_4 FILLER_81_1338 ();
 sg13g2_fill_1 FILLER_81_1342 ();
 sg13g2_decap_8 FILLER_81_1353 ();
 sg13g2_decap_8 FILLER_81_1360 ();
 sg13g2_decap_8 FILLER_81_1367 ();
 sg13g2_decap_4 FILLER_81_1374 ();
 sg13g2_fill_2 FILLER_81_1378 ();
 sg13g2_decap_8 FILLER_81_1402 ();
 sg13g2_decap_8 FILLER_81_1409 ();
 sg13g2_decap_8 FILLER_81_1416 ();
 sg13g2_decap_8 FILLER_81_1423 ();
 sg13g2_fill_2 FILLER_81_1430 ();
 sg13g2_decap_8 FILLER_81_1473 ();
 sg13g2_decap_4 FILLER_81_1480 ();
 sg13g2_fill_2 FILLER_81_1503 ();
 sg13g2_fill_1 FILLER_81_1505 ();
 sg13g2_decap_8 FILLER_81_1519 ();
 sg13g2_decap_8 FILLER_81_1526 ();
 sg13g2_decap_8 FILLER_81_1533 ();
 sg13g2_decap_4 FILLER_81_1540 ();
 sg13g2_fill_2 FILLER_81_1544 ();
 sg13g2_decap_8 FILLER_81_1559 ();
 sg13g2_decap_8 FILLER_81_1566 ();
 sg13g2_decap_8 FILLER_81_1573 ();
 sg13g2_decap_8 FILLER_81_1584 ();
 sg13g2_decap_8 FILLER_81_1591 ();
 sg13g2_decap_8 FILLER_81_1598 ();
 sg13g2_decap_8 FILLER_81_1605 ();
 sg13g2_decap_8 FILLER_81_1612 ();
 sg13g2_decap_8 FILLER_81_1619 ();
 sg13g2_decap_8 FILLER_81_1626 ();
 sg13g2_decap_4 FILLER_81_1633 ();
 sg13g2_decap_8 FILLER_81_1647 ();
 sg13g2_decap_8 FILLER_81_1654 ();
 sg13g2_decap_8 FILLER_81_1661 ();
 sg13g2_decap_8 FILLER_81_1668 ();
 sg13g2_decap_8 FILLER_81_1675 ();
 sg13g2_fill_2 FILLER_81_1682 ();
 sg13g2_fill_1 FILLER_81_1684 ();
 sg13g2_decap_4 FILLER_81_1697 ();
 sg13g2_fill_1 FILLER_81_1701 ();
 sg13g2_decap_8 FILLER_81_1710 ();
 sg13g2_decap_4 FILLER_81_1717 ();
 sg13g2_fill_1 FILLER_81_1721 ();
 sg13g2_decap_8 FILLER_81_1732 ();
 sg13g2_decap_8 FILLER_81_1739 ();
 sg13g2_decap_8 FILLER_81_1750 ();
 sg13g2_decap_8 FILLER_81_1757 ();
 sg13g2_decap_4 FILLER_81_1764 ();
 sg13g2_decap_8 FILLER_82_0 ();
 sg13g2_decap_8 FILLER_82_7 ();
 sg13g2_decap_8 FILLER_82_14 ();
 sg13g2_fill_2 FILLER_82_21 ();
 sg13g2_decap_8 FILLER_82_26 ();
 sg13g2_decap_8 FILLER_82_33 ();
 sg13g2_decap_8 FILLER_82_40 ();
 sg13g2_decap_8 FILLER_82_47 ();
 sg13g2_decap_8 FILLER_82_54 ();
 sg13g2_decap_8 FILLER_82_61 ();
 sg13g2_decap_8 FILLER_82_68 ();
 sg13g2_fill_2 FILLER_82_75 ();
 sg13g2_decap_8 FILLER_82_86 ();
 sg13g2_decap_4 FILLER_82_93 ();
 sg13g2_fill_2 FILLER_82_97 ();
 sg13g2_decap_8 FILLER_82_113 ();
 sg13g2_decap_8 FILLER_82_120 ();
 sg13g2_decap_4 FILLER_82_127 ();
 sg13g2_fill_1 FILLER_82_131 ();
 sg13g2_decap_8 FILLER_82_153 ();
 sg13g2_decap_8 FILLER_82_160 ();
 sg13g2_decap_8 FILLER_82_167 ();
 sg13g2_decap_4 FILLER_82_174 ();
 sg13g2_decap_8 FILLER_82_186 ();
 sg13g2_decap_8 FILLER_82_193 ();
 sg13g2_decap_8 FILLER_82_200 ();
 sg13g2_decap_8 FILLER_82_207 ();
 sg13g2_decap_8 FILLER_82_214 ();
 sg13g2_fill_2 FILLER_82_221 ();
 sg13g2_fill_1 FILLER_82_223 ();
 sg13g2_decap_8 FILLER_82_232 ();
 sg13g2_decap_8 FILLER_82_239 ();
 sg13g2_decap_8 FILLER_82_246 ();
 sg13g2_decap_8 FILLER_82_253 ();
 sg13g2_decap_8 FILLER_82_260 ();
 sg13g2_decap_8 FILLER_82_267 ();
 sg13g2_decap_8 FILLER_82_274 ();
 sg13g2_decap_8 FILLER_82_281 ();
 sg13g2_decap_8 FILLER_82_288 ();
 sg13g2_fill_2 FILLER_82_295 ();
 sg13g2_fill_1 FILLER_82_297 ();
 sg13g2_decap_8 FILLER_82_303 ();
 sg13g2_fill_1 FILLER_82_310 ();
 sg13g2_decap_8 FILLER_82_315 ();
 sg13g2_decap_4 FILLER_82_322 ();
 sg13g2_decap_8 FILLER_82_336 ();
 sg13g2_fill_1 FILLER_82_343 ();
 sg13g2_fill_2 FILLER_82_364 ();
 sg13g2_decap_8 FILLER_82_370 ();
 sg13g2_decap_8 FILLER_82_377 ();
 sg13g2_decap_8 FILLER_82_384 ();
 sg13g2_fill_2 FILLER_82_391 ();
 sg13g2_fill_1 FILLER_82_393 ();
 sg13g2_fill_1 FILLER_82_398 ();
 sg13g2_decap_4 FILLER_82_412 ();
 sg13g2_fill_2 FILLER_82_416 ();
 sg13g2_decap_8 FILLER_82_423 ();
 sg13g2_decap_8 FILLER_82_430 ();
 sg13g2_decap_8 FILLER_82_437 ();
 sg13g2_decap_8 FILLER_82_444 ();
 sg13g2_decap_8 FILLER_82_451 ();
 sg13g2_decap_8 FILLER_82_458 ();
 sg13g2_decap_8 FILLER_82_465 ();
 sg13g2_fill_2 FILLER_82_472 ();
 sg13g2_fill_1 FILLER_82_474 ();
 sg13g2_decap_8 FILLER_82_491 ();
 sg13g2_decap_8 FILLER_82_498 ();
 sg13g2_decap_8 FILLER_82_505 ();
 sg13g2_decap_4 FILLER_82_512 ();
 sg13g2_fill_2 FILLER_82_516 ();
 sg13g2_decap_8 FILLER_82_538 ();
 sg13g2_decap_8 FILLER_82_545 ();
 sg13g2_decap_4 FILLER_82_552 ();
 sg13g2_fill_1 FILLER_82_556 ();
 sg13g2_decap_8 FILLER_82_570 ();
 sg13g2_decap_4 FILLER_82_577 ();
 sg13g2_decap_8 FILLER_82_593 ();
 sg13g2_fill_2 FILLER_82_600 ();
 sg13g2_fill_1 FILLER_82_615 ();
 sg13g2_decap_8 FILLER_82_624 ();
 sg13g2_decap_8 FILLER_82_631 ();
 sg13g2_decap_8 FILLER_82_638 ();
 sg13g2_decap_4 FILLER_82_645 ();
 sg13g2_fill_2 FILLER_82_649 ();
 sg13g2_fill_1 FILLER_82_665 ();
 sg13g2_fill_1 FILLER_82_670 ();
 sg13g2_decap_8 FILLER_82_693 ();
 sg13g2_fill_1 FILLER_82_700 ();
 sg13g2_decap_8 FILLER_82_740 ();
 sg13g2_decap_8 FILLER_82_747 ();
 sg13g2_decap_8 FILLER_82_754 ();
 sg13g2_decap_8 FILLER_82_761 ();
 sg13g2_fill_2 FILLER_82_768 ();
 sg13g2_decap_8 FILLER_82_788 ();
 sg13g2_decap_8 FILLER_82_795 ();
 sg13g2_fill_1 FILLER_82_802 ();
 sg13g2_decap_4 FILLER_82_815 ();
 sg13g2_fill_1 FILLER_82_819 ();
 sg13g2_fill_1 FILLER_82_824 ();
 sg13g2_fill_1 FILLER_82_851 ();
 sg13g2_decap_4 FILLER_82_861 ();
 sg13g2_fill_1 FILLER_82_865 ();
 sg13g2_decap_4 FILLER_82_891 ();
 sg13g2_fill_2 FILLER_82_895 ();
 sg13g2_decap_8 FILLER_82_910 ();
 sg13g2_decap_8 FILLER_82_917 ();
 sg13g2_decap_8 FILLER_82_924 ();
 sg13g2_decap_8 FILLER_82_931 ();
 sg13g2_fill_1 FILLER_82_938 ();
 sg13g2_decap_8 FILLER_82_964 ();
 sg13g2_decap_8 FILLER_82_971 ();
 sg13g2_decap_8 FILLER_82_978 ();
 sg13g2_decap_8 FILLER_82_985 ();
 sg13g2_decap_4 FILLER_82_992 ();
 sg13g2_fill_2 FILLER_82_1005 ();
 sg13g2_fill_1 FILLER_82_1007 ();
 sg13g2_decap_8 FILLER_82_1016 ();
 sg13g2_decap_8 FILLER_82_1023 ();
 sg13g2_decap_8 FILLER_82_1030 ();
 sg13g2_decap_8 FILLER_82_1037 ();
 sg13g2_decap_8 FILLER_82_1048 ();
 sg13g2_decap_8 FILLER_82_1055 ();
 sg13g2_fill_1 FILLER_82_1062 ();
 sg13g2_decap_8 FILLER_82_1071 ();
 sg13g2_decap_4 FILLER_82_1078 ();
 sg13g2_decap_4 FILLER_82_1091 ();
 sg13g2_decap_8 FILLER_82_1103 ();
 sg13g2_decap_4 FILLER_82_1110 ();
 sg13g2_decap_8 FILLER_82_1119 ();
 sg13g2_decap_4 FILLER_82_1126 ();
 sg13g2_decap_8 FILLER_82_1145 ();
 sg13g2_decap_4 FILLER_82_1152 ();
 sg13g2_fill_1 FILLER_82_1178 ();
 sg13g2_decap_8 FILLER_82_1183 ();
 sg13g2_decap_8 FILLER_82_1190 ();
 sg13g2_decap_8 FILLER_82_1197 ();
 sg13g2_decap_8 FILLER_82_1204 ();
 sg13g2_decap_8 FILLER_82_1211 ();
 sg13g2_decap_8 FILLER_82_1218 ();
 sg13g2_fill_1 FILLER_82_1225 ();
 sg13g2_fill_2 FILLER_82_1234 ();
 sg13g2_fill_1 FILLER_82_1236 ();
 sg13g2_fill_1 FILLER_82_1249 ();
 sg13g2_decap_4 FILLER_82_1260 ();
 sg13g2_decap_8 FILLER_82_1272 ();
 sg13g2_fill_2 FILLER_82_1279 ();
 sg13g2_decap_8 FILLER_82_1298 ();
 sg13g2_decap_8 FILLER_82_1305 ();
 sg13g2_decap_8 FILLER_82_1312 ();
 sg13g2_decap_8 FILLER_82_1319 ();
 sg13g2_decap_8 FILLER_82_1326 ();
 sg13g2_decap_8 FILLER_82_1333 ();
 sg13g2_decap_8 FILLER_82_1340 ();
 sg13g2_decap_8 FILLER_82_1347 ();
 sg13g2_decap_8 FILLER_82_1354 ();
 sg13g2_decap_8 FILLER_82_1361 ();
 sg13g2_decap_8 FILLER_82_1368 ();
 sg13g2_fill_1 FILLER_82_1375 ();
 sg13g2_decap_8 FILLER_82_1412 ();
 sg13g2_decap_8 FILLER_82_1419 ();
 sg13g2_decap_4 FILLER_82_1426 ();
 sg13g2_decap_8 FILLER_82_1440 ();
 sg13g2_decap_8 FILLER_82_1447 ();
 sg13g2_decap_8 FILLER_82_1454 ();
 sg13g2_fill_2 FILLER_82_1461 ();
 sg13g2_fill_1 FILLER_82_1463 ();
 sg13g2_fill_2 FILLER_82_1468 ();
 sg13g2_decap_8 FILLER_82_1475 ();
 sg13g2_decap_8 FILLER_82_1482 ();
 sg13g2_decap_4 FILLER_82_1489 ();
 sg13g2_fill_1 FILLER_82_1493 ();
 sg13g2_fill_1 FILLER_82_1511 ();
 sg13g2_decap_8 FILLER_82_1525 ();
 sg13g2_fill_1 FILLER_82_1532 ();
 sg13g2_decap_8 FILLER_82_1541 ();
 sg13g2_decap_8 FILLER_82_1548 ();
 sg13g2_decap_8 FILLER_82_1555 ();
 sg13g2_decap_8 FILLER_82_1562 ();
 sg13g2_decap_8 FILLER_82_1569 ();
 sg13g2_decap_8 FILLER_82_1576 ();
 sg13g2_decap_8 FILLER_82_1583 ();
 sg13g2_decap_8 FILLER_82_1590 ();
 sg13g2_decap_8 FILLER_82_1597 ();
 sg13g2_decap_4 FILLER_82_1604 ();
 sg13g2_fill_1 FILLER_82_1608 ();
 sg13g2_decap_8 FILLER_82_1622 ();
 sg13g2_fill_2 FILLER_82_1629 ();
 sg13g2_fill_1 FILLER_82_1631 ();
 sg13g2_decap_8 FILLER_82_1640 ();
 sg13g2_decap_8 FILLER_82_1647 ();
 sg13g2_decap_8 FILLER_82_1654 ();
 sg13g2_decap_8 FILLER_82_1661 ();
 sg13g2_decap_8 FILLER_82_1668 ();
 sg13g2_decap_8 FILLER_82_1675 ();
 sg13g2_decap_4 FILLER_82_1682 ();
 sg13g2_fill_2 FILLER_82_1686 ();
 sg13g2_fill_1 FILLER_82_1704 ();
 sg13g2_decap_8 FILLER_82_1731 ();
 sg13g2_decap_8 FILLER_82_1738 ();
 sg13g2_decap_8 FILLER_82_1745 ();
 sg13g2_decap_8 FILLER_82_1752 ();
 sg13g2_decap_8 FILLER_82_1759 ();
 sg13g2_fill_2 FILLER_82_1766 ();
 sg13g2_decap_8 FILLER_83_0 ();
 sg13g2_decap_8 FILLER_83_7 ();
 sg13g2_decap_8 FILLER_83_14 ();
 sg13g2_fill_2 FILLER_83_21 ();
 sg13g2_fill_1 FILLER_83_23 ();
 sg13g2_decap_8 FILLER_83_36 ();
 sg13g2_decap_8 FILLER_83_43 ();
 sg13g2_decap_4 FILLER_83_50 ();
 sg13g2_fill_2 FILLER_83_54 ();
 sg13g2_decap_8 FILLER_83_76 ();
 sg13g2_decap_8 FILLER_83_83 ();
 sg13g2_fill_2 FILLER_83_90 ();
 sg13g2_decap_8 FILLER_83_121 ();
 sg13g2_decap_8 FILLER_83_128 ();
 sg13g2_decap_8 FILLER_83_135 ();
 sg13g2_fill_1 FILLER_83_142 ();
 sg13g2_decap_8 FILLER_83_153 ();
 sg13g2_decap_8 FILLER_83_160 ();
 sg13g2_decap_8 FILLER_83_167 ();
 sg13g2_fill_2 FILLER_83_174 ();
 sg13g2_decap_8 FILLER_83_193 ();
 sg13g2_decap_8 FILLER_83_200 ();
 sg13g2_decap_4 FILLER_83_207 ();
 sg13g2_fill_2 FILLER_83_211 ();
 sg13g2_decap_4 FILLER_83_219 ();
 sg13g2_decap_8 FILLER_83_246 ();
 sg13g2_fill_1 FILLER_83_253 ();
 sg13g2_decap_8 FILLER_83_259 ();
 sg13g2_decap_8 FILLER_83_266 ();
 sg13g2_decap_4 FILLER_83_273 ();
 sg13g2_fill_2 FILLER_83_295 ();
 sg13g2_decap_8 FILLER_83_310 ();
 sg13g2_decap_8 FILLER_83_317 ();
 sg13g2_decap_8 FILLER_83_324 ();
 sg13g2_decap_8 FILLER_83_331 ();
 sg13g2_decap_8 FILLER_83_338 ();
 sg13g2_decap_8 FILLER_83_345 ();
 sg13g2_decap_8 FILLER_83_352 ();
 sg13g2_decap_8 FILLER_83_359 ();
 sg13g2_decap_8 FILLER_83_366 ();
 sg13g2_decap_8 FILLER_83_373 ();
 sg13g2_decap_8 FILLER_83_380 ();
 sg13g2_decap_8 FILLER_83_387 ();
 sg13g2_decap_4 FILLER_83_394 ();
 sg13g2_decap_8 FILLER_83_402 ();
 sg13g2_decap_8 FILLER_83_409 ();
 sg13g2_fill_2 FILLER_83_416 ();
 sg13g2_fill_1 FILLER_83_430 ();
 sg13g2_fill_2 FILLER_83_439 ();
 sg13g2_fill_2 FILLER_83_453 ();
 sg13g2_fill_1 FILLER_83_455 ();
 sg13g2_decap_8 FILLER_83_466 ();
 sg13g2_decap_4 FILLER_83_473 ();
 sg13g2_fill_2 FILLER_83_477 ();
 sg13g2_decap_8 FILLER_83_483 ();
 sg13g2_decap_8 FILLER_83_490 ();
 sg13g2_decap_8 FILLER_83_497 ();
 sg13g2_decap_8 FILLER_83_512 ();
 sg13g2_decap_4 FILLER_83_519 ();
 sg13g2_fill_2 FILLER_83_523 ();
 sg13g2_decap_8 FILLER_83_541 ();
 sg13g2_decap_8 FILLER_83_548 ();
 sg13g2_decap_8 FILLER_83_563 ();
 sg13g2_decap_8 FILLER_83_570 ();
 sg13g2_decap_8 FILLER_83_577 ();
 sg13g2_decap_8 FILLER_83_584 ();
 sg13g2_decap_8 FILLER_83_591 ();
 sg13g2_decap_8 FILLER_83_598 ();
 sg13g2_decap_8 FILLER_83_605 ();
 sg13g2_decap_4 FILLER_83_612 ();
 sg13g2_fill_1 FILLER_83_616 ();
 sg13g2_decap_8 FILLER_83_625 ();
 sg13g2_decap_8 FILLER_83_632 ();
 sg13g2_fill_2 FILLER_83_639 ();
 sg13g2_fill_1 FILLER_83_641 ();
 sg13g2_decap_8 FILLER_83_650 ();
 sg13g2_decap_8 FILLER_83_657 ();
 sg13g2_decap_8 FILLER_83_664 ();
 sg13g2_decap_8 FILLER_83_671 ();
 sg13g2_fill_2 FILLER_83_678 ();
 sg13g2_decap_8 FILLER_83_689 ();
 sg13g2_decap_8 FILLER_83_696 ();
 sg13g2_decap_8 FILLER_83_703 ();
 sg13g2_fill_2 FILLER_83_710 ();
 sg13g2_decap_8 FILLER_83_716 ();
 sg13g2_decap_4 FILLER_83_723 ();
 sg13g2_fill_2 FILLER_83_733 ();
 sg13g2_fill_1 FILLER_83_735 ();
 sg13g2_decap_8 FILLER_83_742 ();
 sg13g2_decap_8 FILLER_83_749 ();
 sg13g2_fill_2 FILLER_83_756 ();
 sg13g2_fill_1 FILLER_83_758 ();
 sg13g2_decap_8 FILLER_83_764 ();
 sg13g2_decap_8 FILLER_83_771 ();
 sg13g2_decap_8 FILLER_83_778 ();
 sg13g2_decap_8 FILLER_83_785 ();
 sg13g2_decap_8 FILLER_83_792 ();
 sg13g2_decap_8 FILLER_83_799 ();
 sg13g2_decap_8 FILLER_83_809 ();
 sg13g2_decap_8 FILLER_83_822 ();
 sg13g2_decap_8 FILLER_83_829 ();
 sg13g2_decap_8 FILLER_83_840 ();
 sg13g2_decap_8 FILLER_83_847 ();
 sg13g2_fill_2 FILLER_83_854 ();
 sg13g2_fill_1 FILLER_83_856 ();
 sg13g2_decap_8 FILLER_83_870 ();
 sg13g2_decap_8 FILLER_83_877 ();
 sg13g2_decap_8 FILLER_83_884 ();
 sg13g2_decap_8 FILLER_83_891 ();
 sg13g2_decap_8 FILLER_83_898 ();
 sg13g2_decap_8 FILLER_83_905 ();
 sg13g2_decap_8 FILLER_83_912 ();
 sg13g2_decap_8 FILLER_83_919 ();
 sg13g2_fill_2 FILLER_83_926 ();
 sg13g2_fill_1 FILLER_83_928 ();
 sg13g2_decap_8 FILLER_83_934 ();
 sg13g2_fill_2 FILLER_83_941 ();
 sg13g2_decap_8 FILLER_83_947 ();
 sg13g2_decap_8 FILLER_83_954 ();
 sg13g2_decap_8 FILLER_83_961 ();
 sg13g2_decap_8 FILLER_83_968 ();
 sg13g2_decap_8 FILLER_83_975 ();
 sg13g2_decap_8 FILLER_83_982 ();
 sg13g2_decap_4 FILLER_83_989 ();
 sg13g2_fill_2 FILLER_83_993 ();
 sg13g2_decap_4 FILLER_83_1021 ();
 sg13g2_fill_2 FILLER_83_1025 ();
 sg13g2_decap_8 FILLER_83_1043 ();
 sg13g2_decap_8 FILLER_83_1050 ();
 sg13g2_decap_8 FILLER_83_1057 ();
 sg13g2_decap_8 FILLER_83_1064 ();
 sg13g2_fill_2 FILLER_83_1071 ();
 sg13g2_decap_8 FILLER_83_1079 ();
 sg13g2_decap_8 FILLER_83_1086 ();
 sg13g2_decap_8 FILLER_83_1093 ();
 sg13g2_fill_2 FILLER_83_1100 ();
 sg13g2_decap_8 FILLER_83_1111 ();
 sg13g2_decap_8 FILLER_83_1118 ();
 sg13g2_decap_4 FILLER_83_1125 ();
 sg13g2_fill_2 FILLER_83_1129 ();
 sg13g2_decap_8 FILLER_83_1166 ();
 sg13g2_fill_2 FILLER_83_1173 ();
 sg13g2_fill_1 FILLER_83_1175 ();
 sg13g2_decap_8 FILLER_83_1179 ();
 sg13g2_decap_8 FILLER_83_1186 ();
 sg13g2_decap_8 FILLER_83_1193 ();
 sg13g2_fill_1 FILLER_83_1200 ();
 sg13g2_decap_8 FILLER_83_1206 ();
 sg13g2_decap_8 FILLER_83_1213 ();
 sg13g2_decap_8 FILLER_83_1220 ();
 sg13g2_fill_2 FILLER_83_1227 ();
 sg13g2_fill_1 FILLER_83_1229 ();
 sg13g2_fill_1 FILLER_83_1243 ();
 sg13g2_decap_8 FILLER_83_1250 ();
 sg13g2_decap_8 FILLER_83_1257 ();
 sg13g2_decap_8 FILLER_83_1264 ();
 sg13g2_fill_2 FILLER_83_1271 ();
 sg13g2_fill_1 FILLER_83_1273 ();
 sg13g2_decap_8 FILLER_83_1288 ();
 sg13g2_decap_8 FILLER_83_1295 ();
 sg13g2_decap_8 FILLER_83_1302 ();
 sg13g2_decap_8 FILLER_83_1309 ();
 sg13g2_decap_8 FILLER_83_1316 ();
 sg13g2_decap_8 FILLER_83_1323 ();
 sg13g2_fill_2 FILLER_83_1330 ();
 sg13g2_decap_8 FILLER_83_1348 ();
 sg13g2_decap_8 FILLER_83_1355 ();
 sg13g2_decap_8 FILLER_83_1362 ();
 sg13g2_decap_8 FILLER_83_1369 ();
 sg13g2_decap_8 FILLER_83_1376 ();
 sg13g2_fill_2 FILLER_83_1383 ();
 sg13g2_fill_1 FILLER_83_1385 ();
 sg13g2_fill_1 FILLER_83_1394 ();
 sg13g2_decap_8 FILLER_83_1405 ();
 sg13g2_decap_8 FILLER_83_1412 ();
 sg13g2_decap_8 FILLER_83_1419 ();
 sg13g2_decap_8 FILLER_83_1426 ();
 sg13g2_decap_8 FILLER_83_1433 ();
 sg13g2_decap_8 FILLER_83_1440 ();
 sg13g2_decap_8 FILLER_83_1447 ();
 sg13g2_decap_8 FILLER_83_1454 ();
 sg13g2_decap_4 FILLER_83_1461 ();
 sg13g2_fill_1 FILLER_83_1465 ();
 sg13g2_decap_8 FILLER_83_1492 ();
 sg13g2_decap_8 FILLER_83_1499 ();
 sg13g2_decap_8 FILLER_83_1506 ();
 sg13g2_decap_8 FILLER_83_1513 ();
 sg13g2_decap_8 FILLER_83_1520 ();
 sg13g2_decap_8 FILLER_83_1527 ();
 sg13g2_fill_2 FILLER_83_1534 ();
 sg13g2_decap_8 FILLER_83_1553 ();
 sg13g2_decap_8 FILLER_83_1560 ();
 sg13g2_decap_8 FILLER_83_1567 ();
 sg13g2_decap_8 FILLER_83_1574 ();
 sg13g2_decap_4 FILLER_83_1581 ();
 sg13g2_fill_2 FILLER_83_1585 ();
 sg13g2_decap_8 FILLER_83_1613 ();
 sg13g2_decap_8 FILLER_83_1620 ();
 sg13g2_decap_8 FILLER_83_1627 ();
 sg13g2_fill_2 FILLER_83_1644 ();
 sg13g2_decap_8 FILLER_83_1656 ();
 sg13g2_decap_8 FILLER_83_1663 ();
 sg13g2_decap_8 FILLER_83_1670 ();
 sg13g2_decap_8 FILLER_83_1677 ();
 sg13g2_decap_8 FILLER_83_1697 ();
 sg13g2_decap_8 FILLER_83_1704 ();
 sg13g2_decap_4 FILLER_83_1711 ();
 sg13g2_fill_1 FILLER_83_1715 ();
 sg13g2_decap_8 FILLER_83_1720 ();
 sg13g2_fill_2 FILLER_83_1727 ();
 sg13g2_fill_1 FILLER_83_1729 ();
 sg13g2_decap_8 FILLER_83_1743 ();
 sg13g2_decap_8 FILLER_83_1750 ();
 sg13g2_decap_8 FILLER_83_1757 ();
 sg13g2_decap_4 FILLER_83_1764 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_decap_8 FILLER_84_7 ();
 sg13g2_decap_8 FILLER_84_14 ();
 sg13g2_decap_4 FILLER_84_21 ();
 sg13g2_fill_1 FILLER_84_25 ();
 sg13g2_decap_8 FILLER_84_30 ();
 sg13g2_decap_4 FILLER_84_37 ();
 sg13g2_fill_2 FILLER_84_41 ();
 sg13g2_decap_8 FILLER_84_71 ();
 sg13g2_decap_8 FILLER_84_78 ();
 sg13g2_decap_8 FILLER_84_85 ();
 sg13g2_decap_8 FILLER_84_92 ();
 sg13g2_fill_2 FILLER_84_99 ();
 sg13g2_fill_2 FILLER_84_105 ();
 sg13g2_decap_8 FILLER_84_112 ();
 sg13g2_decap_8 FILLER_84_119 ();
 sg13g2_decap_8 FILLER_84_126 ();
 sg13g2_decap_4 FILLER_84_136 ();
 sg13g2_decap_8 FILLER_84_173 ();
 sg13g2_decap_8 FILLER_84_180 ();
 sg13g2_decap_8 FILLER_84_187 ();
 sg13g2_fill_2 FILLER_84_194 ();
 sg13g2_fill_1 FILLER_84_196 ();
 sg13g2_decap_8 FILLER_84_201 ();
 sg13g2_decap_8 FILLER_84_208 ();
 sg13g2_fill_1 FILLER_84_215 ();
 sg13g2_decap_8 FILLER_84_221 ();
 sg13g2_decap_8 FILLER_84_228 ();
 sg13g2_decap_8 FILLER_84_235 ();
 sg13g2_fill_1 FILLER_84_242 ();
 sg13g2_decap_8 FILLER_84_251 ();
 sg13g2_decap_8 FILLER_84_258 ();
 sg13g2_decap_8 FILLER_84_265 ();
 sg13g2_fill_2 FILLER_84_272 ();
 sg13g2_decap_8 FILLER_84_290 ();
 sg13g2_decap_8 FILLER_84_297 ();
 sg13g2_decap_8 FILLER_84_304 ();
 sg13g2_decap_8 FILLER_84_311 ();
 sg13g2_decap_8 FILLER_84_318 ();
 sg13g2_decap_8 FILLER_84_325 ();
 sg13g2_decap_4 FILLER_84_332 ();
 sg13g2_decap_4 FILLER_84_344 ();
 sg13g2_decap_4 FILLER_84_358 ();
 sg13g2_fill_1 FILLER_84_362 ();
 sg13g2_decap_8 FILLER_84_369 ();
 sg13g2_decap_8 FILLER_84_376 ();
 sg13g2_decap_8 FILLER_84_383 ();
 sg13g2_decap_8 FILLER_84_390 ();
 sg13g2_decap_8 FILLER_84_397 ();
 sg13g2_decap_8 FILLER_84_404 ();
 sg13g2_decap_8 FILLER_84_411 ();
 sg13g2_decap_4 FILLER_84_418 ();
 sg13g2_fill_2 FILLER_84_422 ();
 sg13g2_decap_8 FILLER_84_429 ();
 sg13g2_decap_8 FILLER_84_436 ();
 sg13g2_decap_4 FILLER_84_443 ();
 sg13g2_decap_4 FILLER_84_477 ();
 sg13g2_fill_2 FILLER_84_494 ();
 sg13g2_fill_1 FILLER_84_496 ();
 sg13g2_decap_8 FILLER_84_518 ();
 sg13g2_fill_2 FILLER_84_525 ();
 sg13g2_fill_1 FILLER_84_527 ();
 sg13g2_decap_8 FILLER_84_532 ();
 sg13g2_decap_8 FILLER_84_539 ();
 sg13g2_decap_8 FILLER_84_546 ();
 sg13g2_fill_2 FILLER_84_553 ();
 sg13g2_decap_8 FILLER_84_569 ();
 sg13g2_decap_4 FILLER_84_576 ();
 sg13g2_decap_8 FILLER_84_584 ();
 sg13g2_decap_8 FILLER_84_591 ();
 sg13g2_decap_8 FILLER_84_598 ();
 sg13g2_decap_8 FILLER_84_605 ();
 sg13g2_decap_4 FILLER_84_612 ();
 sg13g2_fill_2 FILLER_84_616 ();
 sg13g2_decap_8 FILLER_84_631 ();
 sg13g2_decap_8 FILLER_84_638 ();
 sg13g2_decap_8 FILLER_84_645 ();
 sg13g2_decap_8 FILLER_84_652 ();
 sg13g2_decap_8 FILLER_84_659 ();
 sg13g2_decap_8 FILLER_84_666 ();
 sg13g2_decap_8 FILLER_84_673 ();
 sg13g2_decap_8 FILLER_84_683 ();
 sg13g2_decap_8 FILLER_84_690 ();
 sg13g2_decap_8 FILLER_84_697 ();
 sg13g2_decap_8 FILLER_84_704 ();
 sg13g2_fill_2 FILLER_84_711 ();
 sg13g2_fill_1 FILLER_84_713 ();
 sg13g2_fill_2 FILLER_84_727 ();
 sg13g2_fill_1 FILLER_84_729 ();
 sg13g2_fill_2 FILLER_84_746 ();
 sg13g2_fill_1 FILLER_84_748 ();
 sg13g2_decap_8 FILLER_84_801 ();
 sg13g2_decap_8 FILLER_84_808 ();
 sg13g2_decap_8 FILLER_84_815 ();
 sg13g2_decap_8 FILLER_84_822 ();
 sg13g2_decap_8 FILLER_84_829 ();
 sg13g2_decap_8 FILLER_84_836 ();
 sg13g2_decap_8 FILLER_84_843 ();
 sg13g2_decap_8 FILLER_84_850 ();
 sg13g2_decap_8 FILLER_84_857 ();
 sg13g2_decap_8 FILLER_84_864 ();
 sg13g2_decap_8 FILLER_84_871 ();
 sg13g2_decap_8 FILLER_84_878 ();
 sg13g2_decap_8 FILLER_84_885 ();
 sg13g2_decap_8 FILLER_84_892 ();
 sg13g2_fill_1 FILLER_84_899 ();
 sg13g2_decap_8 FILLER_84_912 ();
 sg13g2_fill_1 FILLER_84_919 ();
 sg13g2_decap_4 FILLER_84_958 ();
 sg13g2_fill_1 FILLER_84_962 ();
 sg13g2_decap_8 FILLER_84_975 ();
 sg13g2_decap_8 FILLER_84_982 ();
 sg13g2_decap_4 FILLER_84_989 ();
 sg13g2_fill_1 FILLER_84_993 ();
 sg13g2_fill_2 FILLER_84_1003 ();
 sg13g2_decap_8 FILLER_84_1009 ();
 sg13g2_decap_8 FILLER_84_1016 ();
 sg13g2_fill_2 FILLER_84_1023 ();
 sg13g2_fill_2 FILLER_84_1038 ();
 sg13g2_fill_1 FILLER_84_1040 ();
 sg13g2_decap_8 FILLER_84_1049 ();
 sg13g2_decap_8 FILLER_84_1056 ();
 sg13g2_decap_8 FILLER_84_1063 ();
 sg13g2_decap_8 FILLER_84_1070 ();
 sg13g2_decap_8 FILLER_84_1077 ();
 sg13g2_decap_8 FILLER_84_1084 ();
 sg13g2_decap_8 FILLER_84_1091 ();
 sg13g2_fill_2 FILLER_84_1098 ();
 sg13g2_fill_1 FILLER_84_1100 ();
 sg13g2_decap_8 FILLER_84_1107 ();
 sg13g2_decap_8 FILLER_84_1114 ();
 sg13g2_decap_8 FILLER_84_1121 ();
 sg13g2_decap_8 FILLER_84_1128 ();
 sg13g2_decap_8 FILLER_84_1135 ();
 sg13g2_decap_8 FILLER_84_1142 ();
 sg13g2_fill_1 FILLER_84_1149 ();
 sg13g2_decap_8 FILLER_84_1154 ();
 sg13g2_decap_8 FILLER_84_1161 ();
 sg13g2_decap_4 FILLER_84_1168 ();
 sg13g2_fill_1 FILLER_84_1172 ();
 sg13g2_fill_1 FILLER_84_1186 ();
 sg13g2_fill_2 FILLER_84_1213 ();
 sg13g2_decap_8 FILLER_84_1228 ();
 sg13g2_decap_4 FILLER_84_1235 ();
 sg13g2_fill_1 FILLER_84_1239 ();
 sg13g2_decap_8 FILLER_84_1245 ();
 sg13g2_decap_8 FILLER_84_1252 ();
 sg13g2_decap_8 FILLER_84_1259 ();
 sg13g2_decap_8 FILLER_84_1266 ();
 sg13g2_decap_8 FILLER_84_1273 ();
 sg13g2_fill_1 FILLER_84_1280 ();
 sg13g2_decap_8 FILLER_84_1285 ();
 sg13g2_decap_8 FILLER_84_1292 ();
 sg13g2_decap_8 FILLER_84_1299 ();
 sg13g2_decap_8 FILLER_84_1306 ();
 sg13g2_decap_8 FILLER_84_1313 ();
 sg13g2_decap_8 FILLER_84_1320 ();
 sg13g2_decap_4 FILLER_84_1327 ();
 sg13g2_fill_1 FILLER_84_1331 ();
 sg13g2_decap_8 FILLER_84_1348 ();
 sg13g2_decap_8 FILLER_84_1368 ();
 sg13g2_decap_8 FILLER_84_1375 ();
 sg13g2_decap_8 FILLER_84_1382 ();
 sg13g2_decap_8 FILLER_84_1389 ();
 sg13g2_fill_2 FILLER_84_1396 ();
 sg13g2_fill_1 FILLER_84_1398 ();
 sg13g2_decap_8 FILLER_84_1409 ();
 sg13g2_decap_4 FILLER_84_1416 ();
 sg13g2_decap_8 FILLER_84_1424 ();
 sg13g2_decap_8 FILLER_84_1431 ();
 sg13g2_decap_8 FILLER_84_1438 ();
 sg13g2_decap_8 FILLER_84_1445 ();
 sg13g2_decap_8 FILLER_84_1460 ();
 sg13g2_decap_8 FILLER_84_1467 ();
 sg13g2_fill_2 FILLER_84_1474 ();
 sg13g2_fill_1 FILLER_84_1476 ();
 sg13g2_decap_8 FILLER_84_1481 ();
 sg13g2_decap_8 FILLER_84_1488 ();
 sg13g2_decap_8 FILLER_84_1495 ();
 sg13g2_decap_8 FILLER_84_1502 ();
 sg13g2_decap_8 FILLER_84_1509 ();
 sg13g2_decap_8 FILLER_84_1516 ();
 sg13g2_decap_8 FILLER_84_1523 ();
 sg13g2_decap_8 FILLER_84_1530 ();
 sg13g2_decap_8 FILLER_84_1537 ();
 sg13g2_fill_2 FILLER_84_1544 ();
 sg13g2_decap_8 FILLER_84_1564 ();
 sg13g2_fill_1 FILLER_84_1571 ();
 sg13g2_decap_8 FILLER_84_1575 ();
 sg13g2_decap_8 FILLER_84_1582 ();
 sg13g2_decap_8 FILLER_84_1589 ();
 sg13g2_fill_2 FILLER_84_1596 ();
 sg13g2_decap_8 FILLER_84_1602 ();
 sg13g2_decap_8 FILLER_84_1609 ();
 sg13g2_decap_8 FILLER_84_1616 ();
 sg13g2_decap_8 FILLER_84_1623 ();
 sg13g2_decap_8 FILLER_84_1630 ();
 sg13g2_decap_8 FILLER_84_1689 ();
 sg13g2_decap_8 FILLER_84_1696 ();
 sg13g2_decap_8 FILLER_84_1709 ();
 sg13g2_decap_8 FILLER_84_1716 ();
 sg13g2_decap_8 FILLER_84_1723 ();
 sg13g2_decap_8 FILLER_84_1730 ();
 sg13g2_decap_8 FILLER_84_1737 ();
 sg13g2_decap_8 FILLER_84_1744 ();
 sg13g2_decap_8 FILLER_84_1751 ();
 sg13g2_decap_8 FILLER_84_1758 ();
 sg13g2_fill_2 FILLER_84_1765 ();
 sg13g2_fill_1 FILLER_84_1767 ();
 sg13g2_decap_8 FILLER_85_0 ();
 sg13g2_decap_8 FILLER_85_7 ();
 sg13g2_fill_2 FILLER_85_14 ();
 sg13g2_decap_8 FILLER_85_33 ();
 sg13g2_decap_8 FILLER_85_40 ();
 sg13g2_decap_8 FILLER_85_47 ();
 sg13g2_decap_4 FILLER_85_54 ();
 sg13g2_fill_1 FILLER_85_58 ();
 sg13g2_decap_8 FILLER_85_63 ();
 sg13g2_decap_8 FILLER_85_70 ();
 sg13g2_decap_8 FILLER_85_77 ();
 sg13g2_decap_8 FILLER_85_84 ();
 sg13g2_decap_8 FILLER_85_91 ();
 sg13g2_decap_8 FILLER_85_98 ();
 sg13g2_fill_1 FILLER_85_105 ();
 sg13g2_decap_8 FILLER_85_126 ();
 sg13g2_decap_8 FILLER_85_133 ();
 sg13g2_decap_4 FILLER_85_140 ();
 sg13g2_fill_1 FILLER_85_144 ();
 sg13g2_fill_2 FILLER_85_151 ();
 sg13g2_decap_8 FILLER_85_162 ();
 sg13g2_decap_8 FILLER_85_169 ();
 sg13g2_decap_8 FILLER_85_176 ();
 sg13g2_decap_8 FILLER_85_183 ();
 sg13g2_decap_8 FILLER_85_190 ();
 sg13g2_decap_8 FILLER_85_197 ();
 sg13g2_decap_4 FILLER_85_204 ();
 sg13g2_fill_2 FILLER_85_208 ();
 sg13g2_fill_2 FILLER_85_223 ();
 sg13g2_fill_1 FILLER_85_225 ();
 sg13g2_decap_8 FILLER_85_231 ();
 sg13g2_decap_8 FILLER_85_238 ();
 sg13g2_decap_8 FILLER_85_245 ();
 sg13g2_decap_8 FILLER_85_252 ();
 sg13g2_decap_8 FILLER_85_259 ();
 sg13g2_decap_8 FILLER_85_266 ();
 sg13g2_decap_8 FILLER_85_273 ();
 sg13g2_decap_8 FILLER_85_280 ();
 sg13g2_decap_4 FILLER_85_287 ();
 sg13g2_fill_1 FILLER_85_291 ();
 sg13g2_decap_8 FILLER_85_296 ();
 sg13g2_fill_2 FILLER_85_303 ();
 sg13g2_fill_1 FILLER_85_305 ();
 sg13g2_decap_8 FILLER_85_314 ();
 sg13g2_decap_8 FILLER_85_321 ();
 sg13g2_decap_4 FILLER_85_328 ();
 sg13g2_fill_2 FILLER_85_332 ();
 sg13g2_decap_8 FILLER_85_347 ();
 sg13g2_fill_1 FILLER_85_362 ();
 sg13g2_decap_8 FILLER_85_374 ();
 sg13g2_decap_8 FILLER_85_381 ();
 sg13g2_decap_8 FILLER_85_388 ();
 sg13g2_decap_4 FILLER_85_395 ();
 sg13g2_fill_1 FILLER_85_399 ();
 sg13g2_decap_8 FILLER_85_404 ();
 sg13g2_decap_8 FILLER_85_411 ();
 sg13g2_decap_8 FILLER_85_418 ();
 sg13g2_decap_8 FILLER_85_425 ();
 sg13g2_decap_8 FILLER_85_432 ();
 sg13g2_decap_8 FILLER_85_439 ();
 sg13g2_decap_4 FILLER_85_446 ();
 sg13g2_fill_2 FILLER_85_450 ();
 sg13g2_fill_1 FILLER_85_457 ();
 sg13g2_decap_8 FILLER_85_468 ();
 sg13g2_decap_8 FILLER_85_475 ();
 sg13g2_decap_8 FILLER_85_482 ();
 sg13g2_decap_8 FILLER_85_489 ();
 sg13g2_fill_2 FILLER_85_496 ();
 sg13g2_decap_8 FILLER_85_511 ();
 sg13g2_decap_8 FILLER_85_518 ();
 sg13g2_decap_8 FILLER_85_525 ();
 sg13g2_decap_8 FILLER_85_532 ();
 sg13g2_decap_8 FILLER_85_539 ();
 sg13g2_decap_8 FILLER_85_546 ();
 sg13g2_decap_8 FILLER_85_553 ();
 sg13g2_decap_4 FILLER_85_560 ();
 sg13g2_decap_8 FILLER_85_572 ();
 sg13g2_decap_8 FILLER_85_579 ();
 sg13g2_decap_8 FILLER_85_586 ();
 sg13g2_decap_8 FILLER_85_614 ();
 sg13g2_decap_8 FILLER_85_621 ();
 sg13g2_decap_8 FILLER_85_628 ();
 sg13g2_decap_8 FILLER_85_635 ();
 sg13g2_decap_8 FILLER_85_642 ();
 sg13g2_decap_4 FILLER_85_649 ();
 sg13g2_fill_2 FILLER_85_679 ();
 sg13g2_decap_8 FILLER_85_694 ();
 sg13g2_decap_8 FILLER_85_701 ();
 sg13g2_decap_8 FILLER_85_708 ();
 sg13g2_decap_8 FILLER_85_715 ();
 sg13g2_decap_8 FILLER_85_722 ();
 sg13g2_decap_8 FILLER_85_729 ();
 sg13g2_decap_8 FILLER_85_742 ();
 sg13g2_decap_4 FILLER_85_749 ();
 sg13g2_fill_2 FILLER_85_753 ();
 sg13g2_fill_1 FILLER_85_761 ();
 sg13g2_decap_4 FILLER_85_766 ();
 sg13g2_fill_2 FILLER_85_770 ();
 sg13g2_decap_8 FILLER_85_777 ();
 sg13g2_fill_2 FILLER_85_784 ();
 sg13g2_decap_8 FILLER_85_790 ();
 sg13g2_decap_8 FILLER_85_797 ();
 sg13g2_decap_8 FILLER_85_804 ();
 sg13g2_decap_4 FILLER_85_811 ();
 sg13g2_fill_2 FILLER_85_815 ();
 sg13g2_decap_8 FILLER_85_827 ();
 sg13g2_decap_8 FILLER_85_834 ();
 sg13g2_decap_8 FILLER_85_841 ();
 sg13g2_decap_8 FILLER_85_848 ();
 sg13g2_decap_8 FILLER_85_855 ();
 sg13g2_fill_1 FILLER_85_862 ();
 sg13g2_decap_4 FILLER_85_868 ();
 sg13g2_fill_1 FILLER_85_872 ();
 sg13g2_decap_8 FILLER_85_884 ();
 sg13g2_fill_1 FILLER_85_891 ();
 sg13g2_decap_8 FILLER_85_918 ();
 sg13g2_decap_4 FILLER_85_925 ();
 sg13g2_fill_1 FILLER_85_929 ();
 sg13g2_decap_8 FILLER_85_935 ();
 sg13g2_decap_8 FILLER_85_942 ();
 sg13g2_decap_8 FILLER_85_949 ();
 sg13g2_fill_1 FILLER_85_956 ();
 sg13g2_decap_8 FILLER_85_965 ();
 sg13g2_decap_8 FILLER_85_972 ();
 sg13g2_decap_8 FILLER_85_979 ();
 sg13g2_decap_8 FILLER_85_986 ();
 sg13g2_decap_8 FILLER_85_993 ();
 sg13g2_decap_8 FILLER_85_1000 ();
 sg13g2_decap_8 FILLER_85_1007 ();
 sg13g2_decap_8 FILLER_85_1014 ();
 sg13g2_fill_1 FILLER_85_1021 ();
 sg13g2_decap_8 FILLER_85_1030 ();
 sg13g2_decap_8 FILLER_85_1037 ();
 sg13g2_decap_8 FILLER_85_1044 ();
 sg13g2_fill_1 FILLER_85_1056 ();
 sg13g2_decap_8 FILLER_85_1061 ();
 sg13g2_decap_8 FILLER_85_1068 ();
 sg13g2_decap_8 FILLER_85_1075 ();
 sg13g2_decap_8 FILLER_85_1082 ();
 sg13g2_decap_8 FILLER_85_1089 ();
 sg13g2_decap_8 FILLER_85_1096 ();
 sg13g2_decap_8 FILLER_85_1103 ();
 sg13g2_decap_8 FILLER_85_1110 ();
 sg13g2_fill_1 FILLER_85_1121 ();
 sg13g2_decap_8 FILLER_85_1132 ();
 sg13g2_decap_8 FILLER_85_1139 ();
 sg13g2_decap_8 FILLER_85_1146 ();
 sg13g2_decap_8 FILLER_85_1153 ();
 sg13g2_decap_8 FILLER_85_1160 ();
 sg13g2_decap_8 FILLER_85_1167 ();
 sg13g2_fill_2 FILLER_85_1174 ();
 sg13g2_decap_8 FILLER_85_1182 ();
 sg13g2_decap_8 FILLER_85_1189 ();
 sg13g2_fill_2 FILLER_85_1196 ();
 sg13g2_decap_8 FILLER_85_1205 ();
 sg13g2_fill_2 FILLER_85_1212 ();
 sg13g2_decap_8 FILLER_85_1223 ();
 sg13g2_decap_8 FILLER_85_1230 ();
 sg13g2_decap_8 FILLER_85_1237 ();
 sg13g2_decap_8 FILLER_85_1244 ();
 sg13g2_decap_4 FILLER_85_1251 ();
 sg13g2_fill_1 FILLER_85_1255 ();
 sg13g2_decap_8 FILLER_85_1265 ();
 sg13g2_decap_4 FILLER_85_1272 ();
 sg13g2_fill_2 FILLER_85_1281 ();
 sg13g2_decap_8 FILLER_85_1291 ();
 sg13g2_decap_8 FILLER_85_1298 ();
 sg13g2_decap_8 FILLER_85_1305 ();
 sg13g2_decap_8 FILLER_85_1312 ();
 sg13g2_fill_2 FILLER_85_1319 ();
 sg13g2_decap_8 FILLER_85_1325 ();
 sg13g2_fill_1 FILLER_85_1332 ();
 sg13g2_decap_8 FILLER_85_1340 ();
 sg13g2_decap_8 FILLER_85_1347 ();
 sg13g2_decap_8 FILLER_85_1354 ();
 sg13g2_decap_8 FILLER_85_1361 ();
 sg13g2_decap_8 FILLER_85_1368 ();
 sg13g2_decap_4 FILLER_85_1375 ();
 sg13g2_fill_1 FILLER_85_1379 ();
 sg13g2_decap_4 FILLER_85_1386 ();
 sg13g2_fill_2 FILLER_85_1390 ();
 sg13g2_fill_2 FILLER_85_1397 ();
 sg13g2_decap_8 FILLER_85_1408 ();
 sg13g2_fill_2 FILLER_85_1415 ();
 sg13g2_decap_8 FILLER_85_1435 ();
 sg13g2_decap_8 FILLER_85_1442 ();
 sg13g2_decap_8 FILLER_85_1449 ();
 sg13g2_decap_8 FILLER_85_1456 ();
 sg13g2_decap_8 FILLER_85_1463 ();
 sg13g2_decap_8 FILLER_85_1470 ();
 sg13g2_fill_2 FILLER_85_1477 ();
 sg13g2_fill_1 FILLER_85_1479 ();
 sg13g2_decap_8 FILLER_85_1493 ();
 sg13g2_decap_8 FILLER_85_1500 ();
 sg13g2_decap_8 FILLER_85_1507 ();
 sg13g2_decap_8 FILLER_85_1514 ();
 sg13g2_decap_8 FILLER_85_1521 ();
 sg13g2_decap_8 FILLER_85_1528 ();
 sg13g2_decap_8 FILLER_85_1535 ();
 sg13g2_decap_8 FILLER_85_1542 ();
 sg13g2_fill_1 FILLER_85_1549 ();
 sg13g2_decap_8 FILLER_85_1554 ();
 sg13g2_decap_8 FILLER_85_1561 ();
 sg13g2_fill_1 FILLER_85_1568 ();
 sg13g2_fill_1 FILLER_85_1580 ();
 sg13g2_decap_8 FILLER_85_1588 ();
 sg13g2_decap_8 FILLER_85_1595 ();
 sg13g2_decap_8 FILLER_85_1602 ();
 sg13g2_decap_8 FILLER_85_1609 ();
 sg13g2_decap_8 FILLER_85_1616 ();
 sg13g2_decap_8 FILLER_85_1623 ();
 sg13g2_decap_8 FILLER_85_1630 ();
 sg13g2_decap_8 FILLER_85_1637 ();
 sg13g2_decap_4 FILLER_85_1644 ();
 sg13g2_fill_1 FILLER_85_1648 ();
 sg13g2_decap_8 FILLER_85_1658 ();
 sg13g2_decap_4 FILLER_85_1665 ();
 sg13g2_fill_2 FILLER_85_1669 ();
 sg13g2_decap_8 FILLER_85_1675 ();
 sg13g2_decap_8 FILLER_85_1682 ();
 sg13g2_decap_8 FILLER_85_1689 ();
 sg13g2_decap_8 FILLER_85_1696 ();
 sg13g2_decap_8 FILLER_85_1709 ();
 sg13g2_decap_8 FILLER_85_1716 ();
 sg13g2_decap_8 FILLER_85_1723 ();
 sg13g2_decap_8 FILLER_85_1730 ();
 sg13g2_decap_4 FILLER_85_1737 ();
 sg13g2_fill_2 FILLER_85_1766 ();
 sg13g2_decap_8 FILLER_86_0 ();
 sg13g2_decap_8 FILLER_86_7 ();
 sg13g2_decap_8 FILLER_86_14 ();
 sg13g2_decap_8 FILLER_86_21 ();
 sg13g2_fill_2 FILLER_86_28 ();
 sg13g2_decap_8 FILLER_86_38 ();
 sg13g2_decap_8 FILLER_86_45 ();
 sg13g2_decap_8 FILLER_86_52 ();
 sg13g2_decap_8 FILLER_86_59 ();
 sg13g2_decap_4 FILLER_86_66 ();
 sg13g2_fill_1 FILLER_86_70 ();
 sg13g2_fill_1 FILLER_86_79 ();
 sg13g2_decap_8 FILLER_86_85 ();
 sg13g2_decap_8 FILLER_86_92 ();
 sg13g2_decap_8 FILLER_86_99 ();
 sg13g2_decap_8 FILLER_86_106 ();
 sg13g2_decap_8 FILLER_86_113 ();
 sg13g2_fill_2 FILLER_86_120 ();
 sg13g2_fill_1 FILLER_86_122 ();
 sg13g2_decap_8 FILLER_86_133 ();
 sg13g2_decap_8 FILLER_86_140 ();
 sg13g2_decap_4 FILLER_86_147 ();
 sg13g2_fill_2 FILLER_86_151 ();
 sg13g2_decap_8 FILLER_86_165 ();
 sg13g2_decap_8 FILLER_86_172 ();
 sg13g2_decap_8 FILLER_86_179 ();
 sg13g2_decap_8 FILLER_86_186 ();
 sg13g2_decap_8 FILLER_86_193 ();
 sg13g2_decap_8 FILLER_86_200 ();
 sg13g2_decap_8 FILLER_86_207 ();
 sg13g2_decap_8 FILLER_86_214 ();
 sg13g2_decap_8 FILLER_86_229 ();
 sg13g2_decap_8 FILLER_86_236 ();
 sg13g2_decap_8 FILLER_86_243 ();
 sg13g2_decap_8 FILLER_86_250 ();
 sg13g2_decap_8 FILLER_86_257 ();
 sg13g2_decap_8 FILLER_86_264 ();
 sg13g2_fill_2 FILLER_86_271 ();
 sg13g2_decap_4 FILLER_86_277 ();
 sg13g2_fill_1 FILLER_86_281 ();
 sg13g2_decap_8 FILLER_86_290 ();
 sg13g2_decap_8 FILLER_86_297 ();
 sg13g2_decap_8 FILLER_86_304 ();
 sg13g2_decap_8 FILLER_86_311 ();
 sg13g2_decap_4 FILLER_86_318 ();
 sg13g2_fill_2 FILLER_86_322 ();
 sg13g2_decap_8 FILLER_86_328 ();
 sg13g2_decap_8 FILLER_86_335 ();
 sg13g2_fill_2 FILLER_86_342 ();
 sg13g2_decap_8 FILLER_86_382 ();
 sg13g2_decap_4 FILLER_86_389 ();
 sg13g2_fill_1 FILLER_86_407 ();
 sg13g2_decap_8 FILLER_86_420 ();
 sg13g2_decap_8 FILLER_86_427 ();
 sg13g2_decap_8 FILLER_86_434 ();
 sg13g2_decap_8 FILLER_86_441 ();
 sg13g2_decap_8 FILLER_86_448 ();
 sg13g2_decap_8 FILLER_86_455 ();
 sg13g2_decap_8 FILLER_86_462 ();
 sg13g2_decap_8 FILLER_86_469 ();
 sg13g2_decap_8 FILLER_86_476 ();
 sg13g2_decap_8 FILLER_86_483 ();
 sg13g2_decap_8 FILLER_86_490 ();
 sg13g2_decap_4 FILLER_86_505 ();
 sg13g2_fill_1 FILLER_86_509 ();
 sg13g2_fill_2 FILLER_86_518 ();
 sg13g2_fill_1 FILLER_86_520 ();
 sg13g2_decap_8 FILLER_86_529 ();
 sg13g2_decap_8 FILLER_86_536 ();
 sg13g2_decap_8 FILLER_86_543 ();
 sg13g2_decap_8 FILLER_86_550 ();
 sg13g2_decap_8 FILLER_86_557 ();
 sg13g2_decap_8 FILLER_86_564 ();
 sg13g2_decap_8 FILLER_86_571 ();
 sg13g2_decap_8 FILLER_86_578 ();
 sg13g2_decap_8 FILLER_86_585 ();
 sg13g2_fill_1 FILLER_86_592 ();
 sg13g2_fill_1 FILLER_86_601 ();
 sg13g2_decap_8 FILLER_86_610 ();
 sg13g2_fill_1 FILLER_86_617 ();
 sg13g2_decap_8 FILLER_86_622 ();
 sg13g2_decap_8 FILLER_86_629 ();
 sg13g2_decap_8 FILLER_86_636 ();
 sg13g2_decap_8 FILLER_86_643 ();
 sg13g2_decap_8 FILLER_86_671 ();
 sg13g2_fill_2 FILLER_86_678 ();
 sg13g2_fill_1 FILLER_86_694 ();
 sg13g2_decap_8 FILLER_86_699 ();
 sg13g2_fill_2 FILLER_86_706 ();
 sg13g2_fill_1 FILLER_86_708 ();
 sg13g2_fill_1 FILLER_86_713 ();
 sg13g2_decap_8 FILLER_86_722 ();
 sg13g2_decap_8 FILLER_86_729 ();
 sg13g2_decap_8 FILLER_86_736 ();
 sg13g2_decap_8 FILLER_86_743 ();
 sg13g2_decap_4 FILLER_86_750 ();
 sg13g2_fill_1 FILLER_86_754 ();
 sg13g2_decap_8 FILLER_86_761 ();
 sg13g2_decap_8 FILLER_86_768 ();
 sg13g2_decap_8 FILLER_86_775 ();
 sg13g2_decap_8 FILLER_86_782 ();
 sg13g2_decap_8 FILLER_86_789 ();
 sg13g2_decap_8 FILLER_86_796 ();
 sg13g2_decap_8 FILLER_86_803 ();
 sg13g2_decap_4 FILLER_86_823 ();
 sg13g2_decap_8 FILLER_86_840 ();
 sg13g2_fill_2 FILLER_86_847 ();
 sg13g2_fill_1 FILLER_86_849 ();
 sg13g2_fill_2 FILLER_86_863 ();
 sg13g2_decap_8 FILLER_86_888 ();
 sg13g2_decap_8 FILLER_86_895 ();
 sg13g2_fill_1 FILLER_86_902 ();
 sg13g2_decap_8 FILLER_86_920 ();
 sg13g2_decap_8 FILLER_86_927 ();
 sg13g2_decap_8 FILLER_86_947 ();
 sg13g2_decap_8 FILLER_86_954 ();
 sg13g2_fill_1 FILLER_86_961 ();
 sg13g2_decap_8 FILLER_86_972 ();
 sg13g2_decap_8 FILLER_86_979 ();
 sg13g2_decap_8 FILLER_86_986 ();
 sg13g2_decap_8 FILLER_86_993 ();
 sg13g2_decap_8 FILLER_86_1000 ();
 sg13g2_decap_8 FILLER_86_1007 ();
 sg13g2_decap_8 FILLER_86_1014 ();
 sg13g2_fill_2 FILLER_86_1021 ();
 sg13g2_decap_8 FILLER_86_1027 ();
 sg13g2_decap_8 FILLER_86_1034 ();
 sg13g2_fill_2 FILLER_86_1041 ();
 sg13g2_fill_1 FILLER_86_1043 ();
 sg13g2_decap_4 FILLER_86_1052 ();
 sg13g2_decap_4 FILLER_86_1082 ();
 sg13g2_fill_2 FILLER_86_1086 ();
 sg13g2_decap_4 FILLER_86_1101 ();
 sg13g2_fill_2 FILLER_86_1105 ();
 sg13g2_decap_8 FILLER_86_1146 ();
 sg13g2_decap_8 FILLER_86_1153 ();
 sg13g2_decap_8 FILLER_86_1160 ();
 sg13g2_decap_8 FILLER_86_1167 ();
 sg13g2_fill_2 FILLER_86_1174 ();
 sg13g2_decap_8 FILLER_86_1184 ();
 sg13g2_decap_8 FILLER_86_1191 ();
 sg13g2_decap_8 FILLER_86_1198 ();
 sg13g2_decap_4 FILLER_86_1205 ();
 sg13g2_fill_1 FILLER_86_1209 ();
 sg13g2_decap_8 FILLER_86_1218 ();
 sg13g2_decap_8 FILLER_86_1225 ();
 sg13g2_decap_8 FILLER_86_1232 ();
 sg13g2_decap_8 FILLER_86_1239 ();
 sg13g2_decap_8 FILLER_86_1246 ();
 sg13g2_fill_2 FILLER_86_1253 ();
 sg13g2_fill_1 FILLER_86_1255 ();
 sg13g2_fill_1 FILLER_86_1261 ();
 sg13g2_decap_8 FILLER_86_1291 ();
 sg13g2_decap_8 FILLER_86_1298 ();
 sg13g2_decap_8 FILLER_86_1305 ();
 sg13g2_fill_2 FILLER_86_1312 ();
 sg13g2_decap_8 FILLER_86_1326 ();
 sg13g2_decap_8 FILLER_86_1333 ();
 sg13g2_decap_8 FILLER_86_1340 ();
 sg13g2_decap_8 FILLER_86_1347 ();
 sg13g2_decap_8 FILLER_86_1354 ();
 sg13g2_decap_4 FILLER_86_1361 ();
 sg13g2_decap_8 FILLER_86_1391 ();
 sg13g2_decap_4 FILLER_86_1398 ();
 sg13g2_fill_1 FILLER_86_1402 ();
 sg13g2_decap_8 FILLER_86_1411 ();
 sg13g2_fill_1 FILLER_86_1418 ();
 sg13g2_decap_8 FILLER_86_1445 ();
 sg13g2_decap_8 FILLER_86_1452 ();
 sg13g2_decap_8 FILLER_86_1459 ();
 sg13g2_decap_4 FILLER_86_1466 ();
 sg13g2_fill_2 FILLER_86_1470 ();
 sg13g2_fill_2 FILLER_86_1497 ();
 sg13g2_fill_1 FILLER_86_1513 ();
 sg13g2_decap_8 FILLER_86_1518 ();
 sg13g2_fill_2 FILLER_86_1525 ();
 sg13g2_fill_1 FILLER_86_1527 ();
 sg13g2_fill_2 FILLER_86_1536 ();
 sg13g2_fill_2 FILLER_86_1543 ();
 sg13g2_decap_8 FILLER_86_1552 ();
 sg13g2_decap_8 FILLER_86_1559 ();
 sg13g2_fill_2 FILLER_86_1566 ();
 sg13g2_decap_8 FILLER_86_1594 ();
 sg13g2_decap_4 FILLER_86_1601 ();
 sg13g2_fill_2 FILLER_86_1605 ();
 sg13g2_decap_8 FILLER_86_1610 ();
 sg13g2_decap_8 FILLER_86_1617 ();
 sg13g2_fill_1 FILLER_86_1624 ();
 sg13g2_fill_1 FILLER_86_1629 ();
 sg13g2_decap_8 FILLER_86_1655 ();
 sg13g2_decap_8 FILLER_86_1662 ();
 sg13g2_decap_8 FILLER_86_1669 ();
 sg13g2_decap_8 FILLER_86_1676 ();
 sg13g2_decap_8 FILLER_86_1683 ();
 sg13g2_decap_8 FILLER_86_1690 ();
 sg13g2_decap_8 FILLER_86_1719 ();
 sg13g2_decap_8 FILLER_86_1752 ();
 sg13g2_decap_8 FILLER_86_1759 ();
 sg13g2_fill_2 FILLER_86_1766 ();
 sg13g2_decap_8 FILLER_87_0 ();
 sg13g2_decap_8 FILLER_87_7 ();
 sg13g2_decap_4 FILLER_87_14 ();
 sg13g2_decap_8 FILLER_87_26 ();
 sg13g2_fill_2 FILLER_87_33 ();
 sg13g2_fill_1 FILLER_87_35 ();
 sg13g2_decap_8 FILLER_87_46 ();
 sg13g2_decap_8 FILLER_87_53 ();
 sg13g2_decap_4 FILLER_87_60 ();
 sg13g2_fill_1 FILLER_87_64 ();
 sg13g2_fill_2 FILLER_87_79 ();
 sg13g2_decap_4 FILLER_87_86 ();
 sg13g2_fill_1 FILLER_87_90 ();
 sg13g2_decap_8 FILLER_87_99 ();
 sg13g2_decap_8 FILLER_87_106 ();
 sg13g2_decap_8 FILLER_87_113 ();
 sg13g2_decap_8 FILLER_87_120 ();
 sg13g2_decap_8 FILLER_87_127 ();
 sg13g2_decap_8 FILLER_87_134 ();
 sg13g2_decap_8 FILLER_87_141 ();
 sg13g2_fill_2 FILLER_87_148 ();
 sg13g2_decap_8 FILLER_87_158 ();
 sg13g2_decap_8 FILLER_87_173 ();
 sg13g2_decap_8 FILLER_87_180 ();
 sg13g2_decap_8 FILLER_87_187 ();
 sg13g2_decap_8 FILLER_87_194 ();
 sg13g2_fill_2 FILLER_87_201 ();
 sg13g2_decap_8 FILLER_87_211 ();
 sg13g2_decap_4 FILLER_87_218 ();
 sg13g2_decap_8 FILLER_87_226 ();
 sg13g2_fill_2 FILLER_87_233 ();
 sg13g2_fill_1 FILLER_87_235 ();
 sg13g2_decap_8 FILLER_87_244 ();
 sg13g2_decap_8 FILLER_87_251 ();
 sg13g2_decap_8 FILLER_87_258 ();
 sg13g2_fill_1 FILLER_87_265 ();
 sg13g2_fill_1 FILLER_87_279 ();
 sg13g2_decap_8 FILLER_87_288 ();
 sg13g2_decap_8 FILLER_87_304 ();
 sg13g2_decap_8 FILLER_87_323 ();
 sg13g2_decap_8 FILLER_87_330 ();
 sg13g2_decap_8 FILLER_87_337 ();
 sg13g2_decap_8 FILLER_87_344 ();
 sg13g2_fill_2 FILLER_87_351 ();
 sg13g2_fill_1 FILLER_87_353 ();
 sg13g2_fill_1 FILLER_87_362 ();
 sg13g2_fill_1 FILLER_87_366 ();
 sg13g2_decap_8 FILLER_87_378 ();
 sg13g2_decap_4 FILLER_87_385 ();
 sg13g2_fill_2 FILLER_87_389 ();
 sg13g2_decap_8 FILLER_87_403 ();
 sg13g2_decap_8 FILLER_87_425 ();
 sg13g2_decap_8 FILLER_87_432 ();
 sg13g2_fill_2 FILLER_87_439 ();
 sg13g2_fill_1 FILLER_87_441 ();
 sg13g2_fill_2 FILLER_87_449 ();
 sg13g2_decap_8 FILLER_87_455 ();
 sg13g2_decap_8 FILLER_87_462 ();
 sg13g2_decap_8 FILLER_87_469 ();
 sg13g2_decap_8 FILLER_87_476 ();
 sg13g2_decap_8 FILLER_87_483 ();
 sg13g2_decap_8 FILLER_87_490 ();
 sg13g2_decap_8 FILLER_87_497 ();
 sg13g2_decap_8 FILLER_87_504 ();
 sg13g2_decap_8 FILLER_87_511 ();
 sg13g2_fill_2 FILLER_87_518 ();
 sg13g2_fill_1 FILLER_87_520 ();
 sg13g2_decap_8 FILLER_87_526 ();
 sg13g2_decap_4 FILLER_87_533 ();
 sg13g2_fill_1 FILLER_87_537 ();
 sg13g2_decap_8 FILLER_87_554 ();
 sg13g2_decap_8 FILLER_87_561 ();
 sg13g2_decap_8 FILLER_87_568 ();
 sg13g2_decap_8 FILLER_87_575 ();
 sg13g2_decap_8 FILLER_87_582 ();
 sg13g2_decap_8 FILLER_87_589 ();
 sg13g2_decap_8 FILLER_87_596 ();
 sg13g2_decap_8 FILLER_87_603 ();
 sg13g2_decap_8 FILLER_87_628 ();
 sg13g2_fill_2 FILLER_87_635 ();
 sg13g2_decap_4 FILLER_87_650 ();
 sg13g2_decap_8 FILLER_87_666 ();
 sg13g2_decap_8 FILLER_87_673 ();
 sg13g2_decap_4 FILLER_87_680 ();
 sg13g2_fill_2 FILLER_87_710 ();
 sg13g2_fill_1 FILLER_87_712 ();
 sg13g2_decap_4 FILLER_87_726 ();
 sg13g2_fill_2 FILLER_87_730 ();
 sg13g2_decap_8 FILLER_87_737 ();
 sg13g2_decap_4 FILLER_87_744 ();
 sg13g2_fill_1 FILLER_87_748 ();
 sg13g2_decap_8 FILLER_87_769 ();
 sg13g2_decap_8 FILLER_87_776 ();
 sg13g2_decap_4 FILLER_87_783 ();
 sg13g2_fill_1 FILLER_87_787 ();
 sg13g2_decap_8 FILLER_87_801 ();
 sg13g2_fill_2 FILLER_87_808 ();
 sg13g2_fill_1 FILLER_87_810 ();
 sg13g2_decap_8 FILLER_87_829 ();
 sg13g2_decap_8 FILLER_87_836 ();
 sg13g2_fill_1 FILLER_87_843 ();
 sg13g2_decap_8 FILLER_87_852 ();
 sg13g2_decap_8 FILLER_87_859 ();
 sg13g2_decap_8 FILLER_87_866 ();
 sg13g2_decap_8 FILLER_87_884 ();
 sg13g2_decap_8 FILLER_87_891 ();
 sg13g2_decap_4 FILLER_87_898 ();
 sg13g2_fill_1 FILLER_87_902 ();
 sg13g2_decap_8 FILLER_87_912 ();
 sg13g2_decap_8 FILLER_87_919 ();
 sg13g2_decap_8 FILLER_87_926 ();
 sg13g2_decap_8 FILLER_87_933 ();
 sg13g2_decap_8 FILLER_87_940 ();
 sg13g2_decap_8 FILLER_87_947 ();
 sg13g2_decap_8 FILLER_87_954 ();
 sg13g2_decap_8 FILLER_87_1013 ();
 sg13g2_decap_8 FILLER_87_1020 ();
 sg13g2_decap_8 FILLER_87_1027 ();
 sg13g2_decap_8 FILLER_87_1034 ();
 sg13g2_decap_4 FILLER_87_1041 ();
 sg13g2_fill_1 FILLER_87_1045 ();
 sg13g2_decap_8 FILLER_87_1055 ();
 sg13g2_decap_4 FILLER_87_1062 ();
 sg13g2_decap_8 FILLER_87_1070 ();
 sg13g2_decap_8 FILLER_87_1077 ();
 sg13g2_fill_1 FILLER_87_1084 ();
 sg13g2_decap_8 FILLER_87_1098 ();
 sg13g2_decap_8 FILLER_87_1105 ();
 sg13g2_fill_2 FILLER_87_1112 ();
 sg13g2_fill_1 FILLER_87_1114 ();
 sg13g2_decap_4 FILLER_87_1124 ();
 sg13g2_fill_2 FILLER_87_1128 ();
 sg13g2_decap_8 FILLER_87_1139 ();
 sg13g2_decap_8 FILLER_87_1146 ();
 sg13g2_decap_4 FILLER_87_1153 ();
 sg13g2_fill_1 FILLER_87_1157 ();
 sg13g2_decap_4 FILLER_87_1171 ();
 sg13g2_fill_1 FILLER_87_1175 ();
 sg13g2_decap_8 FILLER_87_1184 ();
 sg13g2_fill_2 FILLER_87_1191 ();
 sg13g2_fill_2 FILLER_87_1198 ();
 sg13g2_decap_4 FILLER_87_1203 ();
 sg13g2_fill_1 FILLER_87_1207 ();
 sg13g2_fill_2 FILLER_87_1216 ();
 sg13g2_fill_1 FILLER_87_1218 ();
 sg13g2_decap_8 FILLER_87_1227 ();
 sg13g2_decap_8 FILLER_87_1234 ();
 sg13g2_decap_8 FILLER_87_1241 ();
 sg13g2_decap_8 FILLER_87_1248 ();
 sg13g2_fill_2 FILLER_87_1259 ();
 sg13g2_fill_1 FILLER_87_1261 ();
 sg13g2_decap_8 FILLER_87_1286 ();
 sg13g2_decap_8 FILLER_87_1293 ();
 sg13g2_decap_4 FILLER_87_1300 ();
 sg13g2_fill_1 FILLER_87_1304 ();
 sg13g2_decap_8 FILLER_87_1336 ();
 sg13g2_decap_8 FILLER_87_1343 ();
 sg13g2_fill_1 FILLER_87_1350 ();
 sg13g2_decap_4 FILLER_87_1356 ();
 sg13g2_fill_2 FILLER_87_1360 ();
 sg13g2_decap_4 FILLER_87_1371 ();
 sg13g2_decap_8 FILLER_87_1388 ();
 sg13g2_decap_8 FILLER_87_1395 ();
 sg13g2_decap_8 FILLER_87_1402 ();
 sg13g2_decap_8 FILLER_87_1409 ();
 sg13g2_decap_8 FILLER_87_1416 ();
 sg13g2_decap_8 FILLER_87_1423 ();
 sg13g2_decap_8 FILLER_87_1430 ();
 sg13g2_decap_8 FILLER_87_1437 ();
 sg13g2_decap_8 FILLER_87_1444 ();
 sg13g2_decap_8 FILLER_87_1451 ();
 sg13g2_decap_8 FILLER_87_1458 ();
 sg13g2_decap_8 FILLER_87_1465 ();
 sg13g2_decap_8 FILLER_87_1472 ();
 sg13g2_decap_8 FILLER_87_1479 ();
 sg13g2_fill_2 FILLER_87_1486 ();
 sg13g2_fill_2 FILLER_87_1514 ();
 sg13g2_fill_1 FILLER_87_1516 ();
 sg13g2_fill_1 FILLER_87_1587 ();
 sg13g2_fill_2 FILLER_87_1612 ();
 sg13g2_decap_8 FILLER_87_1649 ();
 sg13g2_decap_8 FILLER_87_1656 ();
 sg13g2_decap_8 FILLER_87_1663 ();
 sg13g2_decap_8 FILLER_87_1670 ();
 sg13g2_fill_2 FILLER_87_1709 ();
 sg13g2_fill_1 FILLER_87_1748 ();
 sg13g2_decap_8 FILLER_87_1758 ();
 sg13g2_fill_2 FILLER_87_1765 ();
 sg13g2_fill_1 FILLER_87_1767 ();
 sg13g2_decap_8 FILLER_88_0 ();
 sg13g2_decap_8 FILLER_88_7 ();
 sg13g2_decap_8 FILLER_88_14 ();
 sg13g2_fill_1 FILLER_88_21 ();
 sg13g2_fill_2 FILLER_88_27 ();
 sg13g2_fill_1 FILLER_88_34 ();
 sg13g2_decap_8 FILLER_88_38 ();
 sg13g2_decap_8 FILLER_88_45 ();
 sg13g2_decap_8 FILLER_88_52 ();
 sg13g2_decap_8 FILLER_88_59 ();
 sg13g2_decap_4 FILLER_88_66 ();
 sg13g2_fill_2 FILLER_88_70 ();
 sg13g2_decap_8 FILLER_88_77 ();
 sg13g2_decap_8 FILLER_88_84 ();
 sg13g2_decap_8 FILLER_88_91 ();
 sg13g2_decap_8 FILLER_88_98 ();
 sg13g2_decap_8 FILLER_88_105 ();
 sg13g2_decap_8 FILLER_88_112 ();
 sg13g2_decap_8 FILLER_88_119 ();
 sg13g2_decap_8 FILLER_88_126 ();
 sg13g2_decap_8 FILLER_88_133 ();
 sg13g2_decap_8 FILLER_88_140 ();
 sg13g2_decap_4 FILLER_88_147 ();
 sg13g2_fill_1 FILLER_88_151 ();
 sg13g2_decap_8 FILLER_88_164 ();
 sg13g2_fill_2 FILLER_88_181 ();
 sg13g2_decap_8 FILLER_88_191 ();
 sg13g2_fill_2 FILLER_88_198 ();
 sg13g2_fill_1 FILLER_88_200 ();
 sg13g2_fill_1 FILLER_88_214 ();
 sg13g2_fill_1 FILLER_88_228 ();
 sg13g2_decap_8 FILLER_88_235 ();
 sg13g2_decap_8 FILLER_88_242 ();
 sg13g2_decap_8 FILLER_88_249 ();
 sg13g2_fill_1 FILLER_88_256 ();
 sg13g2_fill_1 FILLER_88_283 ();
 sg13g2_decap_8 FILLER_88_298 ();
 sg13g2_decap_8 FILLER_88_305 ();
 sg13g2_decap_8 FILLER_88_312 ();
 sg13g2_decap_8 FILLER_88_319 ();
 sg13g2_decap_8 FILLER_88_326 ();
 sg13g2_fill_1 FILLER_88_333 ();
 sg13g2_decap_8 FILLER_88_338 ();
 sg13g2_decap_8 FILLER_88_345 ();
 sg13g2_decap_8 FILLER_88_352 ();
 sg13g2_decap_4 FILLER_88_359 ();
 sg13g2_decap_8 FILLER_88_375 ();
 sg13g2_decap_8 FILLER_88_382 ();
 sg13g2_decap_8 FILLER_88_389 ();
 sg13g2_decap_4 FILLER_88_396 ();
 sg13g2_fill_1 FILLER_88_400 ();
 sg13g2_fill_1 FILLER_88_421 ();
 sg13g2_fill_1 FILLER_88_439 ();
 sg13g2_decap_8 FILLER_88_461 ();
 sg13g2_decap_8 FILLER_88_468 ();
 sg13g2_decap_8 FILLER_88_475 ();
 sg13g2_decap_8 FILLER_88_482 ();
 sg13g2_decap_4 FILLER_88_489 ();
 sg13g2_fill_2 FILLER_88_493 ();
 sg13g2_decap_4 FILLER_88_505 ();
 sg13g2_fill_2 FILLER_88_515 ();
 sg13g2_fill_1 FILLER_88_517 ();
 sg13g2_decap_8 FILLER_88_531 ();
 sg13g2_decap_8 FILLER_88_538 ();
 sg13g2_decap_8 FILLER_88_545 ();
 sg13g2_decap_8 FILLER_88_552 ();
 sg13g2_decap_8 FILLER_88_559 ();
 sg13g2_decap_8 FILLER_88_566 ();
 sg13g2_decap_8 FILLER_88_573 ();
 sg13g2_decap_8 FILLER_88_580 ();
 sg13g2_decap_4 FILLER_88_587 ();
 sg13g2_decap_8 FILLER_88_595 ();
 sg13g2_decap_8 FILLER_88_602 ();
 sg13g2_decap_8 FILLER_88_609 ();
 sg13g2_decap_8 FILLER_88_616 ();
 sg13g2_decap_8 FILLER_88_623 ();
 sg13g2_decap_8 FILLER_88_630 ();
 sg13g2_decap_8 FILLER_88_637 ();
 sg13g2_decap_8 FILLER_88_644 ();
 sg13g2_fill_1 FILLER_88_651 ();
 sg13g2_decap_8 FILLER_88_665 ();
 sg13g2_decap_4 FILLER_88_672 ();
 sg13g2_fill_2 FILLER_88_676 ();
 sg13g2_decap_8 FILLER_88_688 ();
 sg13g2_decap_8 FILLER_88_695 ();
 sg13g2_decap_8 FILLER_88_702 ();
 sg13g2_decap_8 FILLER_88_709 ();
 sg13g2_decap_8 FILLER_88_716 ();
 sg13g2_decap_4 FILLER_88_723 ();
 sg13g2_fill_2 FILLER_88_727 ();
 sg13g2_decap_8 FILLER_88_770 ();
 sg13g2_decap_4 FILLER_88_777 ();
 sg13g2_fill_2 FILLER_88_781 ();
 sg13g2_decap_8 FILLER_88_796 ();
 sg13g2_decap_8 FILLER_88_803 ();
 sg13g2_decap_8 FILLER_88_810 ();
 sg13g2_decap_8 FILLER_88_817 ();
 sg13g2_decap_8 FILLER_88_824 ();
 sg13g2_decap_8 FILLER_88_831 ();
 sg13g2_decap_8 FILLER_88_838 ();
 sg13g2_decap_8 FILLER_88_845 ();
 sg13g2_decap_8 FILLER_88_852 ();
 sg13g2_decap_8 FILLER_88_859 ();
 sg13g2_decap_8 FILLER_88_866 ();
 sg13g2_decap_8 FILLER_88_873 ();
 sg13g2_decap_8 FILLER_88_880 ();
 sg13g2_decap_8 FILLER_88_887 ();
 sg13g2_fill_2 FILLER_88_894 ();
 sg13g2_fill_1 FILLER_88_896 ();
 sg13g2_decap_8 FILLER_88_913 ();
 sg13g2_decap_8 FILLER_88_920 ();
 sg13g2_decap_8 FILLER_88_927 ();
 sg13g2_decap_8 FILLER_88_934 ();
 sg13g2_decap_8 FILLER_88_941 ();
 sg13g2_decap_8 FILLER_88_948 ();
 sg13g2_decap_8 FILLER_88_955 ();
 sg13g2_decap_8 FILLER_88_962 ();
 sg13g2_decap_8 FILLER_88_969 ();
 sg13g2_decap_8 FILLER_88_976 ();
 sg13g2_fill_2 FILLER_88_983 ();
 sg13g2_decap_8 FILLER_88_989 ();
 sg13g2_decap_8 FILLER_88_996 ();
 sg13g2_decap_8 FILLER_88_1003 ();
 sg13g2_decap_8 FILLER_88_1010 ();
 sg13g2_fill_2 FILLER_88_1017 ();
 sg13g2_fill_1 FILLER_88_1019 ();
 sg13g2_decap_8 FILLER_88_1033 ();
 sg13g2_decap_8 FILLER_88_1040 ();
 sg13g2_fill_2 FILLER_88_1047 ();
 sg13g2_fill_1 FILLER_88_1065 ();
 sg13g2_decap_8 FILLER_88_1074 ();
 sg13g2_decap_8 FILLER_88_1081 ();
 sg13g2_decap_8 FILLER_88_1088 ();
 sg13g2_decap_8 FILLER_88_1095 ();
 sg13g2_decap_8 FILLER_88_1102 ();
 sg13g2_decap_8 FILLER_88_1109 ();
 sg13g2_fill_1 FILLER_88_1116 ();
 sg13g2_decap_8 FILLER_88_1125 ();
 sg13g2_fill_2 FILLER_88_1132 ();
 sg13g2_fill_1 FILLER_88_1134 ();
 sg13g2_decap_4 FILLER_88_1143 ();
 sg13g2_decap_4 FILLER_88_1151 ();
 sg13g2_fill_2 FILLER_88_1155 ();
 sg13g2_decap_8 FILLER_88_1183 ();
 sg13g2_decap_8 FILLER_88_1190 ();
 sg13g2_fill_1 FILLER_88_1197 ();
 sg13g2_fill_2 FILLER_88_1233 ();
 sg13g2_fill_1 FILLER_88_1235 ();
 sg13g2_decap_8 FILLER_88_1265 ();
 sg13g2_decap_8 FILLER_88_1272 ();
 sg13g2_decap_8 FILLER_88_1279 ();
 sg13g2_decap_8 FILLER_88_1286 ();
 sg13g2_decap_8 FILLER_88_1293 ();
 sg13g2_decap_8 FILLER_88_1300 ();
 sg13g2_fill_1 FILLER_88_1307 ();
 sg13g2_fill_2 FILLER_88_1325 ();
 sg13g2_fill_1 FILLER_88_1327 ();
 sg13g2_decap_8 FILLER_88_1337 ();
 sg13g2_decap_8 FILLER_88_1344 ();
 sg13g2_decap_8 FILLER_88_1351 ();
 sg13g2_decap_8 FILLER_88_1358 ();
 sg13g2_decap_4 FILLER_88_1365 ();
 sg13g2_fill_2 FILLER_88_1369 ();
 sg13g2_decap_8 FILLER_88_1375 ();
 sg13g2_decap_8 FILLER_88_1382 ();
 sg13g2_decap_8 FILLER_88_1389 ();
 sg13g2_decap_8 FILLER_88_1396 ();
 sg13g2_decap_8 FILLER_88_1403 ();
 sg13g2_decap_4 FILLER_88_1410 ();
 sg13g2_fill_2 FILLER_88_1414 ();
 sg13g2_decap_8 FILLER_88_1429 ();
 sg13g2_decap_4 FILLER_88_1462 ();
 sg13g2_fill_1 FILLER_88_1466 ();
 sg13g2_decap_8 FILLER_88_1471 ();
 sg13g2_decap_8 FILLER_88_1483 ();
 sg13g2_decap_4 FILLER_88_1490 ();
 sg13g2_fill_1 FILLER_88_1494 ();
 sg13g2_decap_8 FILLER_88_1517 ();
 sg13g2_decap_8 FILLER_88_1524 ();
 sg13g2_decap_8 FILLER_88_1531 ();
 sg13g2_decap_8 FILLER_88_1538 ();
 sg13g2_decap_8 FILLER_88_1548 ();
 sg13g2_decap_8 FILLER_88_1555 ();
 sg13g2_decap_8 FILLER_88_1567 ();
 sg13g2_fill_2 FILLER_88_1582 ();
 sg13g2_fill_1 FILLER_88_1587 ();
 sg13g2_decap_8 FILLER_88_1594 ();
 sg13g2_decap_4 FILLER_88_1601 ();
 sg13g2_fill_2 FILLER_88_1605 ();
 sg13g2_decap_8 FILLER_88_1610 ();
 sg13g2_fill_2 FILLER_88_1617 ();
 sg13g2_decap_8 FILLER_88_1631 ();
 sg13g2_decap_8 FILLER_88_1638 ();
 sg13g2_decap_8 FILLER_88_1645 ();
 sg13g2_decap_8 FILLER_88_1652 ();
 sg13g2_decap_8 FILLER_88_1659 ();
 sg13g2_fill_2 FILLER_88_1666 ();
 sg13g2_fill_1 FILLER_88_1668 ();
 sg13g2_decap_8 FILLER_88_1685 ();
 sg13g2_decap_8 FILLER_88_1724 ();
 sg13g2_decap_8 FILLER_88_1731 ();
 sg13g2_decap_8 FILLER_88_1738 ();
 sg13g2_decap_8 FILLER_88_1745 ();
 sg13g2_decap_8 FILLER_88_1752 ();
 sg13g2_decap_8 FILLER_88_1759 ();
 sg13g2_fill_2 FILLER_88_1766 ();
 sg13g2_decap_8 FILLER_89_0 ();
 sg13g2_decap_8 FILLER_89_7 ();
 sg13g2_fill_2 FILLER_89_14 ();
 sg13g2_decap_8 FILLER_89_33 ();
 sg13g2_decap_8 FILLER_89_40 ();
 sg13g2_decap_8 FILLER_89_47 ();
 sg13g2_decap_8 FILLER_89_58 ();
 sg13g2_decap_8 FILLER_89_65 ();
 sg13g2_decap_8 FILLER_89_72 ();
 sg13g2_decap_8 FILLER_89_79 ();
 sg13g2_decap_4 FILLER_89_86 ();
 sg13g2_decap_8 FILLER_89_102 ();
 sg13g2_decap_8 FILLER_89_109 ();
 sg13g2_decap_8 FILLER_89_116 ();
 sg13g2_decap_8 FILLER_89_123 ();
 sg13g2_decap_8 FILLER_89_130 ();
 sg13g2_decap_8 FILLER_89_137 ();
 sg13g2_decap_8 FILLER_89_144 ();
 sg13g2_fill_1 FILLER_89_151 ();
 sg13g2_decap_8 FILLER_89_157 ();
 sg13g2_fill_1 FILLER_89_164 ();
 sg13g2_decap_4 FILLER_89_173 ();
 sg13g2_fill_1 FILLER_89_177 ();
 sg13g2_decap_4 FILLER_89_193 ();
 sg13g2_fill_2 FILLER_89_197 ();
 sg13g2_fill_1 FILLER_89_209 ();
 sg13g2_decap_4 FILLER_89_217 ();
 sg13g2_decap_8 FILLER_89_242 ();
 sg13g2_decap_8 FILLER_89_249 ();
 sg13g2_decap_8 FILLER_89_256 ();
 sg13g2_decap_4 FILLER_89_263 ();
 sg13g2_decap_8 FILLER_89_304 ();
 sg13g2_decap_8 FILLER_89_311 ();
 sg13g2_decap_8 FILLER_89_318 ();
 sg13g2_decap_4 FILLER_89_325 ();
 sg13g2_fill_1 FILLER_89_329 ();
 sg13g2_decap_8 FILLER_89_346 ();
 sg13g2_decap_8 FILLER_89_353 ();
 sg13g2_decap_8 FILLER_89_360 ();
 sg13g2_decap_8 FILLER_89_367 ();
 sg13g2_decap_8 FILLER_89_374 ();
 sg13g2_decap_8 FILLER_89_381 ();
 sg13g2_decap_4 FILLER_89_388 ();
 sg13g2_fill_2 FILLER_89_392 ();
 sg13g2_fill_1 FILLER_89_402 ();
 sg13g2_fill_2 FILLER_89_414 ();
 sg13g2_decap_8 FILLER_89_424 ();
 sg13g2_decap_8 FILLER_89_431 ();
 sg13g2_decap_4 FILLER_89_438 ();
 sg13g2_fill_2 FILLER_89_442 ();
 sg13g2_decap_8 FILLER_89_449 ();
 sg13g2_decap_8 FILLER_89_465 ();
 sg13g2_decap_8 FILLER_89_472 ();
 sg13g2_decap_8 FILLER_89_479 ();
 sg13g2_fill_2 FILLER_89_486 ();
 sg13g2_fill_1 FILLER_89_502 ();
 sg13g2_decap_8 FILLER_89_534 ();
 sg13g2_decap_8 FILLER_89_541 ();
 sg13g2_decap_8 FILLER_89_548 ();
 sg13g2_decap_8 FILLER_89_555 ();
 sg13g2_decap_8 FILLER_89_562 ();
 sg13g2_decap_8 FILLER_89_569 ();
 sg13g2_fill_2 FILLER_89_576 ();
 sg13g2_fill_1 FILLER_89_578 ();
 sg13g2_decap_8 FILLER_89_603 ();
 sg13g2_fill_2 FILLER_89_610 ();
 sg13g2_fill_1 FILLER_89_612 ();
 sg13g2_decap_8 FILLER_89_626 ();
 sg13g2_decap_8 FILLER_89_633 ();
 sg13g2_decap_8 FILLER_89_640 ();
 sg13g2_decap_8 FILLER_89_647 ();
 sg13g2_decap_8 FILLER_89_654 ();
 sg13g2_decap_8 FILLER_89_661 ();
 sg13g2_decap_8 FILLER_89_668 ();
 sg13g2_decap_8 FILLER_89_675 ();
 sg13g2_decap_8 FILLER_89_682 ();
 sg13g2_decap_8 FILLER_89_689 ();
 sg13g2_decap_8 FILLER_89_696 ();
 sg13g2_decap_8 FILLER_89_703 ();
 sg13g2_decap_8 FILLER_89_710 ();
 sg13g2_decap_8 FILLER_89_717 ();
 sg13g2_fill_1 FILLER_89_724 ();
 sg13g2_fill_2 FILLER_89_735 ();
 sg13g2_fill_1 FILLER_89_737 ();
 sg13g2_fill_2 FILLER_89_768 ();
 sg13g2_fill_1 FILLER_89_770 ();
 sg13g2_decap_8 FILLER_89_797 ();
 sg13g2_decap_8 FILLER_89_804 ();
 sg13g2_decap_8 FILLER_89_811 ();
 sg13g2_decap_8 FILLER_89_818 ();
 sg13g2_decap_8 FILLER_89_851 ();
 sg13g2_decap_8 FILLER_89_858 ();
 sg13g2_fill_2 FILLER_89_865 ();
 sg13g2_decap_8 FILLER_89_880 ();
 sg13g2_decap_8 FILLER_89_887 ();
 sg13g2_fill_1 FILLER_89_894 ();
 sg13g2_decap_8 FILLER_89_919 ();
 sg13g2_decap_8 FILLER_89_926 ();
 sg13g2_decap_8 FILLER_89_933 ();
 sg13g2_decap_8 FILLER_89_940 ();
 sg13g2_decap_8 FILLER_89_947 ();
 sg13g2_decap_8 FILLER_89_954 ();
 sg13g2_decap_8 FILLER_89_961 ();
 sg13g2_decap_8 FILLER_89_968 ();
 sg13g2_decap_8 FILLER_89_975 ();
 sg13g2_decap_8 FILLER_89_982 ();
 sg13g2_decap_8 FILLER_89_989 ();
 sg13g2_decap_8 FILLER_89_996 ();
 sg13g2_decap_8 FILLER_89_1003 ();
 sg13g2_fill_2 FILLER_89_1010 ();
 sg13g2_decap_8 FILLER_89_1017 ();
 sg13g2_decap_8 FILLER_89_1024 ();
 sg13g2_decap_8 FILLER_89_1031 ();
 sg13g2_decap_8 FILLER_89_1038 ();
 sg13g2_fill_2 FILLER_89_1045 ();
 sg13g2_decap_8 FILLER_89_1054 ();
 sg13g2_fill_2 FILLER_89_1061 ();
 sg13g2_fill_1 FILLER_89_1063 ();
 sg13g2_decap_8 FILLER_89_1070 ();
 sg13g2_decap_8 FILLER_89_1077 ();
 sg13g2_fill_2 FILLER_89_1084 ();
 sg13g2_fill_1 FILLER_89_1086 ();
 sg13g2_decap_8 FILLER_89_1100 ();
 sg13g2_decap_8 FILLER_89_1107 ();
 sg13g2_decap_8 FILLER_89_1114 ();
 sg13g2_decap_8 FILLER_89_1121 ();
 sg13g2_decap_8 FILLER_89_1128 ();
 sg13g2_decap_4 FILLER_89_1135 ();
 sg13g2_decap_8 FILLER_89_1144 ();
 sg13g2_decap_8 FILLER_89_1151 ();
 sg13g2_decap_8 FILLER_89_1158 ();
 sg13g2_decap_8 FILLER_89_1165 ();
 sg13g2_decap_8 FILLER_89_1172 ();
 sg13g2_decap_4 FILLER_89_1179 ();
 sg13g2_decap_8 FILLER_89_1208 ();
 sg13g2_fill_2 FILLER_89_1215 ();
 sg13g2_fill_1 FILLER_89_1217 ();
 sg13g2_decap_8 FILLER_89_1222 ();
 sg13g2_decap_8 FILLER_89_1229 ();
 sg13g2_decap_8 FILLER_89_1240 ();
 sg13g2_decap_4 FILLER_89_1247 ();
 sg13g2_decap_8 FILLER_89_1259 ();
 sg13g2_decap_8 FILLER_89_1266 ();
 sg13g2_decap_8 FILLER_89_1273 ();
 sg13g2_decap_8 FILLER_89_1280 ();
 sg13g2_decap_8 FILLER_89_1287 ();
 sg13g2_decap_8 FILLER_89_1294 ();
 sg13g2_decap_8 FILLER_89_1301 ();
 sg13g2_decap_4 FILLER_89_1308 ();
 sg13g2_fill_1 FILLER_89_1312 ();
 sg13g2_decap_8 FILLER_89_1317 ();
 sg13g2_decap_8 FILLER_89_1324 ();
 sg13g2_decap_8 FILLER_89_1331 ();
 sg13g2_fill_1 FILLER_89_1338 ();
 sg13g2_decap_8 FILLER_89_1343 ();
 sg13g2_fill_2 FILLER_89_1350 ();
 sg13g2_fill_1 FILLER_89_1352 ();
 sg13g2_fill_2 FILLER_89_1358 ();
 sg13g2_decap_8 FILLER_89_1399 ();
 sg13g2_decap_8 FILLER_89_1406 ();
 sg13g2_decap_8 FILLER_89_1413 ();
 sg13g2_decap_8 FILLER_89_1420 ();
 sg13g2_decap_8 FILLER_89_1427 ();
 sg13g2_decap_8 FILLER_89_1434 ();
 sg13g2_decap_4 FILLER_89_1441 ();
 sg13g2_fill_1 FILLER_89_1445 ();
 sg13g2_decap_8 FILLER_89_1480 ();
 sg13g2_decap_8 FILLER_89_1487 ();
 sg13g2_decap_8 FILLER_89_1494 ();
 sg13g2_decap_8 FILLER_89_1501 ();
 sg13g2_decap_8 FILLER_89_1521 ();
 sg13g2_decap_8 FILLER_89_1528 ();
 sg13g2_decap_4 FILLER_89_1535 ();
 sg13g2_fill_2 FILLER_89_1539 ();
 sg13g2_decap_8 FILLER_89_1550 ();
 sg13g2_decap_4 FILLER_89_1557 ();
 sg13g2_decap_8 FILLER_89_1566 ();
 sg13g2_fill_2 FILLER_89_1573 ();
 sg13g2_fill_1 FILLER_89_1591 ();
 sg13g2_fill_2 FILLER_89_1608 ();
 sg13g2_decap_8 FILLER_89_1619 ();
 sg13g2_decap_8 FILLER_89_1626 ();
 sg13g2_decap_8 FILLER_89_1633 ();
 sg13g2_decap_8 FILLER_89_1640 ();
 sg13g2_decap_8 FILLER_89_1647 ();
 sg13g2_decap_4 FILLER_89_1654 ();
 sg13g2_fill_1 FILLER_89_1658 ();
 sg13g2_fill_1 FILLER_89_1663 ();
 sg13g2_decap_8 FILLER_89_1668 ();
 sg13g2_fill_1 FILLER_89_1675 ();
 sg13g2_decap_8 FILLER_89_1684 ();
 sg13g2_decap_8 FILLER_89_1691 ();
 sg13g2_fill_2 FILLER_89_1698 ();
 sg13g2_decap_8 FILLER_89_1704 ();
 sg13g2_decap_8 FILLER_89_1711 ();
 sg13g2_decap_8 FILLER_89_1718 ();
 sg13g2_decap_8 FILLER_89_1725 ();
 sg13g2_decap_8 FILLER_89_1732 ();
 sg13g2_decap_8 FILLER_89_1739 ();
 sg13g2_decap_8 FILLER_89_1746 ();
 sg13g2_decap_8 FILLER_89_1753 ();
 sg13g2_decap_8 FILLER_89_1760 ();
 sg13g2_fill_1 FILLER_89_1767 ();
 sg13g2_decap_8 FILLER_90_0 ();
 sg13g2_decap_8 FILLER_90_7 ();
 sg13g2_fill_1 FILLER_90_14 ();
 sg13g2_decap_8 FILLER_90_35 ();
 sg13g2_decap_4 FILLER_90_42 ();
 sg13g2_fill_2 FILLER_90_58 ();
 sg13g2_fill_1 FILLER_90_60 ();
 sg13g2_decap_8 FILLER_90_65 ();
 sg13g2_decap_4 FILLER_90_86 ();
 sg13g2_fill_2 FILLER_90_90 ();
 sg13g2_fill_1 FILLER_90_102 ();
 sg13g2_decap_8 FILLER_90_111 ();
 sg13g2_decap_8 FILLER_90_118 ();
 sg13g2_decap_8 FILLER_90_125 ();
 sg13g2_fill_2 FILLER_90_132 ();
 sg13g2_fill_1 FILLER_90_134 ();
 sg13g2_fill_2 FILLER_90_139 ();
 sg13g2_decap_8 FILLER_90_149 ();
 sg13g2_decap_8 FILLER_90_156 ();
 sg13g2_fill_1 FILLER_90_163 ();
 sg13g2_decap_8 FILLER_90_174 ();
 sg13g2_fill_1 FILLER_90_181 ();
 sg13g2_decap_8 FILLER_90_189 ();
 sg13g2_decap_8 FILLER_90_196 ();
 sg13g2_decap_8 FILLER_90_203 ();
 sg13g2_decap_8 FILLER_90_210 ();
 sg13g2_decap_4 FILLER_90_217 ();
 sg13g2_fill_2 FILLER_90_221 ();
 sg13g2_decap_8 FILLER_90_231 ();
 sg13g2_decap_8 FILLER_90_242 ();
 sg13g2_decap_8 FILLER_90_249 ();
 sg13g2_decap_8 FILLER_90_256 ();
 sg13g2_decap_8 FILLER_90_263 ();
 sg13g2_decap_4 FILLER_90_270 ();
 sg13g2_decap_8 FILLER_90_295 ();
 sg13g2_decap_8 FILLER_90_302 ();
 sg13g2_decap_8 FILLER_90_309 ();
 sg13g2_decap_8 FILLER_90_316 ();
 sg13g2_decap_8 FILLER_90_323 ();
 sg13g2_fill_2 FILLER_90_330 ();
 sg13g2_decap_8 FILLER_90_348 ();
 sg13g2_decap_4 FILLER_90_355 ();
 sg13g2_fill_1 FILLER_90_359 ();
 sg13g2_decap_8 FILLER_90_368 ();
 sg13g2_decap_8 FILLER_90_375 ();
 sg13g2_decap_8 FILLER_90_382 ();
 sg13g2_decap_8 FILLER_90_389 ();
 sg13g2_decap_4 FILLER_90_396 ();
 sg13g2_fill_2 FILLER_90_407 ();
 sg13g2_fill_1 FILLER_90_409 ();
 sg13g2_decap_8 FILLER_90_414 ();
 sg13g2_decap_8 FILLER_90_421 ();
 sg13g2_decap_8 FILLER_90_428 ();
 sg13g2_decap_8 FILLER_90_435 ();
 sg13g2_decap_8 FILLER_90_442 ();
 sg13g2_fill_1 FILLER_90_449 ();
 sg13g2_decap_8 FILLER_90_474 ();
 sg13g2_decap_8 FILLER_90_481 ();
 sg13g2_decap_4 FILLER_90_488 ();
 sg13g2_fill_2 FILLER_90_492 ();
 sg13g2_fill_2 FILLER_90_504 ();
 sg13g2_fill_2 FILLER_90_511 ();
 sg13g2_fill_1 FILLER_90_513 ();
 sg13g2_fill_2 FILLER_90_518 ();
 sg13g2_decap_8 FILLER_90_525 ();
 sg13g2_decap_8 FILLER_90_532 ();
 sg13g2_decap_8 FILLER_90_539 ();
 sg13g2_fill_2 FILLER_90_546 ();
 sg13g2_decap_8 FILLER_90_556 ();
 sg13g2_decap_8 FILLER_90_563 ();
 sg13g2_decap_8 FILLER_90_570 ();
 sg13g2_fill_2 FILLER_90_577 ();
 sg13g2_fill_1 FILLER_90_579 ();
 sg13g2_decap_8 FILLER_90_623 ();
 sg13g2_fill_2 FILLER_90_630 ();
 sg13g2_fill_1 FILLER_90_632 ();
 sg13g2_decap_8 FILLER_90_647 ();
 sg13g2_decap_8 FILLER_90_654 ();
 sg13g2_decap_8 FILLER_90_661 ();
 sg13g2_decap_8 FILLER_90_668 ();
 sg13g2_decap_8 FILLER_90_675 ();
 sg13g2_fill_1 FILLER_90_682 ();
 sg13g2_decap_8 FILLER_90_693 ();
 sg13g2_decap_8 FILLER_90_700 ();
 sg13g2_decap_8 FILLER_90_707 ();
 sg13g2_decap_8 FILLER_90_714 ();
 sg13g2_decap_8 FILLER_90_721 ();
 sg13g2_decap_8 FILLER_90_728 ();
 sg13g2_decap_8 FILLER_90_735 ();
 sg13g2_decap_8 FILLER_90_742 ();
 sg13g2_fill_1 FILLER_90_754 ();
 sg13g2_decap_8 FILLER_90_758 ();
 sg13g2_decap_8 FILLER_90_765 ();
 sg13g2_decap_8 FILLER_90_772 ();
 sg13g2_fill_2 FILLER_90_779 ();
 sg13g2_decap_8 FILLER_90_785 ();
 sg13g2_decap_8 FILLER_90_792 ();
 sg13g2_decap_8 FILLER_90_799 ();
 sg13g2_decap_4 FILLER_90_806 ();
 sg13g2_fill_1 FILLER_90_810 ();
 sg13g2_decap_8 FILLER_90_820 ();
 sg13g2_decap_8 FILLER_90_827 ();
 sg13g2_decap_8 FILLER_90_843 ();
 sg13g2_decap_8 FILLER_90_850 ();
 sg13g2_decap_8 FILLER_90_857 ();
 sg13g2_decap_8 FILLER_90_864 ();
 sg13g2_decap_8 FILLER_90_871 ();
 sg13g2_decap_8 FILLER_90_878 ();
 sg13g2_decap_8 FILLER_90_885 ();
 sg13g2_decap_8 FILLER_90_892 ();
 sg13g2_decap_4 FILLER_90_899 ();
 sg13g2_decap_4 FILLER_90_909 ();
 sg13g2_fill_2 FILLER_90_913 ();
 sg13g2_decap_4 FILLER_90_928 ();
 sg13g2_fill_2 FILLER_90_932 ();
 sg13g2_decap_4 FILLER_90_988 ();
 sg13g2_decap_8 FILLER_90_1028 ();
 sg13g2_decap_8 FILLER_90_1035 ();
 sg13g2_decap_8 FILLER_90_1042 ();
 sg13g2_decap_8 FILLER_90_1049 ();
 sg13g2_decap_8 FILLER_90_1056 ();
 sg13g2_fill_2 FILLER_90_1063 ();
 sg13g2_fill_1 FILLER_90_1065 ();
 sg13g2_decap_8 FILLER_90_1075 ();
 sg13g2_decap_4 FILLER_90_1082 ();
 sg13g2_fill_2 FILLER_90_1086 ();
 sg13g2_decap_4 FILLER_90_1114 ();
 sg13g2_fill_2 FILLER_90_1118 ();
 sg13g2_decap_8 FILLER_90_1171 ();
 sg13g2_decap_8 FILLER_90_1182 ();
 sg13g2_decap_8 FILLER_90_1189 ();
 sg13g2_decap_8 FILLER_90_1196 ();
 sg13g2_decap_8 FILLER_90_1203 ();
 sg13g2_decap_8 FILLER_90_1210 ();
 sg13g2_decap_8 FILLER_90_1217 ();
 sg13g2_decap_8 FILLER_90_1224 ();
 sg13g2_decap_8 FILLER_90_1231 ();
 sg13g2_decap_8 FILLER_90_1238 ();
 sg13g2_decap_8 FILLER_90_1245 ();
 sg13g2_decap_8 FILLER_90_1252 ();
 sg13g2_decap_8 FILLER_90_1259 ();
 sg13g2_decap_8 FILLER_90_1266 ();
 sg13g2_fill_1 FILLER_90_1273 ();
 sg13g2_fill_2 FILLER_90_1282 ();
 sg13g2_fill_1 FILLER_90_1284 ();
 sg13g2_fill_2 FILLER_90_1294 ();
 sg13g2_decap_8 FILLER_90_1303 ();
 sg13g2_decap_8 FILLER_90_1310 ();
 sg13g2_decap_8 FILLER_90_1317 ();
 sg13g2_decap_8 FILLER_90_1324 ();
 sg13g2_decap_8 FILLER_90_1331 ();
 sg13g2_decap_4 FILLER_90_1338 ();
 sg13g2_fill_1 FILLER_90_1342 ();
 sg13g2_decap_8 FILLER_90_1347 ();
 sg13g2_decap_4 FILLER_90_1354 ();
 sg13g2_decap_8 FILLER_90_1362 ();
 sg13g2_decap_8 FILLER_90_1374 ();
 sg13g2_decap_8 FILLER_90_1381 ();
 sg13g2_decap_8 FILLER_90_1388 ();
 sg13g2_decap_8 FILLER_90_1395 ();
 sg13g2_decap_8 FILLER_90_1402 ();
 sg13g2_decap_8 FILLER_90_1409 ();
 sg13g2_decap_8 FILLER_90_1416 ();
 sg13g2_decap_8 FILLER_90_1423 ();
 sg13g2_decap_8 FILLER_90_1430 ();
 sg13g2_fill_2 FILLER_90_1437 ();
 sg13g2_fill_1 FILLER_90_1439 ();
 sg13g2_fill_2 FILLER_90_1445 ();
 sg13g2_fill_1 FILLER_90_1447 ();
 sg13g2_decap_8 FILLER_90_1460 ();
 sg13g2_decap_8 FILLER_90_1467 ();
 sg13g2_decap_8 FILLER_90_1474 ();
 sg13g2_decap_8 FILLER_90_1481 ();
 sg13g2_decap_8 FILLER_90_1488 ();
 sg13g2_decap_8 FILLER_90_1495 ();
 sg13g2_decap_8 FILLER_90_1502 ();
 sg13g2_decap_8 FILLER_90_1517 ();
 sg13g2_decap_8 FILLER_90_1524 ();
 sg13g2_decap_8 FILLER_90_1531 ();
 sg13g2_decap_8 FILLER_90_1538 ();
 sg13g2_decap_8 FILLER_90_1545 ();
 sg13g2_decap_4 FILLER_90_1552 ();
 sg13g2_fill_1 FILLER_90_1556 ();
 sg13g2_fill_1 FILLER_90_1583 ();
 sg13g2_fill_2 FILLER_90_1603 ();
 sg13g2_fill_2 FILLER_90_1608 ();
 sg13g2_decap_8 FILLER_90_1619 ();
 sg13g2_decap_8 FILLER_90_1626 ();
 sg13g2_decap_8 FILLER_90_1633 ();
 sg13g2_decap_8 FILLER_90_1640 ();
 sg13g2_fill_1 FILLER_90_1647 ();
 sg13g2_decap_4 FILLER_90_1674 ();
 sg13g2_fill_1 FILLER_90_1678 ();
 sg13g2_decap_4 FILLER_90_1682 ();
 sg13g2_decap_8 FILLER_90_1699 ();
 sg13g2_fill_1 FILLER_90_1706 ();
 sg13g2_decap_8 FILLER_90_1712 ();
 sg13g2_decap_4 FILLER_90_1719 ();
 sg13g2_fill_1 FILLER_90_1723 ();
 sg13g2_decap_8 FILLER_90_1750 ();
 sg13g2_decap_8 FILLER_90_1757 ();
 sg13g2_decap_4 FILLER_90_1764 ();
 sg13g2_decap_8 FILLER_91_0 ();
 sg13g2_decap_8 FILLER_91_7 ();
 sg13g2_fill_2 FILLER_91_14 ();
 sg13g2_fill_1 FILLER_91_16 ();
 sg13g2_decap_8 FILLER_91_35 ();
 sg13g2_decap_4 FILLER_91_42 ();
 sg13g2_fill_2 FILLER_91_46 ();
 sg13g2_fill_2 FILLER_91_60 ();
 sg13g2_fill_1 FILLER_91_62 ();
 sg13g2_decap_8 FILLER_91_71 ();
 sg13g2_decap_8 FILLER_91_78 ();
 sg13g2_decap_8 FILLER_91_118 ();
 sg13g2_fill_1 FILLER_91_125 ();
 sg13g2_decap_4 FILLER_91_158 ();
 sg13g2_fill_2 FILLER_91_162 ();
 sg13g2_decap_8 FILLER_91_172 ();
 sg13g2_decap_8 FILLER_91_179 ();
 sg13g2_decap_8 FILLER_91_186 ();
 sg13g2_decap_8 FILLER_91_193 ();
 sg13g2_decap_8 FILLER_91_200 ();
 sg13g2_decap_8 FILLER_91_207 ();
 sg13g2_decap_8 FILLER_91_214 ();
 sg13g2_decap_8 FILLER_91_221 ();
 sg13g2_decap_8 FILLER_91_228 ();
 sg13g2_decap_8 FILLER_91_235 ();
 sg13g2_decap_8 FILLER_91_242 ();
 sg13g2_decap_8 FILLER_91_249 ();
 sg13g2_decap_8 FILLER_91_256 ();
 sg13g2_decap_8 FILLER_91_263 ();
 sg13g2_decap_8 FILLER_91_270 ();
 sg13g2_decap_8 FILLER_91_277 ();
 sg13g2_decap_8 FILLER_91_284 ();
 sg13g2_decap_8 FILLER_91_291 ();
 sg13g2_decap_8 FILLER_91_298 ();
 sg13g2_decap_8 FILLER_91_305 ();
 sg13g2_decap_8 FILLER_91_312 ();
 sg13g2_decap_8 FILLER_91_319 ();
 sg13g2_fill_2 FILLER_91_326 ();
 sg13g2_fill_1 FILLER_91_328 ();
 sg13g2_fill_2 FILLER_91_345 ();
 sg13g2_decap_8 FILLER_91_354 ();
 sg13g2_decap_8 FILLER_91_361 ();
 sg13g2_decap_8 FILLER_91_368 ();
 sg13g2_decap_8 FILLER_91_375 ();
 sg13g2_decap_8 FILLER_91_382 ();
 sg13g2_decap_8 FILLER_91_389 ();
 sg13g2_decap_8 FILLER_91_396 ();
 sg13g2_decap_8 FILLER_91_406 ();
 sg13g2_decap_8 FILLER_91_413 ();
 sg13g2_decap_8 FILLER_91_420 ();
 sg13g2_decap_8 FILLER_91_427 ();
 sg13g2_decap_8 FILLER_91_434 ();
 sg13g2_decap_8 FILLER_91_441 ();
 sg13g2_decap_4 FILLER_91_448 ();
 sg13g2_decap_8 FILLER_91_466 ();
 sg13g2_decap_8 FILLER_91_481 ();
 sg13g2_decap_4 FILLER_91_488 ();
 sg13g2_fill_2 FILLER_91_492 ();
 sg13g2_decap_8 FILLER_91_498 ();
 sg13g2_decap_4 FILLER_91_505 ();
 sg13g2_decap_8 FILLER_91_517 ();
 sg13g2_decap_8 FILLER_91_524 ();
 sg13g2_fill_2 FILLER_91_531 ();
 sg13g2_fill_1 FILLER_91_547 ();
 sg13g2_decap_8 FILLER_91_558 ();
 sg13g2_decap_8 FILLER_91_565 ();
 sg13g2_decap_8 FILLER_91_572 ();
 sg13g2_decap_8 FILLER_91_579 ();
 sg13g2_fill_2 FILLER_91_586 ();
 sg13g2_fill_2 FILLER_91_593 ();
 sg13g2_decap_4 FILLER_91_600 ();
 sg13g2_fill_2 FILLER_91_604 ();
 sg13g2_decap_4 FILLER_91_619 ();
 sg13g2_fill_1 FILLER_91_623 ();
 sg13g2_decap_4 FILLER_91_652 ();
 sg13g2_fill_1 FILLER_91_656 ();
 sg13g2_fill_1 FILLER_91_692 ();
 sg13g2_decap_8 FILLER_91_706 ();
 sg13g2_decap_8 FILLER_91_713 ();
 sg13g2_decap_8 FILLER_91_720 ();
 sg13g2_decap_8 FILLER_91_727 ();
 sg13g2_decap_4 FILLER_91_734 ();
 sg13g2_fill_1 FILLER_91_738 ();
 sg13g2_decap_8 FILLER_91_743 ();
 sg13g2_decap_8 FILLER_91_755 ();
 sg13g2_decap_8 FILLER_91_762 ();
 sg13g2_decap_8 FILLER_91_769 ();
 sg13g2_decap_8 FILLER_91_776 ();
 sg13g2_decap_8 FILLER_91_783 ();
 sg13g2_decap_8 FILLER_91_790 ();
 sg13g2_decap_4 FILLER_91_797 ();
 sg13g2_decap_8 FILLER_91_805 ();
 sg13g2_decap_8 FILLER_91_812 ();
 sg13g2_fill_2 FILLER_91_819 ();
 sg13g2_fill_1 FILLER_91_834 ();
 sg13g2_decap_8 FILLER_91_861 ();
 sg13g2_decap_8 FILLER_91_868 ();
 sg13g2_decap_8 FILLER_91_875 ();
 sg13g2_decap_8 FILLER_91_882 ();
 sg13g2_decap_4 FILLER_91_928 ();
 sg13g2_fill_2 FILLER_91_932 ();
 sg13g2_fill_2 FILLER_91_944 ();
 sg13g2_decap_8 FILLER_91_963 ();
 sg13g2_decap_8 FILLER_91_970 ();
 sg13g2_decap_8 FILLER_91_977 ();
 sg13g2_decap_4 FILLER_91_984 ();
 sg13g2_decap_8 FILLER_91_1016 ();
 sg13g2_decap_8 FILLER_91_1023 ();
 sg13g2_decap_8 FILLER_91_1030 ();
 sg13g2_decap_8 FILLER_91_1037 ();
 sg13g2_decap_8 FILLER_91_1044 ();
 sg13g2_decap_8 FILLER_91_1051 ();
 sg13g2_decap_8 FILLER_91_1058 ();
 sg13g2_decap_4 FILLER_91_1065 ();
 sg13g2_fill_1 FILLER_91_1073 ();
 sg13g2_decap_8 FILLER_91_1079 ();
 sg13g2_decap_8 FILLER_91_1086 ();
 sg13g2_decap_4 FILLER_91_1093 ();
 sg13g2_fill_2 FILLER_91_1097 ();
 sg13g2_decap_8 FILLER_91_1103 ();
 sg13g2_decap_8 FILLER_91_1110 ();
 sg13g2_fill_2 FILLER_91_1117 ();
 sg13g2_fill_1 FILLER_91_1119 ();
 sg13g2_fill_1 FILLER_91_1137 ();
 sg13g2_decap_8 FILLER_91_1148 ();
 sg13g2_fill_1 FILLER_91_1155 ();
 sg13g2_decap_8 FILLER_91_1160 ();
 sg13g2_decap_8 FILLER_91_1167 ();
 sg13g2_decap_4 FILLER_91_1174 ();
 sg13g2_decap_8 FILLER_91_1191 ();
 sg13g2_decap_8 FILLER_91_1198 ();
 sg13g2_decap_8 FILLER_91_1205 ();
 sg13g2_decap_4 FILLER_91_1212 ();
 sg13g2_fill_1 FILLER_91_1216 ();
 sg13g2_decap_8 FILLER_91_1225 ();
 sg13g2_decap_8 FILLER_91_1232 ();
 sg13g2_decap_8 FILLER_91_1239 ();
 sg13g2_decap_8 FILLER_91_1246 ();
 sg13g2_decap_8 FILLER_91_1253 ();
 sg13g2_decap_8 FILLER_91_1260 ();
 sg13g2_decap_8 FILLER_91_1267 ();
 sg13g2_fill_1 FILLER_91_1274 ();
 sg13g2_decap_8 FILLER_91_1298 ();
 sg13g2_decap_8 FILLER_91_1305 ();
 sg13g2_decap_4 FILLER_91_1312 ();
 sg13g2_fill_2 FILLER_91_1316 ();
 sg13g2_decap_4 FILLER_91_1367 ();
 sg13g2_decap_8 FILLER_91_1384 ();
 sg13g2_decap_4 FILLER_91_1391 ();
 sg13g2_fill_2 FILLER_91_1395 ();
 sg13g2_decap_8 FILLER_91_1401 ();
 sg13g2_decap_8 FILLER_91_1408 ();
 sg13g2_decap_4 FILLER_91_1415 ();
 sg13g2_fill_1 FILLER_91_1419 ();
 sg13g2_decap_8 FILLER_91_1433 ();
 sg13g2_decap_8 FILLER_91_1440 ();
 sg13g2_decap_4 FILLER_91_1447 ();
 sg13g2_decap_8 FILLER_91_1454 ();
 sg13g2_decap_8 FILLER_91_1461 ();
 sg13g2_decap_8 FILLER_91_1468 ();
 sg13g2_decap_8 FILLER_91_1475 ();
 sg13g2_decap_4 FILLER_91_1482 ();
 sg13g2_decap_8 FILLER_91_1490 ();
 sg13g2_decap_8 FILLER_91_1497 ();
 sg13g2_decap_4 FILLER_91_1504 ();
 sg13g2_fill_1 FILLER_91_1508 ();
 sg13g2_decap_8 FILLER_91_1517 ();
 sg13g2_decap_8 FILLER_91_1524 ();
 sg13g2_decap_8 FILLER_91_1531 ();
 sg13g2_decap_8 FILLER_91_1538 ();
 sg13g2_decap_8 FILLER_91_1545 ();
 sg13g2_decap_8 FILLER_91_1552 ();
 sg13g2_decap_8 FILLER_91_1630 ();
 sg13g2_decap_8 FILLER_91_1637 ();
 sg13g2_decap_8 FILLER_91_1644 ();
 sg13g2_decap_8 FILLER_91_1651 ();
 sg13g2_decap_8 FILLER_91_1658 ();
 sg13g2_fill_2 FILLER_91_1665 ();
 sg13g2_fill_1 FILLER_91_1667 ();
 sg13g2_fill_1 FILLER_91_1686 ();
 sg13g2_decap_8 FILLER_91_1700 ();
 sg13g2_decap_8 FILLER_91_1707 ();
 sg13g2_decap_8 FILLER_91_1714 ();
 sg13g2_decap_8 FILLER_91_1721 ();
 sg13g2_fill_2 FILLER_91_1728 ();
 sg13g2_fill_1 FILLER_91_1730 ();
 sg13g2_fill_2 FILLER_91_1744 ();
 sg13g2_decap_8 FILLER_91_1759 ();
 sg13g2_fill_2 FILLER_91_1766 ();
 sg13g2_decap_8 FILLER_92_0 ();
 sg13g2_decap_8 FILLER_92_7 ();
 sg13g2_decap_8 FILLER_92_14 ();
 sg13g2_decap_4 FILLER_92_21 ();
 sg13g2_fill_1 FILLER_92_25 ();
 sg13g2_decap_8 FILLER_92_31 ();
 sg13g2_decap_4 FILLER_92_38 ();
 sg13g2_fill_2 FILLER_92_42 ();
 sg13g2_decap_8 FILLER_92_48 ();
 sg13g2_decap_8 FILLER_92_55 ();
 sg13g2_decap_8 FILLER_92_62 ();
 sg13g2_decap_8 FILLER_92_69 ();
 sg13g2_decap_8 FILLER_92_76 ();
 sg13g2_decap_8 FILLER_92_83 ();
 sg13g2_decap_8 FILLER_92_90 ();
 sg13g2_decap_8 FILLER_92_97 ();
 sg13g2_decap_8 FILLER_92_116 ();
 sg13g2_decap_8 FILLER_92_123 ();
 sg13g2_decap_8 FILLER_92_130 ();
 sg13g2_fill_2 FILLER_92_137 ();
 sg13g2_fill_1 FILLER_92_139 ();
 sg13g2_fill_1 FILLER_92_152 ();
 sg13g2_decap_8 FILLER_92_160 ();
 sg13g2_decap_8 FILLER_92_167 ();
 sg13g2_decap_8 FILLER_92_174 ();
 sg13g2_decap_8 FILLER_92_181 ();
 sg13g2_decap_8 FILLER_92_188 ();
 sg13g2_decap_8 FILLER_92_195 ();
 sg13g2_decap_8 FILLER_92_202 ();
 sg13g2_decap_8 FILLER_92_209 ();
 sg13g2_fill_2 FILLER_92_216 ();
 sg13g2_fill_1 FILLER_92_218 ();
 sg13g2_decap_8 FILLER_92_236 ();
 sg13g2_decap_8 FILLER_92_243 ();
 sg13g2_decap_8 FILLER_92_250 ();
 sg13g2_fill_2 FILLER_92_257 ();
 sg13g2_fill_1 FILLER_92_259 ();
 sg13g2_decap_8 FILLER_92_268 ();
 sg13g2_decap_8 FILLER_92_275 ();
 sg13g2_decap_8 FILLER_92_282 ();
 sg13g2_decap_8 FILLER_92_289 ();
 sg13g2_decap_8 FILLER_92_296 ();
 sg13g2_fill_2 FILLER_92_303 ();
 sg13g2_fill_1 FILLER_92_305 ();
 sg13g2_decap_8 FILLER_92_314 ();
 sg13g2_decap_8 FILLER_92_321 ();
 sg13g2_fill_1 FILLER_92_328 ();
 sg13g2_fill_2 FILLER_92_337 ();
 sg13g2_fill_1 FILLER_92_339 ();
 sg13g2_decap_8 FILLER_92_357 ();
 sg13g2_decap_8 FILLER_92_364 ();
 sg13g2_decap_8 FILLER_92_371 ();
 sg13g2_fill_2 FILLER_92_378 ();
 sg13g2_decap_4 FILLER_92_392 ();
 sg13g2_fill_2 FILLER_92_396 ();
 sg13g2_decap_8 FILLER_92_402 ();
 sg13g2_decap_8 FILLER_92_409 ();
 sg13g2_decap_4 FILLER_92_416 ();
 sg13g2_fill_2 FILLER_92_420 ();
 sg13g2_decap_8 FILLER_92_427 ();
 sg13g2_decap_8 FILLER_92_434 ();
 sg13g2_decap_8 FILLER_92_441 ();
 sg13g2_decap_8 FILLER_92_448 ();
 sg13g2_decap_8 FILLER_92_455 ();
 sg13g2_fill_2 FILLER_92_462 ();
 sg13g2_fill_1 FILLER_92_464 ();
 sg13g2_decap_8 FILLER_92_473 ();
 sg13g2_decap_8 FILLER_92_480 ();
 sg13g2_decap_8 FILLER_92_487 ();
 sg13g2_decap_8 FILLER_92_494 ();
 sg13g2_decap_8 FILLER_92_501 ();
 sg13g2_decap_8 FILLER_92_513 ();
 sg13g2_decap_8 FILLER_92_520 ();
 sg13g2_decap_8 FILLER_92_527 ();
 sg13g2_fill_1 FILLER_92_534 ();
 sg13g2_decap_8 FILLER_92_556 ();
 sg13g2_decap_8 FILLER_92_563 ();
 sg13g2_decap_8 FILLER_92_570 ();
 sg13g2_decap_4 FILLER_92_577 ();
 sg13g2_fill_1 FILLER_92_581 ();
 sg13g2_decap_8 FILLER_92_588 ();
 sg13g2_decap_8 FILLER_92_595 ();
 sg13g2_decap_8 FILLER_92_602 ();
 sg13g2_decap_8 FILLER_92_609 ();
 sg13g2_decap_8 FILLER_92_616 ();
 sg13g2_decap_8 FILLER_92_623 ();
 sg13g2_decap_8 FILLER_92_630 ();
 sg13g2_decap_8 FILLER_92_637 ();
 sg13g2_decap_8 FILLER_92_644 ();
 sg13g2_fill_1 FILLER_92_651 ();
 sg13g2_fill_2 FILLER_92_673 ();
 sg13g2_fill_1 FILLER_92_675 ();
 sg13g2_decap_8 FILLER_92_684 ();
 sg13g2_fill_2 FILLER_92_691 ();
 sg13g2_decap_8 FILLER_92_702 ();
 sg13g2_decap_8 FILLER_92_709 ();
 sg13g2_decap_4 FILLER_92_716 ();
 sg13g2_fill_2 FILLER_92_720 ();
 sg13g2_decap_8 FILLER_92_731 ();
 sg13g2_decap_8 FILLER_92_738 ();
 sg13g2_decap_4 FILLER_92_745 ();
 sg13g2_decap_4 FILLER_92_755 ();
 sg13g2_fill_2 FILLER_92_759 ();
 sg13g2_decap_8 FILLER_92_766 ();
 sg13g2_decap_8 FILLER_92_773 ();
 sg13g2_decap_8 FILLER_92_780 ();
 sg13g2_fill_2 FILLER_92_787 ();
 sg13g2_fill_1 FILLER_92_789 ();
 sg13g2_decap_8 FILLER_92_816 ();
 sg13g2_decap_8 FILLER_92_823 ();
 sg13g2_decap_8 FILLER_92_830 ();
 sg13g2_decap_8 FILLER_92_837 ();
 sg13g2_fill_2 FILLER_92_844 ();
 sg13g2_decap_8 FILLER_92_850 ();
 sg13g2_decap_8 FILLER_92_857 ();
 sg13g2_decap_8 FILLER_92_882 ();
 sg13g2_decap_8 FILLER_92_889 ();
 sg13g2_decap_4 FILLER_92_896 ();
 sg13g2_decap_8 FILLER_92_904 ();
 sg13g2_decap_4 FILLER_92_911 ();
 sg13g2_fill_1 FILLER_92_915 ();
 sg13g2_decap_8 FILLER_92_924 ();
 sg13g2_decap_8 FILLER_92_931 ();
 sg13g2_decap_8 FILLER_92_938 ();
 sg13g2_decap_8 FILLER_92_945 ();
 sg13g2_decap_8 FILLER_92_952 ();
 sg13g2_decap_8 FILLER_92_959 ();
 sg13g2_decap_8 FILLER_92_966 ();
 sg13g2_decap_8 FILLER_92_973 ();
 sg13g2_decap_8 FILLER_92_980 ();
 sg13g2_decap_4 FILLER_92_987 ();
 sg13g2_decap_8 FILLER_92_1013 ();
 sg13g2_decap_8 FILLER_92_1020 ();
 sg13g2_decap_4 FILLER_92_1027 ();
 sg13g2_fill_1 FILLER_92_1031 ();
 sg13g2_decap_8 FILLER_92_1045 ();
 sg13g2_decap_4 FILLER_92_1052 ();
 sg13g2_fill_2 FILLER_92_1056 ();
 sg13g2_decap_8 FILLER_92_1083 ();
 sg13g2_decap_8 FILLER_92_1090 ();
 sg13g2_decap_8 FILLER_92_1097 ();
 sg13g2_decap_8 FILLER_92_1104 ();
 sg13g2_decap_8 FILLER_92_1111 ();
 sg13g2_decap_8 FILLER_92_1118 ();
 sg13g2_decap_8 FILLER_92_1125 ();
 sg13g2_decap_8 FILLER_92_1136 ();
 sg13g2_decap_8 FILLER_92_1143 ();
 sg13g2_fill_2 FILLER_92_1150 ();
 sg13g2_decap_8 FILLER_92_1156 ();
 sg13g2_fill_1 FILLER_92_1163 ();
 sg13g2_decap_4 FILLER_92_1172 ();
 sg13g2_decap_8 FILLER_92_1179 ();
 sg13g2_decap_8 FILLER_92_1186 ();
 sg13g2_decap_8 FILLER_92_1193 ();
 sg13g2_decap_8 FILLER_92_1200 ();
 sg13g2_decap_8 FILLER_92_1207 ();
 sg13g2_decap_4 FILLER_92_1214 ();
 sg13g2_fill_1 FILLER_92_1218 ();
 sg13g2_decap_8 FILLER_92_1245 ();
 sg13g2_decap_8 FILLER_92_1252 ();
 sg13g2_decap_8 FILLER_92_1259 ();
 sg13g2_fill_1 FILLER_92_1266 ();
 sg13g2_decap_8 FILLER_92_1275 ();
 sg13g2_decap_4 FILLER_92_1282 ();
 sg13g2_fill_2 FILLER_92_1286 ();
 sg13g2_decap_8 FILLER_92_1291 ();
 sg13g2_decap_8 FILLER_92_1298 ();
 sg13g2_fill_2 FILLER_92_1305 ();
 sg13g2_fill_2 FILLER_92_1311 ();
 sg13g2_fill_1 FILLER_92_1313 ();
 sg13g2_decap_8 FILLER_92_1340 ();
 sg13g2_decap_8 FILLER_92_1347 ();
 sg13g2_decap_4 FILLER_92_1354 ();
 sg13g2_fill_2 FILLER_92_1358 ();
 sg13g2_fill_2 FILLER_92_1365 ();
 sg13g2_fill_1 FILLER_92_1367 ();
 sg13g2_decap_8 FILLER_92_1412 ();
 sg13g2_decap_8 FILLER_92_1432 ();
 sg13g2_decap_8 FILLER_92_1439 ();
 sg13g2_decap_8 FILLER_92_1446 ();
 sg13g2_fill_2 FILLER_92_1453 ();
 sg13g2_fill_1 FILLER_92_1455 ();
 sg13g2_decap_8 FILLER_92_1461 ();
 sg13g2_decap_4 FILLER_92_1468 ();
 sg13g2_fill_2 FILLER_92_1472 ();
 sg13g2_fill_2 FILLER_92_1478 ();
 sg13g2_fill_1 FILLER_92_1480 ();
 sg13g2_fill_2 FILLER_92_1485 ();
 sg13g2_fill_1 FILLER_92_1487 ();
 sg13g2_decap_8 FILLER_92_1496 ();
 sg13g2_decap_8 FILLER_92_1503 ();
 sg13g2_fill_1 FILLER_92_1510 ();
 sg13g2_fill_2 FILLER_92_1537 ();
 sg13g2_decap_8 FILLER_92_1547 ();
 sg13g2_decap_8 FILLER_92_1554 ();
 sg13g2_fill_2 FILLER_92_1561 ();
 sg13g2_decap_4 FILLER_92_1572 ();
 sg13g2_fill_1 FILLER_92_1576 ();
 sg13g2_decap_8 FILLER_92_1587 ();
 sg13g2_decap_8 FILLER_92_1594 ();
 sg13g2_fill_1 FILLER_92_1601 ();
 sg13g2_fill_2 FILLER_92_1608 ();
 sg13g2_decap_4 FILLER_92_1632 ();
 sg13g2_decap_8 FILLER_92_1640 ();
 sg13g2_decap_8 FILLER_92_1647 ();
 sg13g2_decap_8 FILLER_92_1654 ();
 sg13g2_decap_8 FILLER_92_1661 ();
 sg13g2_decap_8 FILLER_92_1668 ();
 sg13g2_decap_8 FILLER_92_1675 ();
 sg13g2_fill_1 FILLER_92_1687 ();
 sg13g2_decap_8 FILLER_92_1706 ();
 sg13g2_decap_8 FILLER_92_1713 ();
 sg13g2_decap_8 FILLER_92_1720 ();
 sg13g2_fill_1 FILLER_92_1727 ();
 sg13g2_decap_8 FILLER_92_1750 ();
 sg13g2_decap_8 FILLER_92_1757 ();
 sg13g2_decap_4 FILLER_92_1764 ();
 sg13g2_decap_8 FILLER_93_0 ();
 sg13g2_decap_8 FILLER_93_7 ();
 sg13g2_decap_8 FILLER_93_14 ();
 sg13g2_decap_8 FILLER_93_21 ();
 sg13g2_decap_4 FILLER_93_28 ();
 sg13g2_fill_2 FILLER_93_32 ();
 sg13g2_decap_8 FILLER_93_53 ();
 sg13g2_decap_4 FILLER_93_60 ();
 sg13g2_decap_8 FILLER_93_76 ();
 sg13g2_fill_2 FILLER_93_83 ();
 sg13g2_fill_1 FILLER_93_85 ();
 sg13g2_decap_8 FILLER_93_91 ();
 sg13g2_decap_8 FILLER_93_98 ();
 sg13g2_decap_8 FILLER_93_105 ();
 sg13g2_decap_8 FILLER_93_112 ();
 sg13g2_decap_8 FILLER_93_119 ();
 sg13g2_decap_8 FILLER_93_126 ();
 sg13g2_decap_4 FILLER_93_133 ();
 sg13g2_fill_2 FILLER_93_137 ();
 sg13g2_fill_2 FILLER_93_163 ();
 sg13g2_decap_8 FILLER_93_173 ();
 sg13g2_decap_8 FILLER_93_180 ();
 sg13g2_decap_8 FILLER_93_187 ();
 sg13g2_decap_8 FILLER_93_194 ();
 sg13g2_decap_8 FILLER_93_201 ();
 sg13g2_decap_4 FILLER_93_208 ();
 sg13g2_fill_2 FILLER_93_212 ();
 sg13g2_decap_8 FILLER_93_243 ();
 sg13g2_decap_4 FILLER_93_250 ();
 sg13g2_fill_2 FILLER_93_263 ();
 sg13g2_decap_8 FILLER_93_281 ();
 sg13g2_decap_8 FILLER_93_288 ();
 sg13g2_decap_8 FILLER_93_295 ();
 sg13g2_decap_8 FILLER_93_302 ();
 sg13g2_decap_8 FILLER_93_309 ();
 sg13g2_decap_8 FILLER_93_316 ();
 sg13g2_decap_8 FILLER_93_323 ();
 sg13g2_decap_8 FILLER_93_330 ();
 sg13g2_decap_8 FILLER_93_337 ();
 sg13g2_decap_8 FILLER_93_344 ();
 sg13g2_decap_8 FILLER_93_351 ();
 sg13g2_fill_2 FILLER_93_358 ();
 sg13g2_fill_1 FILLER_93_360 ();
 sg13g2_decap_8 FILLER_93_369 ();
 sg13g2_fill_1 FILLER_93_392 ();
 sg13g2_decap_4 FILLER_93_409 ();
 sg13g2_decap_8 FILLER_93_435 ();
 sg13g2_decap_8 FILLER_93_442 ();
 sg13g2_decap_8 FILLER_93_449 ();
 sg13g2_decap_8 FILLER_93_456 ();
 sg13g2_decap_8 FILLER_93_463 ();
 sg13g2_decap_8 FILLER_93_470 ();
 sg13g2_decap_4 FILLER_93_477 ();
 sg13g2_fill_2 FILLER_93_481 ();
 sg13g2_decap_8 FILLER_93_488 ();
 sg13g2_decap_8 FILLER_93_495 ();
 sg13g2_fill_2 FILLER_93_502 ();
 sg13g2_decap_8 FILLER_93_512 ();
 sg13g2_decap_8 FILLER_93_519 ();
 sg13g2_decap_8 FILLER_93_526 ();
 sg13g2_fill_1 FILLER_93_533 ();
 sg13g2_decap_8 FILLER_93_542 ();
 sg13g2_decap_8 FILLER_93_549 ();
 sg13g2_decap_8 FILLER_93_556 ();
 sg13g2_decap_8 FILLER_93_563 ();
 sg13g2_decap_8 FILLER_93_570 ();
 sg13g2_decap_8 FILLER_93_577 ();
 sg13g2_decap_8 FILLER_93_584 ();
 sg13g2_fill_2 FILLER_93_591 ();
 sg13g2_decap_8 FILLER_93_606 ();
 sg13g2_decap_8 FILLER_93_613 ();
 sg13g2_decap_8 FILLER_93_620 ();
 sg13g2_decap_8 FILLER_93_627 ();
 sg13g2_decap_8 FILLER_93_634 ();
 sg13g2_decap_8 FILLER_93_641 ();
 sg13g2_decap_8 FILLER_93_648 ();
 sg13g2_decap_4 FILLER_93_655 ();
 sg13g2_fill_2 FILLER_93_659 ();
 sg13g2_decap_8 FILLER_93_670 ();
 sg13g2_fill_2 FILLER_93_677 ();
 sg13g2_fill_1 FILLER_93_679 ();
 sg13g2_decap_8 FILLER_93_689 ();
 sg13g2_fill_2 FILLER_93_696 ();
 sg13g2_fill_1 FILLER_93_698 ();
 sg13g2_fill_2 FILLER_93_712 ();
 sg13g2_fill_1 FILLER_93_714 ();
 sg13g2_decap_4 FILLER_93_722 ();
 sg13g2_fill_1 FILLER_93_726 ();
 sg13g2_decap_8 FILLER_93_741 ();
 sg13g2_decap_8 FILLER_93_748 ();
 sg13g2_decap_4 FILLER_93_755 ();
 sg13g2_fill_1 FILLER_93_759 ();
 sg13g2_decap_8 FILLER_93_764 ();
 sg13g2_fill_2 FILLER_93_779 ();
 sg13g2_decap_8 FILLER_93_803 ();
 sg13g2_decap_8 FILLER_93_810 ();
 sg13g2_decap_8 FILLER_93_817 ();
 sg13g2_decap_8 FILLER_93_824 ();
 sg13g2_decap_8 FILLER_93_831 ();
 sg13g2_decap_8 FILLER_93_838 ();
 sg13g2_decap_8 FILLER_93_845 ();
 sg13g2_decap_8 FILLER_93_852 ();
 sg13g2_fill_1 FILLER_93_859 ();
 sg13g2_decap_8 FILLER_93_881 ();
 sg13g2_decap_8 FILLER_93_888 ();
 sg13g2_decap_8 FILLER_93_895 ();
 sg13g2_decap_8 FILLER_93_902 ();
 sg13g2_decap_8 FILLER_93_909 ();
 sg13g2_decap_8 FILLER_93_916 ();
 sg13g2_decap_8 FILLER_93_923 ();
 sg13g2_decap_8 FILLER_93_930 ();
 sg13g2_decap_8 FILLER_93_945 ();
 sg13g2_decap_8 FILLER_93_952 ();
 sg13g2_fill_1 FILLER_93_959 ();
 sg13g2_decap_8 FILLER_93_970 ();
 sg13g2_fill_2 FILLER_93_977 ();
 sg13g2_fill_1 FILLER_93_979 ();
 sg13g2_decap_8 FILLER_93_988 ();
 sg13g2_decap_8 FILLER_93_995 ();
 sg13g2_decap_8 FILLER_93_1002 ();
 sg13g2_decap_8 FILLER_93_1009 ();
 sg13g2_decap_8 FILLER_93_1016 ();
 sg13g2_decap_8 FILLER_93_1023 ();
 sg13g2_decap_8 FILLER_93_1030 ();
 sg13g2_decap_8 FILLER_93_1037 ();
 sg13g2_decap_4 FILLER_93_1044 ();
 sg13g2_fill_1 FILLER_93_1048 ();
 sg13g2_decap_8 FILLER_93_1053 ();
 sg13g2_fill_2 FILLER_93_1060 ();
 sg13g2_decap_8 FILLER_93_1079 ();
 sg13g2_decap_8 FILLER_93_1086 ();
 sg13g2_decap_8 FILLER_93_1093 ();
 sg13g2_fill_1 FILLER_93_1100 ();
 sg13g2_decap_8 FILLER_93_1112 ();
 sg13g2_decap_8 FILLER_93_1119 ();
 sg13g2_decap_8 FILLER_93_1126 ();
 sg13g2_decap_8 FILLER_93_1133 ();
 sg13g2_decap_8 FILLER_93_1140 ();
 sg13g2_decap_8 FILLER_93_1147 ();
 sg13g2_decap_8 FILLER_93_1154 ();
 sg13g2_fill_2 FILLER_93_1161 ();
 sg13g2_fill_1 FILLER_93_1163 ();
 sg13g2_fill_1 FILLER_93_1172 ();
 sg13g2_decap_8 FILLER_93_1186 ();
 sg13g2_decap_8 FILLER_93_1193 ();
 sg13g2_decap_4 FILLER_93_1200 ();
 sg13g2_fill_2 FILLER_93_1204 ();
 sg13g2_decap_8 FILLER_93_1242 ();
 sg13g2_fill_2 FILLER_93_1249 ();
 sg13g2_fill_1 FILLER_93_1251 ();
 sg13g2_decap_4 FILLER_93_1287 ();
 sg13g2_fill_2 FILLER_93_1291 ();
 sg13g2_decap_4 FILLER_93_1314 ();
 sg13g2_fill_2 FILLER_93_1323 ();
 sg13g2_decap_8 FILLER_93_1329 ();
 sg13g2_decap_8 FILLER_93_1336 ();
 sg13g2_decap_8 FILLER_93_1343 ();
 sg13g2_decap_8 FILLER_93_1350 ();
 sg13g2_decap_8 FILLER_93_1357 ();
 sg13g2_decap_8 FILLER_93_1364 ();
 sg13g2_decap_8 FILLER_93_1374 ();
 sg13g2_decap_8 FILLER_93_1381 ();
 sg13g2_decap_8 FILLER_93_1388 ();
 sg13g2_decap_8 FILLER_93_1395 ();
 sg13g2_decap_8 FILLER_93_1402 ();
 sg13g2_fill_2 FILLER_93_1409 ();
 sg13g2_decap_8 FILLER_93_1424 ();
 sg13g2_decap_8 FILLER_93_1431 ();
 sg13g2_decap_8 FILLER_93_1438 ();
 sg13g2_decap_8 FILLER_93_1445 ();
 sg13g2_decap_8 FILLER_93_1452 ();
 sg13g2_decap_8 FILLER_93_1459 ();
 sg13g2_fill_1 FILLER_93_1466 ();
 sg13g2_decap_8 FILLER_93_1471 ();
 sg13g2_fill_2 FILLER_93_1490 ();
 sg13g2_decap_8 FILLER_93_1500 ();
 sg13g2_fill_1 FILLER_93_1507 ();
 sg13g2_fill_2 FILLER_93_1516 ();
 sg13g2_fill_1 FILLER_93_1518 ();
 sg13g2_decap_8 FILLER_93_1523 ();
 sg13g2_decap_8 FILLER_93_1530 ();
 sg13g2_decap_8 FILLER_93_1537 ();
 sg13g2_decap_8 FILLER_93_1544 ();
 sg13g2_fill_2 FILLER_93_1551 ();
 sg13g2_fill_1 FILLER_93_1553 ();
 sg13g2_decap_8 FILLER_93_1557 ();
 sg13g2_decap_8 FILLER_93_1564 ();
 sg13g2_decap_8 FILLER_93_1571 ();
 sg13g2_decap_8 FILLER_93_1578 ();
 sg13g2_decap_8 FILLER_93_1585 ();
 sg13g2_fill_2 FILLER_93_1592 ();
 sg13g2_fill_1 FILLER_93_1594 ();
 sg13g2_fill_2 FILLER_93_1603 ();
 sg13g2_fill_2 FILLER_93_1608 ();
 sg13g2_decap_4 FILLER_93_1626 ();
 sg13g2_fill_2 FILLER_93_1630 ();
 sg13g2_decap_8 FILLER_93_1648 ();
 sg13g2_decap_8 FILLER_93_1655 ();
 sg13g2_decap_8 FILLER_93_1662 ();
 sg13g2_decap_8 FILLER_93_1669 ();
 sg13g2_decap_4 FILLER_93_1676 ();
 sg13g2_fill_1 FILLER_93_1680 ();
 sg13g2_fill_2 FILLER_93_1689 ();
 sg13g2_decap_8 FILLER_93_1702 ();
 sg13g2_decap_8 FILLER_93_1709 ();
 sg13g2_decap_8 FILLER_93_1716 ();
 sg13g2_decap_8 FILLER_93_1723 ();
 sg13g2_decap_4 FILLER_93_1730 ();
 sg13g2_fill_1 FILLER_93_1734 ();
 sg13g2_decap_8 FILLER_93_1748 ();
 sg13g2_decap_8 FILLER_93_1755 ();
 sg13g2_decap_4 FILLER_93_1762 ();
 sg13g2_fill_2 FILLER_93_1766 ();
 sg13g2_decap_8 FILLER_94_0 ();
 sg13g2_decap_8 FILLER_94_7 ();
 sg13g2_decap_8 FILLER_94_14 ();
 sg13g2_fill_2 FILLER_94_21 ();
 sg13g2_fill_1 FILLER_94_23 ();
 sg13g2_fill_2 FILLER_94_37 ();
 sg13g2_fill_1 FILLER_94_39 ();
 sg13g2_decap_8 FILLER_94_48 ();
 sg13g2_decap_8 FILLER_94_55 ();
 sg13g2_decap_8 FILLER_94_62 ();
 sg13g2_decap_4 FILLER_94_73 ();
 sg13g2_decap_8 FILLER_94_98 ();
 sg13g2_decap_8 FILLER_94_105 ();
 sg13g2_decap_8 FILLER_94_112 ();
 sg13g2_decap_8 FILLER_94_119 ();
 sg13g2_decap_8 FILLER_94_126 ();
 sg13g2_decap_8 FILLER_94_133 ();
 sg13g2_decap_8 FILLER_94_140 ();
 sg13g2_fill_2 FILLER_94_147 ();
 sg13g2_decap_8 FILLER_94_154 ();
 sg13g2_decap_8 FILLER_94_161 ();
 sg13g2_decap_8 FILLER_94_168 ();
 sg13g2_decap_8 FILLER_94_191 ();
 sg13g2_decap_8 FILLER_94_198 ();
 sg13g2_decap_8 FILLER_94_205 ();
 sg13g2_decap_8 FILLER_94_212 ();
 sg13g2_decap_4 FILLER_94_219 ();
 sg13g2_fill_2 FILLER_94_223 ();
 sg13g2_decap_8 FILLER_94_236 ();
 sg13g2_decap_8 FILLER_94_243 ();
 sg13g2_fill_2 FILLER_94_267 ();
 sg13g2_fill_1 FILLER_94_269 ();
 sg13g2_decap_8 FILLER_94_278 ();
 sg13g2_decap_8 FILLER_94_285 ();
 sg13g2_decap_8 FILLER_94_292 ();
 sg13g2_decap_8 FILLER_94_299 ();
 sg13g2_decap_8 FILLER_94_306 ();
 sg13g2_decap_4 FILLER_94_313 ();
 sg13g2_fill_2 FILLER_94_317 ();
 sg13g2_decap_8 FILLER_94_327 ();
 sg13g2_decap_8 FILLER_94_334 ();
 sg13g2_decap_8 FILLER_94_341 ();
 sg13g2_decap_8 FILLER_94_348 ();
 sg13g2_decap_8 FILLER_94_355 ();
 sg13g2_decap_4 FILLER_94_362 ();
 sg13g2_decap_8 FILLER_94_379 ();
 sg13g2_decap_8 FILLER_94_395 ();
 sg13g2_decap_8 FILLER_94_402 ();
 sg13g2_decap_8 FILLER_94_409 ();
 sg13g2_decap_8 FILLER_94_416 ();
 sg13g2_fill_1 FILLER_94_423 ();
 sg13g2_decap_8 FILLER_94_432 ();
 sg13g2_decap_8 FILLER_94_439 ();
 sg13g2_decap_8 FILLER_94_446 ();
 sg13g2_decap_8 FILLER_94_453 ();
 sg13g2_decap_8 FILLER_94_460 ();
 sg13g2_decap_8 FILLER_94_467 ();
 sg13g2_fill_2 FILLER_94_474 ();
 sg13g2_fill_1 FILLER_94_476 ();
 sg13g2_decap_8 FILLER_94_489 ();
 sg13g2_decap_8 FILLER_94_496 ();
 sg13g2_decap_8 FILLER_94_503 ();
 sg13g2_decap_8 FILLER_94_510 ();
 sg13g2_decap_8 FILLER_94_517 ();
 sg13g2_decap_8 FILLER_94_524 ();
 sg13g2_decap_8 FILLER_94_531 ();
 sg13g2_fill_2 FILLER_94_538 ();
 sg13g2_decap_8 FILLER_94_552 ();
 sg13g2_decap_8 FILLER_94_559 ();
 sg13g2_decap_8 FILLER_94_566 ();
 sg13g2_decap_8 FILLER_94_573 ();
 sg13g2_decap_8 FILLER_94_580 ();
 sg13g2_decap_8 FILLER_94_587 ();
 sg13g2_decap_8 FILLER_94_594 ();
 sg13g2_decap_8 FILLER_94_601 ();
 sg13g2_decap_4 FILLER_94_608 ();
 sg13g2_decap_8 FILLER_94_625 ();
 sg13g2_decap_8 FILLER_94_632 ();
 sg13g2_decap_8 FILLER_94_639 ();
 sg13g2_decap_8 FILLER_94_646 ();
 sg13g2_fill_2 FILLER_94_653 ();
 sg13g2_decap_8 FILLER_94_669 ();
 sg13g2_decap_4 FILLER_94_676 ();
 sg13g2_fill_2 FILLER_94_680 ();
 sg13g2_decap_8 FILLER_94_691 ();
 sg13g2_decap_8 FILLER_94_698 ();
 sg13g2_decap_8 FILLER_94_705 ();
 sg13g2_decap_8 FILLER_94_712 ();
 sg13g2_decap_8 FILLER_94_719 ();
 sg13g2_decap_8 FILLER_94_726 ();
 sg13g2_decap_8 FILLER_94_733 ();
 sg13g2_decap_8 FILLER_94_740 ();
 sg13g2_decap_8 FILLER_94_747 ();
 sg13g2_fill_1 FILLER_94_754 ();
 sg13g2_decap_8 FILLER_94_763 ();
 sg13g2_fill_2 FILLER_94_770 ();
 sg13g2_fill_2 FILLER_94_785 ();
 sg13g2_decap_8 FILLER_94_795 ();
 sg13g2_decap_8 FILLER_94_802 ();
 sg13g2_decap_8 FILLER_94_809 ();
 sg13g2_decap_4 FILLER_94_816 ();
 sg13g2_fill_2 FILLER_94_820 ();
 sg13g2_decap_8 FILLER_94_841 ();
 sg13g2_decap_8 FILLER_94_848 ();
 sg13g2_decap_8 FILLER_94_855 ();
 sg13g2_decap_8 FILLER_94_862 ();
 sg13g2_decap_8 FILLER_94_882 ();
 sg13g2_decap_8 FILLER_94_889 ();
 sg13g2_decap_8 FILLER_94_896 ();
 sg13g2_decap_8 FILLER_94_903 ();
 sg13g2_decap_8 FILLER_94_910 ();
 sg13g2_fill_1 FILLER_94_917 ();
 sg13g2_decap_8 FILLER_94_931 ();
 sg13g2_decap_8 FILLER_94_938 ();
 sg13g2_decap_4 FILLER_94_945 ();
 sg13g2_fill_1 FILLER_94_949 ();
 sg13g2_decap_8 FILLER_94_976 ();
 sg13g2_decap_8 FILLER_94_983 ();
 sg13g2_decap_8 FILLER_94_990 ();
 sg13g2_decap_8 FILLER_94_997 ();
 sg13g2_fill_2 FILLER_94_1004 ();
 sg13g2_decap_4 FILLER_94_1019 ();
 sg13g2_fill_2 FILLER_94_1023 ();
 sg13g2_decap_8 FILLER_94_1064 ();
 sg13g2_decap_8 FILLER_94_1071 ();
 sg13g2_decap_8 FILLER_94_1078 ();
 sg13g2_decap_4 FILLER_94_1085 ();
 sg13g2_fill_1 FILLER_94_1089 ();
 sg13g2_decap_8 FILLER_94_1095 ();
 sg13g2_decap_8 FILLER_94_1102 ();
 sg13g2_fill_1 FILLER_94_1109 ();
 sg13g2_fill_2 FILLER_94_1115 ();
 sg13g2_decap_8 FILLER_94_1121 ();
 sg13g2_decap_8 FILLER_94_1128 ();
 sg13g2_decap_4 FILLER_94_1135 ();
 sg13g2_decap_8 FILLER_94_1155 ();
 sg13g2_decap_4 FILLER_94_1162 ();
 sg13g2_fill_2 FILLER_94_1174 ();
 sg13g2_decap_8 FILLER_94_1183 ();
 sg13g2_decap_8 FILLER_94_1190 ();
 sg13g2_decap_8 FILLER_94_1197 ();
 sg13g2_decap_4 FILLER_94_1204 ();
 sg13g2_decap_8 FILLER_94_1218 ();
 sg13g2_fill_2 FILLER_94_1225 ();
 sg13g2_decap_8 FILLER_94_1235 ();
 sg13g2_decap_8 FILLER_94_1242 ();
 sg13g2_decap_8 FILLER_94_1249 ();
 sg13g2_decap_8 FILLER_94_1256 ();
 sg13g2_decap_8 FILLER_94_1263 ();
 sg13g2_decap_4 FILLER_94_1270 ();
 sg13g2_fill_2 FILLER_94_1274 ();
 sg13g2_decap_8 FILLER_94_1289 ();
 sg13g2_decap_8 FILLER_94_1296 ();
 sg13g2_decap_8 FILLER_94_1303 ();
 sg13g2_decap_4 FILLER_94_1310 ();
 sg13g2_decap_4 FILLER_94_1319 ();
 sg13g2_decap_8 FILLER_94_1327 ();
 sg13g2_decap_8 FILLER_94_1334 ();
 sg13g2_decap_8 FILLER_94_1341 ();
 sg13g2_decap_8 FILLER_94_1348 ();
 sg13g2_decap_8 FILLER_94_1355 ();
 sg13g2_decap_8 FILLER_94_1362 ();
 sg13g2_decap_8 FILLER_94_1369 ();
 sg13g2_decap_8 FILLER_94_1376 ();
 sg13g2_decap_8 FILLER_94_1383 ();
 sg13g2_decap_8 FILLER_94_1390 ();
 sg13g2_decap_8 FILLER_94_1397 ();
 sg13g2_decap_8 FILLER_94_1404 ();
 sg13g2_decap_8 FILLER_94_1411 ();
 sg13g2_decap_8 FILLER_94_1418 ();
 sg13g2_decap_8 FILLER_94_1425 ();
 sg13g2_decap_8 FILLER_94_1432 ();
 sg13g2_fill_2 FILLER_94_1439 ();
 sg13g2_decap_8 FILLER_94_1467 ();
 sg13g2_decap_8 FILLER_94_1474 ();
 sg13g2_decap_8 FILLER_94_1481 ();
 sg13g2_decap_8 FILLER_94_1488 ();
 sg13g2_decap_8 FILLER_94_1495 ();
 sg13g2_decap_8 FILLER_94_1502 ();
 sg13g2_fill_2 FILLER_94_1509 ();
 sg13g2_decap_8 FILLER_94_1515 ();
 sg13g2_fill_1 FILLER_94_1522 ();
 sg13g2_decap_8 FILLER_94_1531 ();
 sg13g2_decap_8 FILLER_94_1538 ();
 sg13g2_decap_8 FILLER_94_1545 ();
 sg13g2_decap_8 FILLER_94_1556 ();
 sg13g2_decap_8 FILLER_94_1563 ();
 sg13g2_decap_8 FILLER_94_1570 ();
 sg13g2_decap_8 FILLER_94_1577 ();
 sg13g2_decap_8 FILLER_94_1584 ();
 sg13g2_decap_8 FILLER_94_1591 ();
 sg13g2_decap_8 FILLER_94_1598 ();
 sg13g2_fill_2 FILLER_94_1608 ();
 sg13g2_decap_8 FILLER_94_1613 ();
 sg13g2_decap_8 FILLER_94_1620 ();
 sg13g2_decap_8 FILLER_94_1627 ();
 sg13g2_fill_2 FILLER_94_1634 ();
 sg13g2_fill_1 FILLER_94_1636 ();
 sg13g2_decap_4 FILLER_94_1641 ();
 sg13g2_fill_1 FILLER_94_1645 ();
 sg13g2_decap_8 FILLER_94_1654 ();
 sg13g2_decap_8 FILLER_94_1661 ();
 sg13g2_decap_4 FILLER_94_1668 ();
 sg13g2_decap_8 FILLER_94_1680 ();
 sg13g2_fill_1 FILLER_94_1687 ();
 sg13g2_fill_2 FILLER_94_1699 ();
 sg13g2_decap_8 FILLER_94_1705 ();
 sg13g2_decap_8 FILLER_94_1712 ();
 sg13g2_decap_8 FILLER_94_1719 ();
 sg13g2_decap_4 FILLER_94_1726 ();
 sg13g2_decap_8 FILLER_94_1756 ();
 sg13g2_decap_4 FILLER_94_1763 ();
 sg13g2_fill_1 FILLER_94_1767 ();
 sg13g2_decap_8 FILLER_95_0 ();
 sg13g2_decap_8 FILLER_95_7 ();
 sg13g2_decap_8 FILLER_95_14 ();
 sg13g2_decap_8 FILLER_95_21 ();
 sg13g2_fill_2 FILLER_95_28 ();
 sg13g2_fill_2 FILLER_95_46 ();
 sg13g2_decap_8 FILLER_95_52 ();
 sg13g2_decap_8 FILLER_95_59 ();
 sg13g2_decap_8 FILLER_95_66 ();
 sg13g2_decap_8 FILLER_95_73 ();
 sg13g2_decap_4 FILLER_95_80 ();
 sg13g2_decap_8 FILLER_95_100 ();
 sg13g2_decap_8 FILLER_95_107 ();
 sg13g2_fill_2 FILLER_95_114 ();
 sg13g2_decap_8 FILLER_95_120 ();
 sg13g2_decap_4 FILLER_95_127 ();
 sg13g2_decap_8 FILLER_95_139 ();
 sg13g2_decap_8 FILLER_95_146 ();
 sg13g2_decap_8 FILLER_95_153 ();
 sg13g2_decap_8 FILLER_95_160 ();
 sg13g2_decap_8 FILLER_95_167 ();
 sg13g2_decap_4 FILLER_95_174 ();
 sg13g2_fill_2 FILLER_95_178 ();
 sg13g2_decap_8 FILLER_95_192 ();
 sg13g2_decap_8 FILLER_95_199 ();
 sg13g2_decap_8 FILLER_95_206 ();
 sg13g2_decap_8 FILLER_95_213 ();
 sg13g2_decap_8 FILLER_95_220 ();
 sg13g2_decap_8 FILLER_95_227 ();
 sg13g2_decap_8 FILLER_95_234 ();
 sg13g2_decap_8 FILLER_95_241 ();
 sg13g2_fill_2 FILLER_95_248 ();
 sg13g2_fill_1 FILLER_95_250 ();
 sg13g2_decap_8 FILLER_95_263 ();
 sg13g2_decap_8 FILLER_95_270 ();
 sg13g2_decap_8 FILLER_95_277 ();
 sg13g2_decap_8 FILLER_95_284 ();
 sg13g2_decap_4 FILLER_95_307 ();
 sg13g2_decap_8 FILLER_95_316 ();
 sg13g2_decap_8 FILLER_95_323 ();
 sg13g2_decap_8 FILLER_95_330 ();
 sg13g2_fill_2 FILLER_95_337 ();
 sg13g2_fill_1 FILLER_95_339 ();
 sg13g2_decap_8 FILLER_95_362 ();
 sg13g2_decap_8 FILLER_95_369 ();
 sg13g2_decap_8 FILLER_95_376 ();
 sg13g2_decap_8 FILLER_95_383 ();
 sg13g2_decap_8 FILLER_95_390 ();
 sg13g2_decap_8 FILLER_95_397 ();
 sg13g2_decap_8 FILLER_95_404 ();
 sg13g2_decap_8 FILLER_95_411 ();
 sg13g2_decap_4 FILLER_95_418 ();
 sg13g2_fill_2 FILLER_95_422 ();
 sg13g2_fill_2 FILLER_95_433 ();
 sg13g2_decap_8 FILLER_95_452 ();
 sg13g2_fill_1 FILLER_95_459 ();
 sg13g2_fill_2 FILLER_95_472 ();
 sg13g2_fill_1 FILLER_95_474 ();
 sg13g2_decap_8 FILLER_95_495 ();
 sg13g2_decap_8 FILLER_95_502 ();
 sg13g2_decap_8 FILLER_95_509 ();
 sg13g2_decap_4 FILLER_95_516 ();
 sg13g2_decap_4 FILLER_95_525 ();
 sg13g2_fill_2 FILLER_95_529 ();
 sg13g2_decap_8 FILLER_95_539 ();
 sg13g2_decap_8 FILLER_95_546 ();
 sg13g2_fill_2 FILLER_95_553 ();
 sg13g2_fill_1 FILLER_95_555 ();
 sg13g2_decap_8 FILLER_95_564 ();
 sg13g2_decap_8 FILLER_95_571 ();
 sg13g2_decap_8 FILLER_95_578 ();
 sg13g2_decap_8 FILLER_95_585 ();
 sg13g2_decap_8 FILLER_95_592 ();
 sg13g2_decap_4 FILLER_95_599 ();
 sg13g2_fill_2 FILLER_95_616 ();
 sg13g2_fill_1 FILLER_95_618 ();
 sg13g2_decap_8 FILLER_95_629 ();
 sg13g2_decap_8 FILLER_95_636 ();
 sg13g2_decap_8 FILLER_95_643 ();
 sg13g2_decap_8 FILLER_95_650 ();
 sg13g2_decap_8 FILLER_95_657 ();
 sg13g2_decap_8 FILLER_95_664 ();
 sg13g2_decap_8 FILLER_95_671 ();
 sg13g2_decap_8 FILLER_95_678 ();
 sg13g2_decap_8 FILLER_95_685 ();
 sg13g2_decap_8 FILLER_95_692 ();
 sg13g2_decap_8 FILLER_95_699 ();
 sg13g2_fill_2 FILLER_95_706 ();
 sg13g2_fill_1 FILLER_95_708 ();
 sg13g2_decap_8 FILLER_95_713 ();
 sg13g2_fill_2 FILLER_95_720 ();
 sg13g2_fill_1 FILLER_95_722 ();
 sg13g2_decap_8 FILLER_95_741 ();
 sg13g2_decap_8 FILLER_95_748 ();
 sg13g2_decap_8 FILLER_95_755 ();
 sg13g2_decap_8 FILLER_95_762 ();
 sg13g2_fill_1 FILLER_95_769 ();
 sg13g2_decap_8 FILLER_95_783 ();
 sg13g2_decap_8 FILLER_95_790 ();
 sg13g2_decap_8 FILLER_95_797 ();
 sg13g2_decap_8 FILLER_95_804 ();
 sg13g2_decap_8 FILLER_95_811 ();
 sg13g2_decap_8 FILLER_95_818 ();
 sg13g2_fill_2 FILLER_95_825 ();
 sg13g2_fill_2 FILLER_95_836 ();
 sg13g2_fill_1 FILLER_95_838 ();
 sg13g2_decap_8 FILLER_95_852 ();
 sg13g2_decap_8 FILLER_95_859 ();
 sg13g2_decap_8 FILLER_95_866 ();
 sg13g2_fill_1 FILLER_95_889 ();
 sg13g2_decap_8 FILLER_95_903 ();
 sg13g2_decap_8 FILLER_95_910 ();
 sg13g2_decap_8 FILLER_95_917 ();
 sg13g2_decap_8 FILLER_95_924 ();
 sg13g2_decap_8 FILLER_95_931 ();
 sg13g2_decap_8 FILLER_95_938 ();
 sg13g2_decap_8 FILLER_95_951 ();
 sg13g2_fill_2 FILLER_95_958 ();
 sg13g2_fill_1 FILLER_95_960 ();
 sg13g2_decap_8 FILLER_95_965 ();
 sg13g2_fill_1 FILLER_95_972 ();
 sg13g2_decap_8 FILLER_95_986 ();
 sg13g2_decap_8 FILLER_95_993 ();
 sg13g2_decap_8 FILLER_95_1000 ();
 sg13g2_decap_4 FILLER_95_1007 ();
 sg13g2_fill_1 FILLER_95_1011 ();
 sg13g2_decap_8 FILLER_95_1042 ();
 sg13g2_decap_8 FILLER_95_1049 ();
 sg13g2_decap_8 FILLER_95_1056 ();
 sg13g2_decap_8 FILLER_95_1063 ();
 sg13g2_decap_8 FILLER_95_1070 ();
 sg13g2_fill_2 FILLER_95_1077 ();
 sg13g2_fill_1 FILLER_95_1079 ();
 sg13g2_decap_8 FILLER_95_1153 ();
 sg13g2_decap_8 FILLER_95_1160 ();
 sg13g2_decap_8 FILLER_95_1167 ();
 sg13g2_decap_8 FILLER_95_1174 ();
 sg13g2_decap_8 FILLER_95_1181 ();
 sg13g2_decap_8 FILLER_95_1188 ();
 sg13g2_fill_2 FILLER_95_1195 ();
 sg13g2_decap_8 FILLER_95_1201 ();
 sg13g2_decap_8 FILLER_95_1208 ();
 sg13g2_decap_8 FILLER_95_1215 ();
 sg13g2_decap_8 FILLER_95_1222 ();
 sg13g2_decap_8 FILLER_95_1229 ();
 sg13g2_decap_8 FILLER_95_1236 ();
 sg13g2_decap_8 FILLER_95_1243 ();
 sg13g2_fill_1 FILLER_95_1250 ();
 sg13g2_decap_8 FILLER_95_1260 ();
 sg13g2_decap_8 FILLER_95_1267 ();
 sg13g2_decap_8 FILLER_95_1274 ();
 sg13g2_decap_8 FILLER_95_1281 ();
 sg13g2_decap_8 FILLER_95_1288 ();
 sg13g2_decap_8 FILLER_95_1295 ();
 sg13g2_decap_8 FILLER_95_1302 ();
 sg13g2_decap_8 FILLER_95_1309 ();
 sg13g2_decap_8 FILLER_95_1320 ();
 sg13g2_decap_4 FILLER_95_1327 ();
 sg13g2_fill_2 FILLER_95_1331 ();
 sg13g2_decap_8 FILLER_95_1341 ();
 sg13g2_decap_8 FILLER_95_1348 ();
 sg13g2_decap_8 FILLER_95_1355 ();
 sg13g2_fill_2 FILLER_95_1366 ();
 sg13g2_fill_1 FILLER_95_1368 ();
 sg13g2_fill_2 FILLER_95_1374 ();
 sg13g2_decap_4 FILLER_95_1402 ();
 sg13g2_fill_2 FILLER_95_1406 ();
 sg13g2_decap_8 FILLER_95_1414 ();
 sg13g2_decap_8 FILLER_95_1421 ();
 sg13g2_decap_8 FILLER_95_1428 ();
 sg13g2_fill_1 FILLER_95_1435 ();
 sg13g2_fill_2 FILLER_95_1444 ();
 sg13g2_fill_1 FILLER_95_1446 ();
 sg13g2_decap_8 FILLER_95_1465 ();
 sg13g2_decap_8 FILLER_95_1472 ();
 sg13g2_decap_8 FILLER_95_1479 ();
 sg13g2_decap_8 FILLER_95_1486 ();
 sg13g2_decap_8 FILLER_95_1505 ();
 sg13g2_decap_8 FILLER_95_1512 ();
 sg13g2_decap_8 FILLER_95_1519 ();
 sg13g2_decap_8 FILLER_95_1526 ();
 sg13g2_decap_8 FILLER_95_1533 ();
 sg13g2_decap_4 FILLER_95_1540 ();
 sg13g2_fill_1 FILLER_95_1544 ();
 sg13g2_decap_8 FILLER_95_1566 ();
 sg13g2_decap_8 FILLER_95_1573 ();
 sg13g2_decap_8 FILLER_95_1580 ();
 sg13g2_decap_4 FILLER_95_1587 ();
 sg13g2_decap_4 FILLER_95_1599 ();
 sg13g2_fill_2 FILLER_95_1616 ();
 sg13g2_fill_1 FILLER_95_1618 ();
 sg13g2_decap_8 FILLER_95_1632 ();
 sg13g2_decap_8 FILLER_95_1639 ();
 sg13g2_decap_8 FILLER_95_1646 ();
 sg13g2_decap_8 FILLER_95_1653 ();
 sg13g2_decap_8 FILLER_95_1660 ();
 sg13g2_decap_8 FILLER_95_1667 ();
 sg13g2_decap_8 FILLER_95_1674 ();
 sg13g2_fill_2 FILLER_95_1681 ();
 sg13g2_decap_8 FILLER_95_1713 ();
 sg13g2_decap_8 FILLER_95_1720 ();
 sg13g2_decap_8 FILLER_95_1727 ();
 sg13g2_decap_8 FILLER_95_1734 ();
 sg13g2_fill_1 FILLER_95_1745 ();
 sg13g2_decap_8 FILLER_95_1759 ();
 sg13g2_fill_2 FILLER_95_1766 ();
 sg13g2_decap_8 FILLER_96_0 ();
 sg13g2_decap_8 FILLER_96_7 ();
 sg13g2_decap_4 FILLER_96_14 ();
 sg13g2_decap_8 FILLER_96_39 ();
 sg13g2_decap_8 FILLER_96_46 ();
 sg13g2_decap_4 FILLER_96_53 ();
 sg13g2_fill_2 FILLER_96_57 ();
 sg13g2_decap_8 FILLER_96_68 ();
 sg13g2_decap_8 FILLER_96_75 ();
 sg13g2_decap_8 FILLER_96_82 ();
 sg13g2_decap_8 FILLER_96_89 ();
 sg13g2_decap_4 FILLER_96_96 ();
 sg13g2_fill_2 FILLER_96_121 ();
 sg13g2_fill_1 FILLER_96_123 ();
 sg13g2_decap_8 FILLER_96_129 ();
 sg13g2_decap_8 FILLER_96_136 ();
 sg13g2_decap_8 FILLER_96_143 ();
 sg13g2_decap_8 FILLER_96_150 ();
 sg13g2_decap_8 FILLER_96_157 ();
 sg13g2_decap_4 FILLER_96_164 ();
 sg13g2_fill_2 FILLER_96_171 ();
 sg13g2_fill_1 FILLER_96_173 ();
 sg13g2_decap_8 FILLER_96_182 ();
 sg13g2_decap_8 FILLER_96_189 ();
 sg13g2_decap_4 FILLER_96_196 ();
 sg13g2_fill_1 FILLER_96_200 ();
 sg13g2_decap_8 FILLER_96_207 ();
 sg13g2_decap_8 FILLER_96_214 ();
 sg13g2_decap_8 FILLER_96_221 ();
 sg13g2_decap_8 FILLER_96_228 ();
 sg13g2_decap_8 FILLER_96_235 ();
 sg13g2_decap_8 FILLER_96_242 ();
 sg13g2_decap_8 FILLER_96_249 ();
 sg13g2_decap_8 FILLER_96_256 ();
 sg13g2_decap_8 FILLER_96_263 ();
 sg13g2_decap_8 FILLER_96_270 ();
 sg13g2_decap_8 FILLER_96_277 ();
 sg13g2_fill_1 FILLER_96_284 ();
 sg13g2_decap_4 FILLER_96_290 ();
 sg13g2_decap_8 FILLER_96_302 ();
 sg13g2_decap_8 FILLER_96_309 ();
 sg13g2_decap_8 FILLER_96_316 ();
 sg13g2_fill_1 FILLER_96_323 ();
 sg13g2_decap_8 FILLER_96_342 ();
 sg13g2_decap_8 FILLER_96_349 ();
 sg13g2_decap_8 FILLER_96_356 ();
 sg13g2_decap_8 FILLER_96_363 ();
 sg13g2_decap_8 FILLER_96_370 ();
 sg13g2_decap_8 FILLER_96_377 ();
 sg13g2_fill_2 FILLER_96_384 ();
 sg13g2_fill_1 FILLER_96_386 ();
 sg13g2_decap_8 FILLER_96_399 ();
 sg13g2_decap_8 FILLER_96_406 ();
 sg13g2_decap_8 FILLER_96_413 ();
 sg13g2_decap_8 FILLER_96_420 ();
 sg13g2_decap_8 FILLER_96_427 ();
 sg13g2_decap_8 FILLER_96_434 ();
 sg13g2_decap_8 FILLER_96_441 ();
 sg13g2_decap_8 FILLER_96_448 ();
 sg13g2_fill_2 FILLER_96_459 ();
 sg13g2_fill_1 FILLER_96_461 ();
 sg13g2_decap_8 FILLER_96_492 ();
 sg13g2_decap_8 FILLER_96_499 ();
 sg13g2_decap_8 FILLER_96_506 ();
 sg13g2_fill_2 FILLER_96_513 ();
 sg13g2_fill_2 FILLER_96_523 ();
 sg13g2_fill_1 FILLER_96_525 ();
 sg13g2_decap_8 FILLER_96_532 ();
 sg13g2_decap_8 FILLER_96_539 ();
 sg13g2_fill_2 FILLER_96_546 ();
 sg13g2_fill_1 FILLER_96_548 ();
 sg13g2_decap_4 FILLER_96_555 ();
 sg13g2_decap_8 FILLER_96_574 ();
 sg13g2_decap_8 FILLER_96_581 ();
 sg13g2_fill_1 FILLER_96_588 ();
 sg13g2_decap_8 FILLER_96_598 ();
 sg13g2_fill_2 FILLER_96_605 ();
 sg13g2_fill_1 FILLER_96_607 ();
 sg13g2_decap_8 FILLER_96_621 ();
 sg13g2_decap_8 FILLER_96_628 ();
 sg13g2_decap_8 FILLER_96_635 ();
 sg13g2_fill_2 FILLER_96_642 ();
 sg13g2_decap_4 FILLER_96_660 ();
 sg13g2_fill_2 FILLER_96_664 ();
 sg13g2_decap_8 FILLER_96_674 ();
 sg13g2_decap_8 FILLER_96_681 ();
 sg13g2_fill_1 FILLER_96_688 ();
 sg13g2_decap_4 FILLER_96_724 ();
 sg13g2_fill_1 FILLER_96_728 ();
 sg13g2_fill_2 FILLER_96_737 ();
 sg13g2_fill_1 FILLER_96_739 ();
 sg13g2_decap_8 FILLER_96_745 ();
 sg13g2_decap_8 FILLER_96_752 ();
 sg13g2_decap_8 FILLER_96_759 ();
 sg13g2_decap_8 FILLER_96_766 ();
 sg13g2_decap_8 FILLER_96_773 ();
 sg13g2_decap_8 FILLER_96_780 ();
 sg13g2_fill_2 FILLER_96_787 ();
 sg13g2_decap_8 FILLER_96_815 ();
 sg13g2_fill_1 FILLER_96_822 ();
 sg13g2_decap_8 FILLER_96_836 ();
 sg13g2_decap_8 FILLER_96_843 ();
 sg13g2_decap_8 FILLER_96_850 ();
 sg13g2_decap_8 FILLER_96_857 ();
 sg13g2_decap_8 FILLER_96_864 ();
 sg13g2_decap_8 FILLER_96_871 ();
 sg13g2_decap_4 FILLER_96_878 ();
 sg13g2_decap_4 FILLER_96_886 ();
 sg13g2_fill_2 FILLER_96_890 ();
 sg13g2_decap_8 FILLER_96_904 ();
 sg13g2_decap_8 FILLER_96_911 ();
 sg13g2_decap_8 FILLER_96_918 ();
 sg13g2_fill_2 FILLER_96_925 ();
 sg13g2_fill_1 FILLER_96_927 ();
 sg13g2_decap_8 FILLER_96_941 ();
 sg13g2_fill_1 FILLER_96_948 ();
 sg13g2_decap_4 FILLER_96_962 ();
 sg13g2_decap_8 FILLER_96_979 ();
 sg13g2_decap_8 FILLER_96_986 ();
 sg13g2_fill_2 FILLER_96_993 ();
 sg13g2_decap_8 FILLER_96_1000 ();
 sg13g2_decap_8 FILLER_96_1007 ();
 sg13g2_decap_8 FILLER_96_1014 ();
 sg13g2_decap_8 FILLER_96_1021 ();
 sg13g2_decap_8 FILLER_96_1032 ();
 sg13g2_decap_8 FILLER_96_1039 ();
 sg13g2_decap_8 FILLER_96_1046 ();
 sg13g2_decap_8 FILLER_96_1053 ();
 sg13g2_fill_2 FILLER_96_1060 ();
 sg13g2_fill_1 FILLER_96_1062 ();
 sg13g2_decap_8 FILLER_96_1069 ();
 sg13g2_decap_8 FILLER_96_1076 ();
 sg13g2_decap_4 FILLER_96_1083 ();
 sg13g2_decap_4 FILLER_96_1109 ();
 sg13g2_decap_8 FILLER_96_1117 ();
 sg13g2_decap_8 FILLER_96_1124 ();
 sg13g2_fill_1 FILLER_96_1131 ();
 sg13g2_decap_8 FILLER_96_1141 ();
 sg13g2_decap_4 FILLER_96_1148 ();
 sg13g2_fill_1 FILLER_96_1152 ();
 sg13g2_decap_8 FILLER_96_1166 ();
 sg13g2_decap_8 FILLER_96_1173 ();
 sg13g2_decap_8 FILLER_96_1180 ();
 sg13g2_decap_8 FILLER_96_1187 ();
 sg13g2_decap_4 FILLER_96_1194 ();
 sg13g2_fill_2 FILLER_96_1198 ();
 sg13g2_decap_8 FILLER_96_1212 ();
 sg13g2_decap_8 FILLER_96_1219 ();
 sg13g2_decap_4 FILLER_96_1226 ();
 sg13g2_decap_4 FILLER_96_1233 ();
 sg13g2_fill_1 FILLER_96_1237 ();
 sg13g2_decap_8 FILLER_96_1247 ();
 sg13g2_decap_8 FILLER_96_1254 ();
 sg13g2_decap_8 FILLER_96_1261 ();
 sg13g2_decap_8 FILLER_96_1268 ();
 sg13g2_fill_2 FILLER_96_1275 ();
 sg13g2_decap_8 FILLER_96_1281 ();
 sg13g2_decap_8 FILLER_96_1288 ();
 sg13g2_decap_8 FILLER_96_1295 ();
 sg13g2_fill_2 FILLER_96_1302 ();
 sg13g2_decap_8 FILLER_96_1338 ();
 sg13g2_decap_4 FILLER_96_1345 ();
 sg13g2_fill_2 FILLER_96_1349 ();
 sg13g2_decap_4 FILLER_96_1355 ();
 sg13g2_fill_1 FILLER_96_1359 ();
 sg13g2_decap_8 FILLER_96_1391 ();
 sg13g2_decap_8 FILLER_96_1398 ();
 sg13g2_decap_8 FILLER_96_1405 ();
 sg13g2_decap_8 FILLER_96_1412 ();
 sg13g2_decap_8 FILLER_96_1419 ();
 sg13g2_decap_8 FILLER_96_1432 ();
 sg13g2_decap_4 FILLER_96_1439 ();
 sg13g2_fill_2 FILLER_96_1443 ();
 sg13g2_decap_8 FILLER_96_1449 ();
 sg13g2_decap_8 FILLER_96_1456 ();
 sg13g2_decap_8 FILLER_96_1463 ();
 sg13g2_decap_8 FILLER_96_1470 ();
 sg13g2_decap_8 FILLER_96_1477 ();
 sg13g2_decap_8 FILLER_96_1484 ();
 sg13g2_decap_8 FILLER_96_1491 ();
 sg13g2_decap_8 FILLER_96_1498 ();
 sg13g2_fill_1 FILLER_96_1505 ();
 sg13g2_fill_1 FILLER_96_1510 ();
 sg13g2_decap_8 FILLER_96_1519 ();
 sg13g2_fill_2 FILLER_96_1526 ();
 sg13g2_fill_1 FILLER_96_1528 ();
 sg13g2_decap_8 FILLER_96_1534 ();
 sg13g2_decap_8 FILLER_96_1541 ();
 sg13g2_decap_8 FILLER_96_1548 ();
 sg13g2_decap_4 FILLER_96_1555 ();
 sg13g2_decap_8 FILLER_96_1563 ();
 sg13g2_decap_8 FILLER_96_1570 ();
 sg13g2_decap_8 FILLER_96_1597 ();
 sg13g2_decap_8 FILLER_96_1604 ();
 sg13g2_fill_2 FILLER_96_1611 ();
 sg13g2_fill_1 FILLER_96_1613 ();
 sg13g2_fill_1 FILLER_96_1620 ();
 sg13g2_decap_8 FILLER_96_1634 ();
 sg13g2_decap_8 FILLER_96_1641 ();
 sg13g2_fill_2 FILLER_96_1648 ();
 sg13g2_decap_8 FILLER_96_1659 ();
 sg13g2_decap_8 FILLER_96_1666 ();
 sg13g2_decap_8 FILLER_96_1673 ();
 sg13g2_decap_8 FILLER_96_1698 ();
 sg13g2_decap_8 FILLER_96_1705 ();
 sg13g2_decap_8 FILLER_96_1712 ();
 sg13g2_decap_8 FILLER_96_1719 ();
 sg13g2_decap_8 FILLER_96_1726 ();
 sg13g2_decap_8 FILLER_96_1733 ();
 sg13g2_decap_8 FILLER_96_1740 ();
 sg13g2_decap_8 FILLER_96_1747 ();
 sg13g2_decap_8 FILLER_96_1754 ();
 sg13g2_decap_8 FILLER_96_1761 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_8 FILLER_97_7 ();
 sg13g2_decap_4 FILLER_97_14 ();
 sg13g2_fill_2 FILLER_97_22 ();
 sg13g2_fill_1 FILLER_97_31 ();
 sg13g2_fill_2 FILLER_97_40 ();
 sg13g2_decap_8 FILLER_97_48 ();
 sg13g2_decap_8 FILLER_97_55 ();
 sg13g2_decap_8 FILLER_97_62 ();
 sg13g2_decap_8 FILLER_97_69 ();
 sg13g2_decap_8 FILLER_97_76 ();
 sg13g2_decap_8 FILLER_97_83 ();
 sg13g2_decap_8 FILLER_97_90 ();
 sg13g2_decap_8 FILLER_97_97 ();
 sg13g2_decap_8 FILLER_97_104 ();
 sg13g2_fill_2 FILLER_97_111 ();
 sg13g2_fill_1 FILLER_97_113 ();
 sg13g2_fill_2 FILLER_97_118 ();
 sg13g2_decap_8 FILLER_97_138 ();
 sg13g2_decap_8 FILLER_97_145 ();
 sg13g2_decap_8 FILLER_97_152 ();
 sg13g2_decap_8 FILLER_97_159 ();
 sg13g2_decap_4 FILLER_97_166 ();
 sg13g2_fill_2 FILLER_97_170 ();
 sg13g2_decap_8 FILLER_97_184 ();
 sg13g2_decap_4 FILLER_97_191 ();
 sg13g2_decap_8 FILLER_97_203 ();
 sg13g2_decap_8 FILLER_97_210 ();
 sg13g2_decap_8 FILLER_97_217 ();
 sg13g2_decap_4 FILLER_97_224 ();
 sg13g2_fill_2 FILLER_97_233 ();
 sg13g2_decap_8 FILLER_97_245 ();
 sg13g2_decap_8 FILLER_97_252 ();
 sg13g2_fill_2 FILLER_97_259 ();
 sg13g2_fill_1 FILLER_97_261 ();
 sg13g2_decap_8 FILLER_97_270 ();
 sg13g2_decap_8 FILLER_97_277 ();
 sg13g2_fill_1 FILLER_97_284 ();
 sg13g2_decap_8 FILLER_97_290 ();
 sg13g2_decap_4 FILLER_97_297 ();
 sg13g2_fill_2 FILLER_97_301 ();
 sg13g2_decap_8 FILLER_97_324 ();
 sg13g2_decap_8 FILLER_97_331 ();
 sg13g2_decap_8 FILLER_97_338 ();
 sg13g2_decap_8 FILLER_97_345 ();
 sg13g2_decap_8 FILLER_97_352 ();
 sg13g2_decap_8 FILLER_97_359 ();
 sg13g2_decap_4 FILLER_97_366 ();
 sg13g2_decap_8 FILLER_97_374 ();
 sg13g2_decap_8 FILLER_97_381 ();
 sg13g2_decap_8 FILLER_97_388 ();
 sg13g2_decap_8 FILLER_97_395 ();
 sg13g2_decap_8 FILLER_97_402 ();
 sg13g2_decap_8 FILLER_97_409 ();
 sg13g2_decap_8 FILLER_97_416 ();
 sg13g2_decap_8 FILLER_97_423 ();
 sg13g2_decap_8 FILLER_97_430 ();
 sg13g2_decap_8 FILLER_97_437 ();
 sg13g2_decap_8 FILLER_97_444 ();
 sg13g2_decap_8 FILLER_97_451 ();
 sg13g2_decap_8 FILLER_97_458 ();
 sg13g2_fill_2 FILLER_97_465 ();
 sg13g2_fill_2 FILLER_97_476 ();
 sg13g2_fill_1 FILLER_97_483 ();
 sg13g2_decap_8 FILLER_97_492 ();
 sg13g2_decap_8 FILLER_97_499 ();
 sg13g2_decap_8 FILLER_97_506 ();
 sg13g2_decap_8 FILLER_97_513 ();
 sg13g2_decap_8 FILLER_97_520 ();
 sg13g2_decap_8 FILLER_97_535 ();
 sg13g2_fill_1 FILLER_97_542 ();
 sg13g2_fill_2 FILLER_97_553 ();
 sg13g2_decap_4 FILLER_97_563 ();
 sg13g2_fill_2 FILLER_97_567 ();
 sg13g2_fill_2 FILLER_97_616 ();
 sg13g2_fill_1 FILLER_97_618 ();
 sg13g2_decap_8 FILLER_97_666 ();
 sg13g2_decap_8 FILLER_97_673 ();
 sg13g2_decap_8 FILLER_97_680 ();
 sg13g2_decap_8 FILLER_97_687 ();
 sg13g2_decap_8 FILLER_97_694 ();
 sg13g2_decap_8 FILLER_97_701 ();
 sg13g2_decap_8 FILLER_97_708 ();
 sg13g2_decap_8 FILLER_97_715 ();
 sg13g2_decap_8 FILLER_97_722 ();
 sg13g2_decap_8 FILLER_97_729 ();
 sg13g2_decap_8 FILLER_97_736 ();
 sg13g2_decap_8 FILLER_97_743 ();
 sg13g2_decap_8 FILLER_97_750 ();
 sg13g2_decap_8 FILLER_97_757 ();
 sg13g2_decap_8 FILLER_97_764 ();
 sg13g2_decap_8 FILLER_97_779 ();
 sg13g2_decap_8 FILLER_97_786 ();
 sg13g2_decap_8 FILLER_97_793 ();
 sg13g2_decap_8 FILLER_97_804 ();
 sg13g2_decap_8 FILLER_97_811 ();
 sg13g2_fill_2 FILLER_97_818 ();
 sg13g2_fill_1 FILLER_97_820 ();
 sg13g2_decap_8 FILLER_97_829 ();
 sg13g2_decap_8 FILLER_97_836 ();
 sg13g2_decap_8 FILLER_97_843 ();
 sg13g2_decap_8 FILLER_97_850 ();
 sg13g2_decap_8 FILLER_97_857 ();
 sg13g2_decap_4 FILLER_97_864 ();
 sg13g2_fill_2 FILLER_97_868 ();
 sg13g2_decap_4 FILLER_97_892 ();
 sg13g2_decap_4 FILLER_97_904 ();
 sg13g2_fill_2 FILLER_97_908 ();
 sg13g2_fill_2 FILLER_97_923 ();
 sg13g2_fill_1 FILLER_97_925 ();
 sg13g2_decap_4 FILLER_97_932 ();
 sg13g2_fill_2 FILLER_97_936 ();
 sg13g2_decap_4 FILLER_97_964 ();
 sg13g2_fill_1 FILLER_97_968 ();
 sg13g2_decap_8 FILLER_97_974 ();
 sg13g2_decap_8 FILLER_97_981 ();
 sg13g2_decap_8 FILLER_97_988 ();
 sg13g2_decap_8 FILLER_97_995 ();
 sg13g2_decap_8 FILLER_97_1002 ();
 sg13g2_decap_8 FILLER_97_1009 ();
 sg13g2_fill_1 FILLER_97_1016 ();
 sg13g2_decap_8 FILLER_97_1022 ();
 sg13g2_decap_8 FILLER_97_1029 ();
 sg13g2_decap_8 FILLER_97_1036 ();
 sg13g2_decap_8 FILLER_97_1043 ();
 sg13g2_decap_8 FILLER_97_1050 ();
 sg13g2_decap_8 FILLER_97_1057 ();
 sg13g2_decap_8 FILLER_97_1064 ();
 sg13g2_decap_8 FILLER_97_1071 ();
 sg13g2_fill_1 FILLER_97_1078 ();
 sg13g2_decap_8 FILLER_97_1084 ();
 sg13g2_decap_8 FILLER_97_1103 ();
 sg13g2_decap_8 FILLER_97_1110 ();
 sg13g2_decap_8 FILLER_97_1117 ();
 sg13g2_decap_8 FILLER_97_1124 ();
 sg13g2_decap_8 FILLER_97_1131 ();
 sg13g2_decap_8 FILLER_97_1138 ();
 sg13g2_fill_1 FILLER_97_1145 ();
 sg13g2_decap_8 FILLER_97_1149 ();
 sg13g2_fill_2 FILLER_97_1164 ();
 sg13g2_fill_1 FILLER_97_1166 ();
 sg13g2_fill_2 FILLER_97_1170 ();
 sg13g2_decap_8 FILLER_97_1182 ();
 sg13g2_fill_2 FILLER_97_1189 ();
 sg13g2_fill_2 FILLER_97_1222 ();
 sg13g2_fill_1 FILLER_97_1224 ();
 sg13g2_decap_4 FILLER_97_1245 ();
 sg13g2_decap_4 FILLER_97_1262 ();
 sg13g2_decap_8 FILLER_97_1281 ();
 sg13g2_decap_8 FILLER_97_1288 ();
 sg13g2_decap_8 FILLER_97_1295 ();
 sg13g2_decap_8 FILLER_97_1302 ();
 sg13g2_fill_2 FILLER_97_1319 ();
 sg13g2_fill_1 FILLER_97_1321 ();
 sg13g2_decap_8 FILLER_97_1335 ();
 sg13g2_decap_8 FILLER_97_1342 ();
 sg13g2_decap_4 FILLER_97_1349 ();
 sg13g2_decap_8 FILLER_97_1358 ();
 sg13g2_decap_8 FILLER_97_1365 ();
 sg13g2_fill_2 FILLER_97_1372 ();
 sg13g2_fill_2 FILLER_97_1387 ();
 sg13g2_fill_1 FILLER_97_1389 ();
 sg13g2_fill_2 FILLER_97_1403 ();
 sg13g2_fill_1 FILLER_97_1405 ();
 sg13g2_decap_8 FILLER_97_1419 ();
 sg13g2_decap_8 FILLER_97_1426 ();
 sg13g2_decap_8 FILLER_97_1433 ();
 sg13g2_decap_4 FILLER_97_1440 ();
 sg13g2_fill_1 FILLER_97_1444 ();
 sg13g2_decap_8 FILLER_97_1458 ();
 sg13g2_decap_8 FILLER_97_1465 ();
 sg13g2_decap_8 FILLER_97_1472 ();
 sg13g2_decap_8 FILLER_97_1479 ();
 sg13g2_fill_2 FILLER_97_1486 ();
 sg13g2_fill_2 FILLER_97_1496 ();
 sg13g2_fill_1 FILLER_97_1498 ();
 sg13g2_decap_8 FILLER_97_1542 ();
 sg13g2_decap_8 FILLER_97_1549 ();
 sg13g2_decap_8 FILLER_97_1556 ();
 sg13g2_decap_8 FILLER_97_1563 ();
 sg13g2_decap_8 FILLER_97_1570 ();
 sg13g2_decap_8 FILLER_97_1577 ();
 sg13g2_decap_8 FILLER_97_1584 ();
 sg13g2_decap_8 FILLER_97_1591 ();
 sg13g2_decap_4 FILLER_97_1598 ();
 sg13g2_fill_2 FILLER_97_1602 ();
 sg13g2_decap_8 FILLER_97_1626 ();
 sg13g2_decap_8 FILLER_97_1633 ();
 sg13g2_decap_8 FILLER_97_1640 ();
 sg13g2_fill_2 FILLER_97_1647 ();
 sg13g2_fill_1 FILLER_97_1649 ();
 sg13g2_decap_8 FILLER_97_1663 ();
 sg13g2_decap_8 FILLER_97_1670 ();
 sg13g2_fill_1 FILLER_97_1677 ();
 sg13g2_decap_8 FILLER_97_1694 ();
 sg13g2_decap_8 FILLER_97_1701 ();
 sg13g2_decap_4 FILLER_97_1708 ();
 sg13g2_decap_8 FILLER_97_1721 ();
 sg13g2_decap_8 FILLER_97_1728 ();
 sg13g2_decap_8 FILLER_97_1735 ();
 sg13g2_decap_8 FILLER_97_1742 ();
 sg13g2_decap_8 FILLER_97_1749 ();
 sg13g2_decap_8 FILLER_97_1756 ();
 sg13g2_decap_4 FILLER_97_1763 ();
 sg13g2_fill_1 FILLER_97_1767 ();
 sg13g2_decap_8 FILLER_98_0 ();
 sg13g2_decap_8 FILLER_98_7 ();
 sg13g2_fill_1 FILLER_98_14 ();
 sg13g2_decap_8 FILLER_98_40 ();
 sg13g2_decap_8 FILLER_98_47 ();
 sg13g2_decap_8 FILLER_98_54 ();
 sg13g2_decap_4 FILLER_98_61 ();
 sg13g2_fill_1 FILLER_98_65 ();
 sg13g2_decap_8 FILLER_98_70 ();
 sg13g2_decap_8 FILLER_98_77 ();
 sg13g2_decap_8 FILLER_98_84 ();
 sg13g2_decap_8 FILLER_98_91 ();
 sg13g2_decap_8 FILLER_98_98 ();
 sg13g2_decap_8 FILLER_98_105 ();
 sg13g2_decap_8 FILLER_98_112 ();
 sg13g2_decap_8 FILLER_98_119 ();
 sg13g2_decap_8 FILLER_98_126 ();
 sg13g2_decap_8 FILLER_98_133 ();
 sg13g2_decap_8 FILLER_98_140 ();
 sg13g2_decap_8 FILLER_98_147 ();
 sg13g2_decap_8 FILLER_98_154 ();
 sg13g2_decap_8 FILLER_98_161 ();
 sg13g2_fill_2 FILLER_98_168 ();
 sg13g2_fill_1 FILLER_98_170 ();
 sg13g2_fill_1 FILLER_98_175 ();
 sg13g2_decap_8 FILLER_98_181 ();
 sg13g2_decap_8 FILLER_98_188 ();
 sg13g2_fill_2 FILLER_98_195 ();
 sg13g2_fill_1 FILLER_98_197 ();
 sg13g2_decap_4 FILLER_98_212 ();
 sg13g2_decap_8 FILLER_98_220 ();
 sg13g2_fill_2 FILLER_98_227 ();
 sg13g2_fill_1 FILLER_98_229 ();
 sg13g2_decap_8 FILLER_98_235 ();
 sg13g2_decap_8 FILLER_98_242 ();
 sg13g2_decap_8 FILLER_98_249 ();
 sg13g2_decap_8 FILLER_98_256 ();
 sg13g2_decap_8 FILLER_98_263 ();
 sg13g2_decap_8 FILLER_98_270 ();
 sg13g2_fill_1 FILLER_98_277 ();
 sg13g2_decap_8 FILLER_98_286 ();
 sg13g2_decap_8 FILLER_98_293 ();
 sg13g2_decap_8 FILLER_98_300 ();
 sg13g2_decap_8 FILLER_98_307 ();
 sg13g2_fill_2 FILLER_98_314 ();
 sg13g2_decap_8 FILLER_98_333 ();
 sg13g2_decap_8 FILLER_98_340 ();
 sg13g2_decap_8 FILLER_98_347 ();
 sg13g2_decap_8 FILLER_98_354 ();
 sg13g2_decap_8 FILLER_98_361 ();
 sg13g2_fill_2 FILLER_98_368 ();
 sg13g2_fill_1 FILLER_98_370 ();
 sg13g2_decap_4 FILLER_98_376 ();
 sg13g2_decap_8 FILLER_98_385 ();
 sg13g2_fill_2 FILLER_98_392 ();
 sg13g2_fill_1 FILLER_98_394 ();
 sg13g2_decap_4 FILLER_98_400 ();
 sg13g2_decap_8 FILLER_98_426 ();
 sg13g2_decap_8 FILLER_98_433 ();
 sg13g2_decap_8 FILLER_98_440 ();
 sg13g2_decap_8 FILLER_98_447 ();
 sg13g2_decap_8 FILLER_98_454 ();
 sg13g2_fill_2 FILLER_98_461 ();
 sg13g2_fill_1 FILLER_98_463 ();
 sg13g2_decap_8 FILLER_98_471 ();
 sg13g2_decap_8 FILLER_98_478 ();
 sg13g2_decap_8 FILLER_98_485 ();
 sg13g2_decap_8 FILLER_98_492 ();
 sg13g2_decap_8 FILLER_98_499 ();
 sg13g2_decap_8 FILLER_98_506 ();
 sg13g2_decap_8 FILLER_98_516 ();
 sg13g2_decap_8 FILLER_98_523 ();
 sg13g2_fill_2 FILLER_98_530 ();
 sg13g2_fill_1 FILLER_98_532 ();
 sg13g2_decap_8 FILLER_98_537 ();
 sg13g2_decap_4 FILLER_98_544 ();
 sg13g2_fill_1 FILLER_98_548 ();
 sg13g2_decap_8 FILLER_98_552 ();
 sg13g2_decap_8 FILLER_98_559 ();
 sg13g2_decap_8 FILLER_98_566 ();
 sg13g2_decap_8 FILLER_98_573 ();
 sg13g2_decap_8 FILLER_98_580 ();
 sg13g2_decap_4 FILLER_98_587 ();
 sg13g2_decap_8 FILLER_98_595 ();
 sg13g2_decap_8 FILLER_98_602 ();
 sg13g2_decap_8 FILLER_98_609 ();
 sg13g2_decap_4 FILLER_98_616 ();
 sg13g2_decap_8 FILLER_98_626 ();
 sg13g2_decap_8 FILLER_98_633 ();
 sg13g2_fill_2 FILLER_98_640 ();
 sg13g2_fill_1 FILLER_98_642 ();
 sg13g2_decap_8 FILLER_98_647 ();
 sg13g2_fill_1 FILLER_98_654 ();
 sg13g2_decap_4 FILLER_98_660 ();
 sg13g2_decap_8 FILLER_98_672 ();
 sg13g2_decap_8 FILLER_98_679 ();
 sg13g2_decap_4 FILLER_98_686 ();
 sg13g2_fill_1 FILLER_98_690 ();
 sg13g2_decap_4 FILLER_98_695 ();
 sg13g2_fill_2 FILLER_98_699 ();
 sg13g2_decap_8 FILLER_98_706 ();
 sg13g2_decap_4 FILLER_98_713 ();
 sg13g2_fill_1 FILLER_98_717 ();
 sg13g2_decap_8 FILLER_98_739 ();
 sg13g2_decap_8 FILLER_98_746 ();
 sg13g2_fill_2 FILLER_98_753 ();
 sg13g2_decap_8 FILLER_98_759 ();
 sg13g2_decap_8 FILLER_98_766 ();
 sg13g2_decap_8 FILLER_98_773 ();
 sg13g2_decap_8 FILLER_98_780 ();
 sg13g2_decap_8 FILLER_98_787 ();
 sg13g2_decap_8 FILLER_98_794 ();
 sg13g2_decap_8 FILLER_98_801 ();
 sg13g2_decap_8 FILLER_98_808 ();
 sg13g2_decap_4 FILLER_98_815 ();
 sg13g2_fill_2 FILLER_98_819 ();
 sg13g2_decap_8 FILLER_98_825 ();
 sg13g2_decap_8 FILLER_98_832 ();
 sg13g2_decap_8 FILLER_98_839 ();
 sg13g2_decap_8 FILLER_98_846 ();
 sg13g2_decap_4 FILLER_98_853 ();
 sg13g2_decap_8 FILLER_98_896 ();
 sg13g2_decap_8 FILLER_98_906 ();
 sg13g2_decap_8 FILLER_98_913 ();
 sg13g2_decap_8 FILLER_98_920 ();
 sg13g2_decap_8 FILLER_98_927 ();
 sg13g2_decap_4 FILLER_98_934 ();
 sg13g2_fill_1 FILLER_98_938 ();
 sg13g2_decap_8 FILLER_98_948 ();
 sg13g2_decap_8 FILLER_98_955 ();
 sg13g2_decap_8 FILLER_98_962 ();
 sg13g2_decap_4 FILLER_98_969 ();
 sg13g2_fill_1 FILLER_98_973 ();
 sg13g2_fill_1 FILLER_98_978 ();
 sg13g2_decap_8 FILLER_98_992 ();
 sg13g2_decap_8 FILLER_98_999 ();
 sg13g2_decap_8 FILLER_98_1006 ();
 sg13g2_fill_2 FILLER_98_1013 ();
 sg13g2_decap_8 FILLER_98_1023 ();
 sg13g2_decap_8 FILLER_98_1030 ();
 sg13g2_fill_2 FILLER_98_1037 ();
 sg13g2_decap_4 FILLER_98_1047 ();
 sg13g2_fill_1 FILLER_98_1051 ();
 sg13g2_decap_8 FILLER_98_1056 ();
 sg13g2_decap_8 FILLER_98_1063 ();
 sg13g2_fill_2 FILLER_98_1070 ();
 sg13g2_fill_1 FILLER_98_1072 ();
 sg13g2_fill_1 FILLER_98_1079 ();
 sg13g2_decap_8 FILLER_98_1105 ();
 sg13g2_decap_4 FILLER_98_1112 ();
 sg13g2_fill_1 FILLER_98_1116 ();
 sg13g2_decap_8 FILLER_98_1121 ();
 sg13g2_decap_8 FILLER_98_1128 ();
 sg13g2_decap_4 FILLER_98_1135 ();
 sg13g2_fill_1 FILLER_98_1139 ();
 sg13g2_decap_8 FILLER_98_1153 ();
 sg13g2_decap_8 FILLER_98_1160 ();
 sg13g2_fill_2 FILLER_98_1175 ();
 sg13g2_decap_4 FILLER_98_1195 ();
 sg13g2_fill_1 FILLER_98_1199 ();
 sg13g2_decap_4 FILLER_98_1208 ();
 sg13g2_fill_2 FILLER_98_1212 ();
 sg13g2_decap_4 FILLER_98_1240 ();
 sg13g2_fill_1 FILLER_98_1244 ();
 sg13g2_fill_1 FILLER_98_1271 ();
 sg13g2_decap_8 FILLER_98_1285 ();
 sg13g2_decap_8 FILLER_98_1292 ();
 sg13g2_decap_8 FILLER_98_1299 ();
 sg13g2_decap_8 FILLER_98_1306 ();
 sg13g2_decap_8 FILLER_98_1313 ();
 sg13g2_decap_8 FILLER_98_1320 ();
 sg13g2_decap_8 FILLER_98_1327 ();
 sg13g2_decap_8 FILLER_98_1334 ();
 sg13g2_decap_8 FILLER_98_1341 ();
 sg13g2_decap_8 FILLER_98_1348 ();
 sg13g2_decap_8 FILLER_98_1355 ();
 sg13g2_decap_8 FILLER_98_1362 ();
 sg13g2_decap_8 FILLER_98_1369 ();
 sg13g2_decap_8 FILLER_98_1376 ();
 sg13g2_fill_2 FILLER_98_1383 ();
 sg13g2_fill_1 FILLER_98_1385 ();
 sg13g2_fill_1 FILLER_98_1390 ();
 sg13g2_decap_8 FILLER_98_1404 ();
 sg13g2_fill_2 FILLER_98_1411 ();
 sg13g2_decap_8 FILLER_98_1453 ();
 sg13g2_fill_2 FILLER_98_1460 ();
 sg13g2_decap_8 FILLER_98_1473 ();
 sg13g2_decap_8 FILLER_98_1480 ();
 sg13g2_decap_8 FILLER_98_1487 ();
 sg13g2_decap_8 FILLER_98_1494 ();
 sg13g2_fill_2 FILLER_98_1501 ();
 sg13g2_fill_1 FILLER_98_1503 ();
 sg13g2_fill_2 FILLER_98_1508 ();
 sg13g2_decap_8 FILLER_98_1520 ();
 sg13g2_decap_8 FILLER_98_1527 ();
 sg13g2_decap_4 FILLER_98_1534 ();
 sg13g2_fill_1 FILLER_98_1538 ();
 sg13g2_decap_8 FILLER_98_1551 ();
 sg13g2_decap_4 FILLER_98_1558 ();
 sg13g2_decap_8 FILLER_98_1571 ();
 sg13g2_fill_1 FILLER_98_1578 ();
 sg13g2_decap_8 FILLER_98_1587 ();
 sg13g2_decap_8 FILLER_98_1594 ();
 sg13g2_decap_8 FILLER_98_1601 ();
 sg13g2_decap_8 FILLER_98_1608 ();
 sg13g2_decap_4 FILLER_98_1615 ();
 sg13g2_decap_8 FILLER_98_1627 ();
 sg13g2_decap_4 FILLER_98_1634 ();
 sg13g2_fill_2 FILLER_98_1646 ();
 sg13g2_fill_1 FILLER_98_1648 ();
 sg13g2_decap_8 FILLER_98_1659 ();
 sg13g2_decap_8 FILLER_98_1666 ();
 sg13g2_decap_8 FILLER_98_1673 ();
 sg13g2_decap_8 FILLER_98_1680 ();
 sg13g2_decap_8 FILLER_98_1687 ();
 sg13g2_decap_8 FILLER_98_1694 ();
 sg13g2_decap_4 FILLER_98_1701 ();
 sg13g2_fill_2 FILLER_98_1705 ();
 sg13g2_decap_8 FILLER_98_1727 ();
 sg13g2_decap_8 FILLER_98_1734 ();
 sg13g2_decap_8 FILLER_98_1741 ();
 sg13g2_decap_8 FILLER_98_1748 ();
 sg13g2_decap_8 FILLER_98_1755 ();
 sg13g2_decap_4 FILLER_98_1762 ();
 sg13g2_fill_2 FILLER_98_1766 ();
 sg13g2_decap_8 FILLER_99_0 ();
 sg13g2_decap_8 FILLER_99_7 ();
 sg13g2_decap_8 FILLER_99_14 ();
 sg13g2_decap_8 FILLER_99_21 ();
 sg13g2_decap_8 FILLER_99_28 ();
 sg13g2_decap_8 FILLER_99_35 ();
 sg13g2_decap_8 FILLER_99_42 ();
 sg13g2_decap_4 FILLER_99_49 ();
 sg13g2_fill_2 FILLER_99_53 ();
 sg13g2_fill_1 FILLER_99_63 ();
 sg13g2_decap_8 FILLER_99_83 ();
 sg13g2_decap_8 FILLER_99_90 ();
 sg13g2_decap_8 FILLER_99_97 ();
 sg13g2_decap_8 FILLER_99_112 ();
 sg13g2_decap_8 FILLER_99_119 ();
 sg13g2_fill_2 FILLER_99_146 ();
 sg13g2_decap_8 FILLER_99_156 ();
 sg13g2_fill_2 FILLER_99_163 ();
 sg13g2_fill_1 FILLER_99_165 ();
 sg13g2_decap_8 FILLER_99_174 ();
 sg13g2_decap_8 FILLER_99_181 ();
 sg13g2_decap_8 FILLER_99_188 ();
 sg13g2_decap_8 FILLER_99_195 ();
 sg13g2_fill_2 FILLER_99_202 ();
 sg13g2_decap_8 FILLER_99_234 ();
 sg13g2_decap_4 FILLER_99_241 ();
 sg13g2_fill_1 FILLER_99_245 ();
 sg13g2_decap_8 FILLER_99_262 ();
 sg13g2_fill_1 FILLER_99_269 ();
 sg13g2_decap_8 FILLER_99_275 ();
 sg13g2_decap_8 FILLER_99_282 ();
 sg13g2_decap_8 FILLER_99_289 ();
 sg13g2_decap_8 FILLER_99_296 ();
 sg13g2_fill_2 FILLER_99_303 ();
 sg13g2_fill_1 FILLER_99_305 ();
 sg13g2_decap_8 FILLER_99_341 ();
 sg13g2_decap_8 FILLER_99_348 ();
 sg13g2_fill_2 FILLER_99_355 ();
 sg13g2_fill_1 FILLER_99_357 ();
 sg13g2_fill_2 FILLER_99_403 ();
 sg13g2_fill_1 FILLER_99_405 ();
 sg13g2_decap_8 FILLER_99_434 ();
 sg13g2_decap_8 FILLER_99_441 ();
 sg13g2_decap_8 FILLER_99_448 ();
 sg13g2_decap_8 FILLER_99_479 ();
 sg13g2_decap_8 FILLER_99_486 ();
 sg13g2_decap_8 FILLER_99_493 ();
 sg13g2_decap_8 FILLER_99_500 ();
 sg13g2_fill_1 FILLER_99_507 ();
 sg13g2_fill_1 FILLER_99_512 ();
 sg13g2_fill_2 FILLER_99_521 ();
 sg13g2_decap_8 FILLER_99_543 ();
 sg13g2_decap_8 FILLER_99_550 ();
 sg13g2_decap_8 FILLER_99_557 ();
 sg13g2_decap_8 FILLER_99_564 ();
 sg13g2_decap_8 FILLER_99_571 ();
 sg13g2_decap_8 FILLER_99_578 ();
 sg13g2_decap_8 FILLER_99_585 ();
 sg13g2_fill_2 FILLER_99_592 ();
 sg13g2_decap_8 FILLER_99_602 ();
 sg13g2_decap_4 FILLER_99_609 ();
 sg13g2_fill_1 FILLER_99_613 ();
 sg13g2_decap_8 FILLER_99_619 ();
 sg13g2_decap_8 FILLER_99_626 ();
 sg13g2_decap_8 FILLER_99_633 ();
 sg13g2_decap_8 FILLER_99_640 ();
 sg13g2_decap_8 FILLER_99_647 ();
 sg13g2_fill_2 FILLER_99_654 ();
 sg13g2_fill_1 FILLER_99_656 ();
 sg13g2_decap_8 FILLER_99_665 ();
 sg13g2_decap_8 FILLER_99_680 ();
 sg13g2_decap_8 FILLER_99_687 ();
 sg13g2_decap_8 FILLER_99_694 ();
 sg13g2_decap_8 FILLER_99_701 ();
 sg13g2_decap_8 FILLER_99_708 ();
 sg13g2_fill_2 FILLER_99_715 ();
 sg13g2_fill_1 FILLER_99_717 ();
 sg13g2_decap_4 FILLER_99_740 ();
 sg13g2_decap_8 FILLER_99_770 ();
 sg13g2_decap_8 FILLER_99_777 ();
 sg13g2_decap_8 FILLER_99_784 ();
 sg13g2_decap_8 FILLER_99_791 ();
 sg13g2_decap_8 FILLER_99_798 ();
 sg13g2_decap_4 FILLER_99_805 ();
 sg13g2_fill_2 FILLER_99_809 ();
 sg13g2_decap_8 FILLER_99_837 ();
 sg13g2_decap_8 FILLER_99_844 ();
 sg13g2_decap_8 FILLER_99_851 ();
 sg13g2_decap_8 FILLER_99_858 ();
 sg13g2_fill_2 FILLER_99_865 ();
 sg13g2_fill_1 FILLER_99_867 ();
 sg13g2_decap_8 FILLER_99_872 ();
 sg13g2_decap_8 FILLER_99_879 ();
 sg13g2_decap_8 FILLER_99_886 ();
 sg13g2_fill_2 FILLER_99_898 ();
 sg13g2_decap_8 FILLER_99_910 ();
 sg13g2_decap_8 FILLER_99_917 ();
 sg13g2_decap_8 FILLER_99_924 ();
 sg13g2_decap_8 FILLER_99_931 ();
 sg13g2_decap_8 FILLER_99_938 ();
 sg13g2_decap_8 FILLER_99_945 ();
 sg13g2_decap_8 FILLER_99_952 ();
 sg13g2_decap_8 FILLER_99_959 ();
 sg13g2_decap_8 FILLER_99_966 ();
 sg13g2_decap_8 FILLER_99_973 ();
 sg13g2_decap_8 FILLER_99_988 ();
 sg13g2_decap_8 FILLER_99_995 ();
 sg13g2_decap_4 FILLER_99_1002 ();
 sg13g2_fill_1 FILLER_99_1006 ();
 sg13g2_decap_8 FILLER_99_1020 ();
 sg13g2_decap_8 FILLER_99_1027 ();
 sg13g2_decap_4 FILLER_99_1034 ();
 sg13g2_decap_4 FILLER_99_1042 ();
 sg13g2_fill_2 FILLER_99_1046 ();
 sg13g2_decap_8 FILLER_99_1079 ();
 sg13g2_decap_4 FILLER_99_1086 ();
 sg13g2_decap_8 FILLER_99_1096 ();
 sg13g2_decap_8 FILLER_99_1103 ();
 sg13g2_fill_2 FILLER_99_1110 ();
 sg13g2_decap_8 FILLER_99_1143 ();
 sg13g2_decap_8 FILLER_99_1163 ();
 sg13g2_decap_8 FILLER_99_1170 ();
 sg13g2_decap_8 FILLER_99_1177 ();
 sg13g2_decap_4 FILLER_99_1184 ();
 sg13g2_fill_2 FILLER_99_1188 ();
 sg13g2_decap_8 FILLER_99_1203 ();
 sg13g2_decap_8 FILLER_99_1210 ();
 sg13g2_decap_8 FILLER_99_1217 ();
 sg13g2_fill_2 FILLER_99_1224 ();
 sg13g2_fill_1 FILLER_99_1226 ();
 sg13g2_decap_8 FILLER_99_1236 ();
 sg13g2_decap_8 FILLER_99_1243 ();
 sg13g2_decap_4 FILLER_99_1250 ();
 sg13g2_fill_1 FILLER_99_1254 ();
 sg13g2_decap_8 FILLER_99_1259 ();
 sg13g2_decap_8 FILLER_99_1266 ();
 sg13g2_decap_8 FILLER_99_1273 ();
 sg13g2_decap_8 FILLER_99_1280 ();
 sg13g2_decap_8 FILLER_99_1287 ();
 sg13g2_decap_8 FILLER_99_1294 ();
 sg13g2_decap_4 FILLER_99_1301 ();
 sg13g2_decap_8 FILLER_99_1308 ();
 sg13g2_fill_2 FILLER_99_1315 ();
 sg13g2_decap_8 FILLER_99_1323 ();
 sg13g2_decap_8 FILLER_99_1330 ();
 sg13g2_decap_8 FILLER_99_1337 ();
 sg13g2_decap_8 FILLER_99_1344 ();
 sg13g2_decap_4 FILLER_99_1351 ();
 sg13g2_decap_4 FILLER_99_1368 ();
 sg13g2_fill_2 FILLER_99_1372 ();
 sg13g2_decap_8 FILLER_99_1379 ();
 sg13g2_decap_8 FILLER_99_1386 ();
 sg13g2_fill_2 FILLER_99_1393 ();
 sg13g2_fill_1 FILLER_99_1395 ();
 sg13g2_decap_8 FILLER_99_1405 ();
 sg13g2_decap_8 FILLER_99_1412 ();
 sg13g2_decap_4 FILLER_99_1419 ();
 sg13g2_fill_1 FILLER_99_1423 ();
 sg13g2_decap_8 FILLER_99_1428 ();
 sg13g2_decap_8 FILLER_99_1435 ();
 sg13g2_decap_8 FILLER_99_1442 ();
 sg13g2_decap_8 FILLER_99_1449 ();
 sg13g2_fill_1 FILLER_99_1456 ();
 sg13g2_decap_8 FILLER_99_1465 ();
 sg13g2_decap_8 FILLER_99_1472 ();
 sg13g2_fill_2 FILLER_99_1479 ();
 sg13g2_decap_8 FILLER_99_1489 ();
 sg13g2_decap_8 FILLER_99_1496 ();
 sg13g2_decap_8 FILLER_99_1503 ();
 sg13g2_decap_8 FILLER_99_1510 ();
 sg13g2_decap_8 FILLER_99_1517 ();
 sg13g2_decap_8 FILLER_99_1524 ();
 sg13g2_decap_8 FILLER_99_1531 ();
 sg13g2_decap_4 FILLER_99_1538 ();
 sg13g2_fill_2 FILLER_99_1545 ();
 sg13g2_decap_8 FILLER_99_1582 ();
 sg13g2_decap_8 FILLER_99_1589 ();
 sg13g2_decap_8 FILLER_99_1596 ();
 sg13g2_fill_2 FILLER_99_1603 ();
 sg13g2_fill_1 FILLER_99_1605 ();
 sg13g2_decap_8 FILLER_99_1610 ();
 sg13g2_decap_8 FILLER_99_1617 ();
 sg13g2_decap_4 FILLER_99_1624 ();
 sg13g2_decap_8 FILLER_99_1632 ();
 sg13g2_decap_4 FILLER_99_1647 ();
 sg13g2_fill_2 FILLER_99_1651 ();
 sg13g2_decap_8 FILLER_99_1658 ();
 sg13g2_decap_8 FILLER_99_1665 ();
 sg13g2_decap_8 FILLER_99_1672 ();
 sg13g2_decap_8 FILLER_99_1679 ();
 sg13g2_decap_4 FILLER_99_1686 ();
 sg13g2_fill_2 FILLER_99_1690 ();
 sg13g2_decap_8 FILLER_99_1708 ();
 sg13g2_decap_8 FILLER_99_1715 ();
 sg13g2_decap_4 FILLER_99_1722 ();
 sg13g2_fill_2 FILLER_99_1726 ();
 sg13g2_decap_8 FILLER_99_1737 ();
 sg13g2_decap_8 FILLER_99_1744 ();
 sg13g2_decap_8 FILLER_99_1751 ();
 sg13g2_decap_8 FILLER_99_1758 ();
 sg13g2_fill_2 FILLER_99_1765 ();
 sg13g2_fill_1 FILLER_99_1767 ();
 sg13g2_decap_8 FILLER_100_0 ();
 sg13g2_decap_8 FILLER_100_7 ();
 sg13g2_decap_8 FILLER_100_14 ();
 sg13g2_decap_8 FILLER_100_21 ();
 sg13g2_decap_8 FILLER_100_28 ();
 sg13g2_decap_8 FILLER_100_35 ();
 sg13g2_decap_8 FILLER_100_42 ();
 sg13g2_decap_4 FILLER_100_49 ();
 sg13g2_decap_8 FILLER_100_82 ();
 sg13g2_decap_8 FILLER_100_89 ();
 sg13g2_decap_8 FILLER_100_96 ();
 sg13g2_decap_8 FILLER_100_103 ();
 sg13g2_fill_2 FILLER_100_110 ();
 sg13g2_decap_4 FILLER_100_125 ();
 sg13g2_decap_4 FILLER_100_146 ();
 sg13g2_decap_8 FILLER_100_170 ();
 sg13g2_decap_8 FILLER_100_177 ();
 sg13g2_decap_8 FILLER_100_184 ();
 sg13g2_decap_8 FILLER_100_191 ();
 sg13g2_decap_8 FILLER_100_198 ();
 sg13g2_decap_4 FILLER_100_205 ();
 sg13g2_fill_2 FILLER_100_209 ();
 sg13g2_fill_1 FILLER_100_217 ();
 sg13g2_decap_8 FILLER_100_229 ();
 sg13g2_decap_8 FILLER_100_236 ();
 sg13g2_decap_8 FILLER_100_243 ();
 sg13g2_decap_8 FILLER_100_250 ();
 sg13g2_decap_4 FILLER_100_257 ();
 sg13g2_fill_2 FILLER_100_261 ();
 sg13g2_decap_8 FILLER_100_291 ();
 sg13g2_decap_8 FILLER_100_298 ();
 sg13g2_decap_8 FILLER_100_305 ();
 sg13g2_fill_2 FILLER_100_312 ();
 sg13g2_fill_2 FILLER_100_322 ();
 sg13g2_decap_8 FILLER_100_332 ();
 sg13g2_decap_8 FILLER_100_339 ();
 sg13g2_decap_8 FILLER_100_346 ();
 sg13g2_decap_8 FILLER_100_353 ();
 sg13g2_decap_4 FILLER_100_360 ();
 sg13g2_decap_8 FILLER_100_380 ();
 sg13g2_decap_8 FILLER_100_387 ();
 sg13g2_fill_2 FILLER_100_394 ();
 sg13g2_fill_1 FILLER_100_396 ();
 sg13g2_decap_8 FILLER_100_405 ();
 sg13g2_fill_1 FILLER_100_412 ();
 sg13g2_decap_4 FILLER_100_425 ();
 sg13g2_fill_1 FILLER_100_429 ();
 sg13g2_decap_8 FILLER_100_434 ();
 sg13g2_decap_8 FILLER_100_441 ();
 sg13g2_decap_8 FILLER_100_448 ();
 sg13g2_decap_8 FILLER_100_458 ();
 sg13g2_decap_4 FILLER_100_465 ();
 sg13g2_fill_2 FILLER_100_469 ();
 sg13g2_decap_8 FILLER_100_475 ();
 sg13g2_decap_8 FILLER_100_482 ();
 sg13g2_decap_4 FILLER_100_489 ();
 sg13g2_fill_2 FILLER_100_509 ();
 sg13g2_fill_1 FILLER_100_511 ();
 sg13g2_decap_8 FILLER_100_528 ();
 sg13g2_decap_8 FILLER_100_535 ();
 sg13g2_decap_8 FILLER_100_542 ();
 sg13g2_fill_2 FILLER_100_549 ();
 sg13g2_fill_1 FILLER_100_551 ();
 sg13g2_decap_8 FILLER_100_565 ();
 sg13g2_decap_8 FILLER_100_572 ();
 sg13g2_decap_8 FILLER_100_579 ();
 sg13g2_decap_8 FILLER_100_586 ();
 sg13g2_decap_8 FILLER_100_593 ();
 sg13g2_decap_8 FILLER_100_600 ();
 sg13g2_decap_8 FILLER_100_607 ();
 sg13g2_decap_8 FILLER_100_614 ();
 sg13g2_decap_8 FILLER_100_621 ();
 sg13g2_decap_8 FILLER_100_628 ();
 sg13g2_decap_8 FILLER_100_635 ();
 sg13g2_decap_8 FILLER_100_642 ();
 sg13g2_fill_2 FILLER_100_649 ();
 sg13g2_fill_1 FILLER_100_651 ();
 sg13g2_fill_2 FILLER_100_665 ();
 sg13g2_decap_8 FILLER_100_684 ();
 sg13g2_decap_8 FILLER_100_691 ();
 sg13g2_decap_8 FILLER_100_698 ();
 sg13g2_decap_8 FILLER_100_705 ();
 sg13g2_decap_8 FILLER_100_712 ();
 sg13g2_decap_4 FILLER_100_719 ();
 sg13g2_fill_1 FILLER_100_723 ();
 sg13g2_decap_4 FILLER_100_730 ();
 sg13g2_fill_2 FILLER_100_734 ();
 sg13g2_decap_8 FILLER_100_741 ();
 sg13g2_decap_8 FILLER_100_748 ();
 sg13g2_decap_8 FILLER_100_755 ();
 sg13g2_fill_1 FILLER_100_762 ();
 sg13g2_fill_2 FILLER_100_771 ();
 sg13g2_fill_1 FILLER_100_773 ();
 sg13g2_decap_8 FILLER_100_782 ();
 sg13g2_decap_8 FILLER_100_789 ();
 sg13g2_decap_8 FILLER_100_796 ();
 sg13g2_decap_8 FILLER_100_803 ();
 sg13g2_decap_4 FILLER_100_810 ();
 sg13g2_fill_2 FILLER_100_814 ();
 sg13g2_decap_8 FILLER_100_820 ();
 sg13g2_decap_8 FILLER_100_827 ();
 sg13g2_decap_8 FILLER_100_834 ();
 sg13g2_decap_8 FILLER_100_841 ();
 sg13g2_decap_4 FILLER_100_848 ();
 sg13g2_decap_8 FILLER_100_860 ();
 sg13g2_decap_8 FILLER_100_867 ();
 sg13g2_decap_8 FILLER_100_874 ();
 sg13g2_decap_8 FILLER_100_881 ();
 sg13g2_decap_8 FILLER_100_888 ();
 sg13g2_decap_8 FILLER_100_895 ();
 sg13g2_fill_1 FILLER_100_902 ();
 sg13g2_decap_8 FILLER_100_920 ();
 sg13g2_decap_8 FILLER_100_927 ();
 sg13g2_decap_8 FILLER_100_934 ();
 sg13g2_decap_8 FILLER_100_941 ();
 sg13g2_decap_8 FILLER_100_948 ();
 sg13g2_fill_2 FILLER_100_955 ();
 sg13g2_decap_8 FILLER_100_965 ();
 sg13g2_decap_8 FILLER_100_972 ();
 sg13g2_decap_8 FILLER_100_979 ();
 sg13g2_decap_8 FILLER_100_986 ();
 sg13g2_decap_8 FILLER_100_993 ();
 sg13g2_decap_8 FILLER_100_1000 ();
 sg13g2_decap_8 FILLER_100_1007 ();
 sg13g2_fill_2 FILLER_100_1014 ();
 sg13g2_decap_8 FILLER_100_1029 ();
 sg13g2_decap_8 FILLER_100_1036 ();
 sg13g2_decap_8 FILLER_100_1043 ();
 sg13g2_decap_8 FILLER_100_1050 ();
 sg13g2_decap_8 FILLER_100_1057 ();
 sg13g2_decap_8 FILLER_100_1068 ();
 sg13g2_fill_2 FILLER_100_1075 ();
 sg13g2_fill_1 FILLER_100_1077 ();
 sg13g2_decap_4 FILLER_100_1097 ();
 sg13g2_fill_1 FILLER_100_1101 ();
 sg13g2_decap_8 FILLER_100_1119 ();
 sg13g2_fill_2 FILLER_100_1126 ();
 sg13g2_decap_8 FILLER_100_1132 ();
 sg13g2_decap_8 FILLER_100_1139 ();
 sg13g2_fill_1 FILLER_100_1146 ();
 sg13g2_decap_8 FILLER_100_1156 ();
 sg13g2_decap_8 FILLER_100_1163 ();
 sg13g2_decap_8 FILLER_100_1170 ();
 sg13g2_decap_4 FILLER_100_1177 ();
 sg13g2_fill_2 FILLER_100_1190 ();
 sg13g2_fill_1 FILLER_100_1192 ();
 sg13g2_decap_8 FILLER_100_1201 ();
 sg13g2_decap_8 FILLER_100_1208 ();
 sg13g2_decap_8 FILLER_100_1215 ();
 sg13g2_decap_8 FILLER_100_1222 ();
 sg13g2_decap_8 FILLER_100_1229 ();
 sg13g2_decap_8 FILLER_100_1236 ();
 sg13g2_decap_8 FILLER_100_1243 ();
 sg13g2_decap_8 FILLER_100_1250 ();
 sg13g2_decap_8 FILLER_100_1257 ();
 sg13g2_decap_8 FILLER_100_1264 ();
 sg13g2_decap_8 FILLER_100_1271 ();
 sg13g2_decap_8 FILLER_100_1278 ();
 sg13g2_decap_4 FILLER_100_1285 ();
 sg13g2_fill_1 FILLER_100_1289 ();
 sg13g2_decap_8 FILLER_100_1293 ();
 sg13g2_fill_2 FILLER_100_1300 ();
 sg13g2_fill_1 FILLER_100_1313 ();
 sg13g2_decap_8 FILLER_100_1335 ();
 sg13g2_decap_8 FILLER_100_1342 ();
 sg13g2_fill_2 FILLER_100_1349 ();
 sg13g2_fill_1 FILLER_100_1351 ();
 sg13g2_decap_4 FILLER_100_1387 ();
 sg13g2_fill_2 FILLER_100_1391 ();
 sg13g2_decap_8 FILLER_100_1409 ();
 sg13g2_decap_8 FILLER_100_1416 ();
 sg13g2_decap_8 FILLER_100_1423 ();
 sg13g2_decap_8 FILLER_100_1430 ();
 sg13g2_decap_8 FILLER_100_1437 ();
 sg13g2_decap_8 FILLER_100_1444 ();
 sg13g2_fill_2 FILLER_100_1451 ();
 sg13g2_fill_1 FILLER_100_1453 ();
 sg13g2_decap_8 FILLER_100_1478 ();
 sg13g2_decap_8 FILLER_100_1485 ();
 sg13g2_decap_8 FILLER_100_1492 ();
 sg13g2_decap_8 FILLER_100_1499 ();
 sg13g2_decap_8 FILLER_100_1529 ();
 sg13g2_decap_8 FILLER_100_1536 ();
 sg13g2_decap_8 FILLER_100_1543 ();
 sg13g2_decap_8 FILLER_100_1550 ();
 sg13g2_decap_4 FILLER_100_1557 ();
 sg13g2_fill_1 FILLER_100_1561 ();
 sg13g2_decap_8 FILLER_100_1566 ();
 sg13g2_decap_8 FILLER_100_1573 ();
 sg13g2_decap_8 FILLER_100_1580 ();
 sg13g2_decap_8 FILLER_100_1587 ();
 sg13g2_decap_8 FILLER_100_1594 ();
 sg13g2_decap_8 FILLER_100_1601 ();
 sg13g2_decap_8 FILLER_100_1608 ();
 sg13g2_decap_4 FILLER_100_1615 ();
 sg13g2_fill_1 FILLER_100_1619 ();
 sg13g2_decap_4 FILLER_100_1624 ();
 sg13g2_fill_2 FILLER_100_1628 ();
 sg13g2_decap_8 FILLER_100_1635 ();
 sg13g2_decap_4 FILLER_100_1642 ();
 sg13g2_fill_2 FILLER_100_1646 ();
 sg13g2_fill_2 FILLER_100_1661 ();
 sg13g2_fill_1 FILLER_100_1663 ();
 sg13g2_decap_8 FILLER_100_1672 ();
 sg13g2_decap_8 FILLER_100_1679 ();
 sg13g2_decap_8 FILLER_100_1686 ();
 sg13g2_decap_8 FILLER_100_1693 ();
 sg13g2_fill_2 FILLER_100_1709 ();
 sg13g2_fill_1 FILLER_100_1711 ();
 sg13g2_fill_1 FILLER_100_1730 ();
 sg13g2_fill_1 FILLER_100_1741 ();
 sg13g2_decap_8 FILLER_100_1750 ();
 sg13g2_decap_8 FILLER_100_1757 ();
 sg13g2_decap_4 FILLER_100_1764 ();
 sg13g2_decap_8 FILLER_101_0 ();
 sg13g2_decap_8 FILLER_101_7 ();
 sg13g2_decap_8 FILLER_101_14 ();
 sg13g2_fill_1 FILLER_101_21 ();
 sg13g2_fill_2 FILLER_101_31 ();
 sg13g2_decap_8 FILLER_101_38 ();
 sg13g2_decap_4 FILLER_101_45 ();
 sg13g2_fill_2 FILLER_101_49 ();
 sg13g2_decap_8 FILLER_101_55 ();
 sg13g2_decap_4 FILLER_101_62 ();
 sg13g2_fill_2 FILLER_101_66 ();
 sg13g2_decap_8 FILLER_101_93 ();
 sg13g2_decap_8 FILLER_101_100 ();
 sg13g2_decap_8 FILLER_101_107 ();
 sg13g2_decap_8 FILLER_101_114 ();
 sg13g2_decap_4 FILLER_101_129 ();
 sg13g2_fill_1 FILLER_101_133 ();
 sg13g2_decap_8 FILLER_101_141 ();
 sg13g2_decap_8 FILLER_101_148 ();
 sg13g2_decap_8 FILLER_101_155 ();
 sg13g2_decap_4 FILLER_101_162 ();
 sg13g2_decap_8 FILLER_101_178 ();
 sg13g2_decap_8 FILLER_101_185 ();
 sg13g2_decap_8 FILLER_101_192 ();
 sg13g2_decap_8 FILLER_101_199 ();
 sg13g2_decap_8 FILLER_101_206 ();
 sg13g2_decap_8 FILLER_101_213 ();
 sg13g2_decap_4 FILLER_101_220 ();
 sg13g2_fill_2 FILLER_101_224 ();
 sg13g2_decap_8 FILLER_101_232 ();
 sg13g2_decap_8 FILLER_101_239 ();
 sg13g2_decap_8 FILLER_101_246 ();
 sg13g2_decap_8 FILLER_101_253 ();
 sg13g2_decap_8 FILLER_101_260 ();
 sg13g2_decap_8 FILLER_101_267 ();
 sg13g2_fill_2 FILLER_101_274 ();
 sg13g2_fill_1 FILLER_101_276 ();
 sg13g2_decap_8 FILLER_101_286 ();
 sg13g2_decap_8 FILLER_101_293 ();
 sg13g2_decap_8 FILLER_101_300 ();
 sg13g2_decap_8 FILLER_101_307 ();
 sg13g2_decap_8 FILLER_101_314 ();
 sg13g2_decap_8 FILLER_101_321 ();
 sg13g2_fill_2 FILLER_101_328 ();
 sg13g2_fill_1 FILLER_101_330 ();
 sg13g2_decap_8 FILLER_101_339 ();
 sg13g2_decap_8 FILLER_101_346 ();
 sg13g2_decap_4 FILLER_101_353 ();
 sg13g2_fill_2 FILLER_101_357 ();
 sg13g2_decap_8 FILLER_101_379 ();
 sg13g2_decap_8 FILLER_101_386 ();
 sg13g2_decap_8 FILLER_101_393 ();
 sg13g2_decap_8 FILLER_101_400 ();
 sg13g2_decap_8 FILLER_101_407 ();
 sg13g2_decap_8 FILLER_101_414 ();
 sg13g2_decap_8 FILLER_101_421 ();
 sg13g2_decap_8 FILLER_101_428 ();
 sg13g2_decap_8 FILLER_101_435 ();
 sg13g2_decap_4 FILLER_101_442 ();
 sg13g2_fill_1 FILLER_101_446 ();
 sg13g2_decap_8 FILLER_101_463 ();
 sg13g2_decap_4 FILLER_101_470 ();
 sg13g2_decap_8 FILLER_101_482 ();
 sg13g2_decap_8 FILLER_101_489 ();
 sg13g2_fill_2 FILLER_101_504 ();
 sg13g2_decap_8 FILLER_101_534 ();
 sg13g2_decap_8 FILLER_101_541 ();
 sg13g2_decap_8 FILLER_101_548 ();
 sg13g2_decap_8 FILLER_101_555 ();
 sg13g2_decap_4 FILLER_101_562 ();
 sg13g2_fill_2 FILLER_101_566 ();
 sg13g2_decap_4 FILLER_101_582 ();
 sg13g2_decap_8 FILLER_101_607 ();
 sg13g2_decap_8 FILLER_101_614 ();
 sg13g2_decap_8 FILLER_101_621 ();
 sg13g2_decap_8 FILLER_101_628 ();
 sg13g2_decap_8 FILLER_101_635 ();
 sg13g2_decap_8 FILLER_101_642 ();
 sg13g2_fill_2 FILLER_101_649 ();
 sg13g2_fill_1 FILLER_101_651 ();
 sg13g2_decap_8 FILLER_101_664 ();
 sg13g2_decap_8 FILLER_101_671 ();
 sg13g2_decap_8 FILLER_101_678 ();
 sg13g2_decap_4 FILLER_101_685 ();
 sg13g2_decap_8 FILLER_101_693 ();
 sg13g2_decap_8 FILLER_101_700 ();
 sg13g2_decap_4 FILLER_101_707 ();
 sg13g2_fill_2 FILLER_101_711 ();
 sg13g2_decap_8 FILLER_101_754 ();
 sg13g2_decap_8 FILLER_101_761 ();
 sg13g2_decap_8 FILLER_101_768 ();
 sg13g2_decap_8 FILLER_101_775 ();
 sg13g2_decap_8 FILLER_101_782 ();
 sg13g2_decap_8 FILLER_101_789 ();
 sg13g2_decap_8 FILLER_101_796 ();
 sg13g2_decap_8 FILLER_101_839 ();
 sg13g2_decap_4 FILLER_101_846 ();
 sg13g2_fill_1 FILLER_101_850 ();
 sg13g2_fill_2 FILLER_101_855 ();
 sg13g2_decap_8 FILLER_101_870 ();
 sg13g2_decap_8 FILLER_101_877 ();
 sg13g2_decap_8 FILLER_101_884 ();
 sg13g2_decap_8 FILLER_101_891 ();
 sg13g2_fill_2 FILLER_101_898 ();
 sg13g2_fill_1 FILLER_101_900 ();
 sg13g2_decap_8 FILLER_101_940 ();
 sg13g2_fill_2 FILLER_101_947 ();
 sg13g2_fill_1 FILLER_101_949 ();
 sg13g2_fill_2 FILLER_101_959 ();
 sg13g2_fill_1 FILLER_101_961 ();
 sg13g2_decap_8 FILLER_101_975 ();
 sg13g2_decap_8 FILLER_101_982 ();
 sg13g2_decap_8 FILLER_101_989 ();
 sg13g2_decap_8 FILLER_101_996 ();
 sg13g2_fill_2 FILLER_101_1003 ();
 sg13g2_fill_1 FILLER_101_1005 ();
 sg13g2_decap_8 FILLER_101_1040 ();
 sg13g2_decap_8 FILLER_101_1047 ();
 sg13g2_decap_4 FILLER_101_1054 ();
 sg13g2_decap_8 FILLER_101_1071 ();
 sg13g2_decap_8 FILLER_101_1078 ();
 sg13g2_fill_2 FILLER_101_1085 ();
 sg13g2_decap_8 FILLER_101_1101 ();
 sg13g2_decap_8 FILLER_101_1108 ();
 sg13g2_decap_8 FILLER_101_1115 ();
 sg13g2_decap_8 FILLER_101_1122 ();
 sg13g2_decap_8 FILLER_101_1129 ();
 sg13g2_decap_8 FILLER_101_1136 ();
 sg13g2_decap_8 FILLER_101_1143 ();
 sg13g2_decap_8 FILLER_101_1150 ();
 sg13g2_decap_8 FILLER_101_1157 ();
 sg13g2_decap_8 FILLER_101_1164 ();
 sg13g2_decap_8 FILLER_101_1171 ();
 sg13g2_decap_8 FILLER_101_1178 ();
 sg13g2_decap_8 FILLER_101_1185 ();
 sg13g2_decap_8 FILLER_101_1192 ();
 sg13g2_decap_8 FILLER_101_1199 ();
 sg13g2_decap_8 FILLER_101_1206 ();
 sg13g2_decap_8 FILLER_101_1213 ();
 sg13g2_decap_8 FILLER_101_1220 ();
 sg13g2_decap_8 FILLER_101_1227 ();
 sg13g2_decap_8 FILLER_101_1234 ();
 sg13g2_decap_4 FILLER_101_1245 ();
 sg13g2_decap_8 FILLER_101_1272 ();
 sg13g2_decap_8 FILLER_101_1279 ();
 sg13g2_decap_4 FILLER_101_1286 ();
 sg13g2_decap_4 FILLER_101_1299 ();
 sg13g2_fill_2 FILLER_101_1303 ();
 sg13g2_fill_2 FILLER_101_1324 ();
 sg13g2_fill_1 FILLER_101_1326 ();
 sg13g2_decap_8 FILLER_101_1341 ();
 sg13g2_decap_4 FILLER_101_1348 ();
 sg13g2_decap_8 FILLER_101_1369 ();
 sg13g2_decap_8 FILLER_101_1376 ();
 sg13g2_decap_8 FILLER_101_1383 ();
 sg13g2_decap_8 FILLER_101_1390 ();
 sg13g2_decap_8 FILLER_101_1397 ();
 sg13g2_decap_8 FILLER_101_1404 ();
 sg13g2_decap_8 FILLER_101_1411 ();
 sg13g2_decap_8 FILLER_101_1418 ();
 sg13g2_decap_8 FILLER_101_1425 ();
 sg13g2_decap_8 FILLER_101_1432 ();
 sg13g2_decap_8 FILLER_101_1439 ();
 sg13g2_decap_8 FILLER_101_1446 ();
 sg13g2_decap_8 FILLER_101_1453 ();
 sg13g2_decap_8 FILLER_101_1460 ();
 sg13g2_decap_8 FILLER_101_1467 ();
 sg13g2_decap_8 FILLER_101_1474 ();
 sg13g2_decap_8 FILLER_101_1481 ();
 sg13g2_decap_8 FILLER_101_1488 ();
 sg13g2_decap_8 FILLER_101_1495 ();
 sg13g2_decap_8 FILLER_101_1502 ();
 sg13g2_fill_2 FILLER_101_1509 ();
 sg13g2_fill_1 FILLER_101_1511 ();
 sg13g2_decap_8 FILLER_101_1525 ();
 sg13g2_decap_8 FILLER_101_1532 ();
 sg13g2_decap_8 FILLER_101_1539 ();
 sg13g2_fill_2 FILLER_101_1546 ();
 sg13g2_fill_1 FILLER_101_1548 ();
 sg13g2_decap_8 FILLER_101_1552 ();
 sg13g2_decap_8 FILLER_101_1559 ();
 sg13g2_decap_8 FILLER_101_1566 ();
 sg13g2_decap_8 FILLER_101_1573 ();
 sg13g2_decap_8 FILLER_101_1580 ();
 sg13g2_decap_8 FILLER_101_1587 ();
 sg13g2_decap_8 FILLER_101_1594 ();
 sg13g2_decap_8 FILLER_101_1601 ();
 sg13g2_decap_8 FILLER_101_1636 ();
 sg13g2_decap_8 FILLER_101_1643 ();
 sg13g2_decap_4 FILLER_101_1650 ();
 sg13g2_fill_1 FILLER_101_1654 ();
 sg13g2_decap_8 FILLER_101_1660 ();
 sg13g2_decap_8 FILLER_101_1667 ();
 sg13g2_decap_8 FILLER_101_1674 ();
 sg13g2_decap_8 FILLER_101_1681 ();
 sg13g2_fill_1 FILLER_101_1688 ();
 sg13g2_decap_8 FILLER_101_1697 ();
 sg13g2_decap_8 FILLER_101_1708 ();
 sg13g2_decap_8 FILLER_101_1715 ();
 sg13g2_decap_8 FILLER_101_1722 ();
 sg13g2_fill_1 FILLER_101_1729 ();
 sg13g2_decap_8 FILLER_101_1758 ();
 sg13g2_fill_2 FILLER_101_1765 ();
 sg13g2_fill_1 FILLER_101_1767 ();
 sg13g2_decap_8 FILLER_102_0 ();
 sg13g2_decap_8 FILLER_102_7 ();
 sg13g2_fill_2 FILLER_102_14 ();
 sg13g2_fill_1 FILLER_102_16 ();
 sg13g2_decap_4 FILLER_102_47 ();
 sg13g2_decap_8 FILLER_102_56 ();
 sg13g2_decap_8 FILLER_102_63 ();
 sg13g2_fill_2 FILLER_102_70 ();
 sg13g2_fill_1 FILLER_102_72 ();
 sg13g2_decap_8 FILLER_102_98 ();
 sg13g2_decap_8 FILLER_102_105 ();
 sg13g2_fill_2 FILLER_102_112 ();
 sg13g2_decap_4 FILLER_102_134 ();
 sg13g2_fill_1 FILLER_102_138 ();
 sg13g2_decap_8 FILLER_102_147 ();
 sg13g2_decap_8 FILLER_102_154 ();
 sg13g2_decap_4 FILLER_102_161 ();
 sg13g2_fill_1 FILLER_102_165 ();
 sg13g2_decap_4 FILLER_102_178 ();
 sg13g2_fill_2 FILLER_102_182 ();
 sg13g2_decap_8 FILLER_102_191 ();
 sg13g2_decap_8 FILLER_102_198 ();
 sg13g2_decap_8 FILLER_102_205 ();
 sg13g2_fill_1 FILLER_102_212 ();
 sg13g2_fill_2 FILLER_102_234 ();
 sg13g2_fill_1 FILLER_102_236 ();
 sg13g2_decap_8 FILLER_102_253 ();
 sg13g2_decap_4 FILLER_102_260 ();
 sg13g2_fill_1 FILLER_102_264 ();
 sg13g2_fill_2 FILLER_102_269 ();
 sg13g2_decap_8 FILLER_102_277 ();
 sg13g2_decap_8 FILLER_102_284 ();
 sg13g2_fill_1 FILLER_102_291 ();
 sg13g2_decap_8 FILLER_102_309 ();
 sg13g2_decap_4 FILLER_102_316 ();
 sg13g2_decap_4 FILLER_102_328 ();
 sg13g2_fill_2 FILLER_102_332 ();
 sg13g2_decap_8 FILLER_102_339 ();
 sg13g2_decap_8 FILLER_102_346 ();
 sg13g2_decap_8 FILLER_102_353 ();
 sg13g2_decap_4 FILLER_102_360 ();
 sg13g2_fill_2 FILLER_102_364 ();
 sg13g2_decap_8 FILLER_102_371 ();
 sg13g2_fill_2 FILLER_102_378 ();
 sg13g2_decap_8 FILLER_102_395 ();
 sg13g2_decap_8 FILLER_102_406 ();
 sg13g2_decap_8 FILLER_102_413 ();
 sg13g2_decap_8 FILLER_102_420 ();
 sg13g2_decap_8 FILLER_102_427 ();
 sg13g2_fill_2 FILLER_102_434 ();
 sg13g2_fill_1 FILLER_102_436 ();
 sg13g2_decap_8 FILLER_102_447 ();
 sg13g2_decap_8 FILLER_102_454 ();
 sg13g2_decap_8 FILLER_102_461 ();
 sg13g2_decap_8 FILLER_102_468 ();
 sg13g2_decap_8 FILLER_102_475 ();
 sg13g2_decap_8 FILLER_102_482 ();
 sg13g2_decap_8 FILLER_102_489 ();
 sg13g2_decap_8 FILLER_102_496 ();
 sg13g2_decap_4 FILLER_102_503 ();
 sg13g2_fill_1 FILLER_102_507 ();
 sg13g2_fill_1 FILLER_102_513 ();
 sg13g2_decap_8 FILLER_102_527 ();
 sg13g2_decap_8 FILLER_102_534 ();
 sg13g2_fill_2 FILLER_102_541 ();
 sg13g2_fill_1 FILLER_102_543 ();
 sg13g2_decap_8 FILLER_102_564 ();
 sg13g2_decap_8 FILLER_102_571 ();
 sg13g2_decap_8 FILLER_102_578 ();
 sg13g2_fill_1 FILLER_102_585 ();
 sg13g2_fill_2 FILLER_102_611 ();
 sg13g2_fill_1 FILLER_102_613 ();
 sg13g2_decap_8 FILLER_102_648 ();
 sg13g2_decap_8 FILLER_102_655 ();
 sg13g2_decap_8 FILLER_102_662 ();
 sg13g2_decap_8 FILLER_102_669 ();
 sg13g2_decap_4 FILLER_102_676 ();
 sg13g2_fill_2 FILLER_102_680 ();
 sg13g2_fill_2 FILLER_102_728 ();
 sg13g2_decap_8 FILLER_102_734 ();
 sg13g2_decap_8 FILLER_102_741 ();
 sg13g2_decap_8 FILLER_102_748 ();
 sg13g2_fill_2 FILLER_102_755 ();
 sg13g2_fill_1 FILLER_102_757 ();
 sg13g2_decap_8 FILLER_102_761 ();
 sg13g2_fill_2 FILLER_102_768 ();
 sg13g2_fill_1 FILLER_102_770 ();
 sg13g2_decap_8 FILLER_102_783 ();
 sg13g2_decap_8 FILLER_102_790 ();
 sg13g2_decap_8 FILLER_102_797 ();
 sg13g2_decap_8 FILLER_102_804 ();
 sg13g2_fill_2 FILLER_102_811 ();
 sg13g2_decap_4 FILLER_102_817 ();
 sg13g2_decap_4 FILLER_102_835 ();
 sg13g2_fill_2 FILLER_102_839 ();
 sg13g2_decap_8 FILLER_102_867 ();
 sg13g2_decap_8 FILLER_102_874 ();
 sg13g2_decap_8 FILLER_102_881 ();
 sg13g2_decap_8 FILLER_102_888 ();
 sg13g2_decap_4 FILLER_102_895 ();
 sg13g2_fill_2 FILLER_102_899 ();
 sg13g2_decap_8 FILLER_102_904 ();
 sg13g2_decap_8 FILLER_102_911 ();
 sg13g2_fill_1 FILLER_102_918 ();
 sg13g2_decap_8 FILLER_102_936 ();
 sg13g2_decap_4 FILLER_102_943 ();
 sg13g2_fill_1 FILLER_102_947 ();
 sg13g2_decap_8 FILLER_102_974 ();
 sg13g2_decap_8 FILLER_102_981 ();
 sg13g2_decap_8 FILLER_102_988 ();
 sg13g2_decap_8 FILLER_102_995 ();
 sg13g2_decap_4 FILLER_102_1002 ();
 sg13g2_decap_4 FILLER_102_1011 ();
 sg13g2_fill_1 FILLER_102_1015 ();
 sg13g2_decap_8 FILLER_102_1028 ();
 sg13g2_decap_8 FILLER_102_1035 ();
 sg13g2_decap_8 FILLER_102_1042 ();
 sg13g2_decap_8 FILLER_102_1049 ();
 sg13g2_decap_8 FILLER_102_1056 ();
 sg13g2_decap_8 FILLER_102_1063 ();
 sg13g2_decap_8 FILLER_102_1070 ();
 sg13g2_decap_8 FILLER_102_1077 ();
 sg13g2_fill_1 FILLER_102_1084 ();
 sg13g2_decap_8 FILLER_102_1089 ();
 sg13g2_decap_8 FILLER_102_1096 ();
 sg13g2_fill_1 FILLER_102_1103 ();
 sg13g2_fill_1 FILLER_102_1108 ();
 sg13g2_decap_8 FILLER_102_1117 ();
 sg13g2_decap_8 FILLER_102_1124 ();
 sg13g2_decap_8 FILLER_102_1131 ();
 sg13g2_decap_8 FILLER_102_1138 ();
 sg13g2_decap_8 FILLER_102_1145 ();
 sg13g2_decap_8 FILLER_102_1152 ();
 sg13g2_fill_1 FILLER_102_1159 ();
 sg13g2_fill_2 FILLER_102_1186 ();
 sg13g2_fill_1 FILLER_102_1188 ();
 sg13g2_decap_8 FILLER_102_1202 ();
 sg13g2_decap_8 FILLER_102_1209 ();
 sg13g2_fill_2 FILLER_102_1216 ();
 sg13g2_fill_1 FILLER_102_1218 ();
 sg13g2_fill_2 FILLER_102_1302 ();
 sg13g2_decap_4 FILLER_102_1314 ();
 sg13g2_decap_8 FILLER_102_1323 ();
 sg13g2_decap_8 FILLER_102_1330 ();
 sg13g2_decap_8 FILLER_102_1337 ();
 sg13g2_decap_8 FILLER_102_1344 ();
 sg13g2_decap_8 FILLER_102_1351 ();
 sg13g2_decap_4 FILLER_102_1358 ();
 sg13g2_fill_2 FILLER_102_1362 ();
 sg13g2_decap_8 FILLER_102_1368 ();
 sg13g2_decap_8 FILLER_102_1375 ();
 sg13g2_decap_8 FILLER_102_1382 ();
 sg13g2_decap_8 FILLER_102_1389 ();
 sg13g2_fill_2 FILLER_102_1396 ();
 sg13g2_decap_8 FILLER_102_1420 ();
 sg13g2_decap_8 FILLER_102_1427 ();
 sg13g2_decap_8 FILLER_102_1434 ();
 sg13g2_decap_8 FILLER_102_1441 ();
 sg13g2_decap_8 FILLER_102_1448 ();
 sg13g2_decap_8 FILLER_102_1455 ();
 sg13g2_decap_8 FILLER_102_1462 ();
 sg13g2_decap_4 FILLER_102_1469 ();
 sg13g2_fill_1 FILLER_102_1473 ();
 sg13g2_decap_8 FILLER_102_1485 ();
 sg13g2_decap_8 FILLER_102_1492 ();
 sg13g2_fill_2 FILLER_102_1499 ();
 sg13g2_decap_8 FILLER_102_1521 ();
 sg13g2_fill_2 FILLER_102_1528 ();
 sg13g2_fill_1 FILLER_102_1530 ();
 sg13g2_decap_4 FILLER_102_1539 ();
 sg13g2_fill_1 FILLER_102_1543 ();
 sg13g2_decap_8 FILLER_102_1547 ();
 sg13g2_decap_8 FILLER_102_1554 ();
 sg13g2_fill_1 FILLER_102_1561 ();
 sg13g2_decap_4 FILLER_102_1570 ();
 sg13g2_decap_8 FILLER_102_1582 ();
 sg13g2_decap_4 FILLER_102_1589 ();
 sg13g2_decap_8 FILLER_102_1600 ();
 sg13g2_decap_8 FILLER_102_1607 ();
 sg13g2_fill_2 FILLER_102_1614 ();
 sg13g2_decap_8 FILLER_102_1627 ();
 sg13g2_decap_8 FILLER_102_1634 ();
 sg13g2_decap_8 FILLER_102_1641 ();
 sg13g2_decap_8 FILLER_102_1648 ();
 sg13g2_decap_8 FILLER_102_1655 ();
 sg13g2_decap_8 FILLER_102_1662 ();
 sg13g2_decap_8 FILLER_102_1669 ();
 sg13g2_decap_8 FILLER_102_1676 ();
 sg13g2_decap_8 FILLER_102_1683 ();
 sg13g2_decap_8 FILLER_102_1690 ();
 sg13g2_fill_2 FILLER_102_1697 ();
 sg13g2_fill_1 FILLER_102_1699 ();
 sg13g2_decap_8 FILLER_102_1710 ();
 sg13g2_decap_8 FILLER_102_1717 ();
 sg13g2_decap_8 FILLER_102_1724 ();
 sg13g2_fill_2 FILLER_102_1731 ();
 sg13g2_fill_2 FILLER_102_1738 ();
 sg13g2_decap_8 FILLER_102_1751 ();
 sg13g2_decap_8 FILLER_102_1758 ();
 sg13g2_fill_2 FILLER_102_1765 ();
 sg13g2_fill_1 FILLER_102_1767 ();
 sg13g2_decap_8 FILLER_103_0 ();
 sg13g2_decap_8 FILLER_103_7 ();
 sg13g2_decap_8 FILLER_103_14 ();
 sg13g2_decap_8 FILLER_103_21 ();
 sg13g2_decap_8 FILLER_103_28 ();
 sg13g2_decap_8 FILLER_103_35 ();
 sg13g2_fill_2 FILLER_103_42 ();
 sg13g2_fill_1 FILLER_103_44 ();
 sg13g2_decap_8 FILLER_103_53 ();
 sg13g2_decap_8 FILLER_103_60 ();
 sg13g2_decap_4 FILLER_103_67 ();
 sg13g2_fill_1 FILLER_103_71 ();
 sg13g2_decap_8 FILLER_103_76 ();
 sg13g2_fill_2 FILLER_103_83 ();
 sg13g2_decap_4 FILLER_103_90 ();
 sg13g2_fill_2 FILLER_103_94 ();
 sg13g2_decap_8 FILLER_103_104 ();
 sg13g2_decap_8 FILLER_103_111 ();
 sg13g2_decap_4 FILLER_103_118 ();
 sg13g2_decap_8 FILLER_103_127 ();
 sg13g2_decap_8 FILLER_103_134 ();
 sg13g2_decap_8 FILLER_103_141 ();
 sg13g2_decap_8 FILLER_103_148 ();
 sg13g2_decap_8 FILLER_103_155 ();
 sg13g2_decap_8 FILLER_103_199 ();
 sg13g2_decap_8 FILLER_103_206 ();
 sg13g2_decap_8 FILLER_103_213 ();
 sg13g2_decap_4 FILLER_103_220 ();
 sg13g2_fill_2 FILLER_103_224 ();
 sg13g2_decap_8 FILLER_103_230 ();
 sg13g2_fill_2 FILLER_103_237 ();
 sg13g2_decap_8 FILLER_103_244 ();
 sg13g2_decap_8 FILLER_103_251 ();
 sg13g2_decap_8 FILLER_103_258 ();
 sg13g2_decap_8 FILLER_103_265 ();
 sg13g2_decap_8 FILLER_103_272 ();
 sg13g2_decap_8 FILLER_103_279 ();
 sg13g2_decap_8 FILLER_103_286 ();
 sg13g2_decap_8 FILLER_103_293 ();
 sg13g2_decap_8 FILLER_103_300 ();
 sg13g2_decap_8 FILLER_103_307 ();
 sg13g2_fill_2 FILLER_103_314 ();
 sg13g2_decap_8 FILLER_103_322 ();
 sg13g2_decap_4 FILLER_103_329 ();
 sg13g2_fill_2 FILLER_103_338 ();
 sg13g2_decap_8 FILLER_103_348 ();
 sg13g2_decap_8 FILLER_103_355 ();
 sg13g2_decap_8 FILLER_103_362 ();
 sg13g2_fill_2 FILLER_103_369 ();
 sg13g2_decap_8 FILLER_103_403 ();
 sg13g2_decap_8 FILLER_103_410 ();
 sg13g2_decap_8 FILLER_103_417 ();
 sg13g2_decap_8 FILLER_103_424 ();
 sg13g2_decap_8 FILLER_103_431 ();
 sg13g2_fill_1 FILLER_103_438 ();
 sg13g2_decap_8 FILLER_103_443 ();
 sg13g2_decap_8 FILLER_103_450 ();
 sg13g2_decap_8 FILLER_103_457 ();
 sg13g2_decap_4 FILLER_103_464 ();
 sg13g2_decap_8 FILLER_103_474 ();
 sg13g2_decap_8 FILLER_103_481 ();
 sg13g2_decap_8 FILLER_103_488 ();
 sg13g2_decap_8 FILLER_103_495 ();
 sg13g2_decap_8 FILLER_103_502 ();
 sg13g2_decap_8 FILLER_103_509 ();
 sg13g2_decap_8 FILLER_103_516 ();
 sg13g2_decap_8 FILLER_103_523 ();
 sg13g2_decap_8 FILLER_103_530 ();
 sg13g2_fill_1 FILLER_103_561 ();
 sg13g2_decap_8 FILLER_103_567 ();
 sg13g2_decap_8 FILLER_103_574 ();
 sg13g2_decap_8 FILLER_103_581 ();
 sg13g2_decap_8 FILLER_103_607 ();
 sg13g2_decap_8 FILLER_103_614 ();
 sg13g2_decap_4 FILLER_103_621 ();
 sg13g2_decap_8 FILLER_103_629 ();
 sg13g2_decap_8 FILLER_103_636 ();
 sg13g2_fill_2 FILLER_103_643 ();
 sg13g2_decap_8 FILLER_103_658 ();
 sg13g2_decap_8 FILLER_103_665 ();
 sg13g2_decap_8 FILLER_103_672 ();
 sg13g2_decap_4 FILLER_103_679 ();
 sg13g2_fill_1 FILLER_103_683 ();
 sg13g2_decap_4 FILLER_103_695 ();
 sg13g2_decap_8 FILLER_103_703 ();
 sg13g2_decap_8 FILLER_103_710 ();
 sg13g2_fill_2 FILLER_103_717 ();
 sg13g2_fill_2 FILLER_103_722 ();
 sg13g2_fill_1 FILLER_103_724 ();
 sg13g2_fill_1 FILLER_103_729 ();
 sg13g2_decap_8 FILLER_103_738 ();
 sg13g2_decap_8 FILLER_103_745 ();
 sg13g2_decap_4 FILLER_103_752 ();
 sg13g2_fill_2 FILLER_103_756 ();
 sg13g2_decap_8 FILLER_103_794 ();
 sg13g2_fill_2 FILLER_103_801 ();
 sg13g2_decap_8 FILLER_103_806 ();
 sg13g2_decap_8 FILLER_103_813 ();
 sg13g2_decap_8 FILLER_103_820 ();
 sg13g2_decap_8 FILLER_103_827 ();
 sg13g2_decap_4 FILLER_103_859 ();
 sg13g2_fill_2 FILLER_103_863 ();
 sg13g2_decap_8 FILLER_103_873 ();
 sg13g2_decap_8 FILLER_103_880 ();
 sg13g2_decap_8 FILLER_103_887 ();
 sg13g2_decap_4 FILLER_103_894 ();
 sg13g2_decap_8 FILLER_103_917 ();
 sg13g2_decap_8 FILLER_103_924 ();
 sg13g2_decap_8 FILLER_103_931 ();
 sg13g2_decap_8 FILLER_103_938 ();
 sg13g2_decap_8 FILLER_103_945 ();
 sg13g2_decap_4 FILLER_103_952 ();
 sg13g2_fill_2 FILLER_103_956 ();
 sg13g2_decap_8 FILLER_103_962 ();
 sg13g2_decap_8 FILLER_103_969 ();
 sg13g2_decap_4 FILLER_103_976 ();
 sg13g2_fill_2 FILLER_103_980 ();
 sg13g2_decap_8 FILLER_103_987 ();
 sg13g2_decap_8 FILLER_103_994 ();
 sg13g2_decap_8 FILLER_103_1001 ();
 sg13g2_fill_2 FILLER_103_1008 ();
 sg13g2_decap_8 FILLER_103_1015 ();
 sg13g2_decap_8 FILLER_103_1027 ();
 sg13g2_decap_8 FILLER_103_1034 ();
 sg13g2_decap_8 FILLER_103_1041 ();
 sg13g2_decap_8 FILLER_103_1048 ();
 sg13g2_decap_8 FILLER_103_1055 ();
 sg13g2_decap_8 FILLER_103_1062 ();
 sg13g2_decap_8 FILLER_103_1069 ();
 sg13g2_decap_8 FILLER_103_1076 ();
 sg13g2_decap_8 FILLER_103_1083 ();
 sg13g2_decap_8 FILLER_103_1134 ();
 sg13g2_fill_2 FILLER_103_1141 ();
 sg13g2_fill_1 FILLER_103_1143 ();
 sg13g2_decap_8 FILLER_103_1148 ();
 sg13g2_fill_2 FILLER_103_1155 ();
 sg13g2_fill_1 FILLER_103_1157 ();
 sg13g2_decap_8 FILLER_103_1163 ();
 sg13g2_fill_1 FILLER_103_1170 ();
 sg13g2_decap_8 FILLER_103_1175 ();
 sg13g2_decap_8 FILLER_103_1182 ();
 sg13g2_fill_2 FILLER_103_1189 ();
 sg13g2_fill_1 FILLER_103_1191 ();
 sg13g2_decap_8 FILLER_103_1207 ();
 sg13g2_decap_8 FILLER_103_1214 ();
 sg13g2_decap_8 FILLER_103_1225 ();
 sg13g2_fill_2 FILLER_103_1232 ();
 sg13g2_fill_1 FILLER_103_1234 ();
 sg13g2_decap_8 FILLER_103_1240 ();
 sg13g2_decap_8 FILLER_103_1247 ();
 sg13g2_decap_8 FILLER_103_1254 ();
 sg13g2_decap_8 FILLER_103_1261 ();
 sg13g2_decap_8 FILLER_103_1268 ();
 sg13g2_decap_8 FILLER_103_1275 ();
 sg13g2_decap_8 FILLER_103_1282 ();
 sg13g2_fill_1 FILLER_103_1289 ();
 sg13g2_decap_8 FILLER_103_1305 ();
 sg13g2_decap_8 FILLER_103_1312 ();
 sg13g2_decap_8 FILLER_103_1319 ();
 sg13g2_decap_8 FILLER_103_1326 ();
 sg13g2_decap_8 FILLER_103_1337 ();
 sg13g2_decap_8 FILLER_103_1344 ();
 sg13g2_decap_8 FILLER_103_1351 ();
 sg13g2_decap_4 FILLER_103_1358 ();
 sg13g2_decap_8 FILLER_103_1369 ();
 sg13g2_decap_8 FILLER_103_1376 ();
 sg13g2_fill_2 FILLER_103_1383 ();
 sg13g2_decap_8 FILLER_103_1397 ();
 sg13g2_decap_8 FILLER_103_1404 ();
 sg13g2_fill_1 FILLER_103_1411 ();
 sg13g2_decap_8 FILLER_103_1420 ();
 sg13g2_decap_4 FILLER_103_1427 ();
 sg13g2_fill_1 FILLER_103_1431 ();
 sg13g2_decap_8 FILLER_103_1440 ();
 sg13g2_decap_8 FILLER_103_1447 ();
 sg13g2_decap_4 FILLER_103_1454 ();
 sg13g2_decap_8 FILLER_103_1462 ();
 sg13g2_fill_1 FILLER_103_1469 ();
 sg13g2_decap_8 FILLER_103_1475 ();
 sg13g2_decap_8 FILLER_103_1482 ();
 sg13g2_decap_4 FILLER_103_1489 ();
 sg13g2_fill_2 FILLER_103_1493 ();
 sg13g2_fill_2 FILLER_103_1503 ();
 sg13g2_fill_1 FILLER_103_1505 ();
 sg13g2_decap_8 FILLER_103_1514 ();
 sg13g2_decap_8 FILLER_103_1521 ();
 sg13g2_decap_8 FILLER_103_1528 ();
 sg13g2_fill_2 FILLER_103_1535 ();
 sg13g2_fill_1 FILLER_103_1537 ();
 sg13g2_fill_2 FILLER_103_1549 ();
 sg13g2_decap_8 FILLER_103_1559 ();
 sg13g2_decap_4 FILLER_103_1566 ();
 sg13g2_fill_1 FILLER_103_1570 ();
 sg13g2_decap_8 FILLER_103_1604 ();
 sg13g2_decap_4 FILLER_103_1611 ();
 sg13g2_fill_1 FILLER_103_1615 ();
 sg13g2_decap_8 FILLER_103_1633 ();
 sg13g2_decap_8 FILLER_103_1640 ();
 sg13g2_decap_8 FILLER_103_1647 ();
 sg13g2_fill_2 FILLER_103_1670 ();
 sg13g2_decap_8 FILLER_103_1676 ();
 sg13g2_decap_8 FILLER_103_1683 ();
 sg13g2_decap_8 FILLER_103_1690 ();
 sg13g2_decap_8 FILLER_103_1697 ();
 sg13g2_decap_8 FILLER_103_1704 ();
 sg13g2_decap_8 FILLER_103_1711 ();
 sg13g2_fill_2 FILLER_103_1726 ();
 sg13g2_decap_8 FILLER_103_1736 ();
 sg13g2_decap_8 FILLER_103_1743 ();
 sg13g2_decap_8 FILLER_103_1750 ();
 sg13g2_decap_8 FILLER_103_1757 ();
 sg13g2_decap_4 FILLER_103_1764 ();
 sg13g2_decap_8 FILLER_104_0 ();
 sg13g2_decap_8 FILLER_104_7 ();
 sg13g2_decap_8 FILLER_104_14 ();
 sg13g2_decap_8 FILLER_104_21 ();
 sg13g2_decap_8 FILLER_104_28 ();
 sg13g2_decap_8 FILLER_104_35 ();
 sg13g2_decap_8 FILLER_104_42 ();
 sg13g2_decap_8 FILLER_104_49 ();
 sg13g2_decap_8 FILLER_104_56 ();
 sg13g2_decap_8 FILLER_104_63 ();
 sg13g2_decap_8 FILLER_104_70 ();
 sg13g2_decap_8 FILLER_104_77 ();
 sg13g2_decap_8 FILLER_104_84 ();
 sg13g2_decap_8 FILLER_104_91 ();
 sg13g2_decap_8 FILLER_104_98 ();
 sg13g2_decap_8 FILLER_104_105 ();
 sg13g2_decap_8 FILLER_104_112 ();
 sg13g2_decap_8 FILLER_104_119 ();
 sg13g2_decap_8 FILLER_104_126 ();
 sg13g2_decap_8 FILLER_104_133 ();
 sg13g2_decap_8 FILLER_104_140 ();
 sg13g2_decap_8 FILLER_104_147 ();
 sg13g2_decap_8 FILLER_104_158 ();
 sg13g2_decap_8 FILLER_104_165 ();
 sg13g2_decap_8 FILLER_104_172 ();
 sg13g2_decap_4 FILLER_104_179 ();
 sg13g2_fill_2 FILLER_104_183 ();
 sg13g2_fill_1 FILLER_104_197 ();
 sg13g2_decap_8 FILLER_104_204 ();
 sg13g2_fill_2 FILLER_104_211 ();
 sg13g2_fill_1 FILLER_104_213 ();
 sg13g2_decap_8 FILLER_104_222 ();
 sg13g2_decap_4 FILLER_104_229 ();
 sg13g2_fill_2 FILLER_104_233 ();
 sg13g2_fill_1 FILLER_104_258 ();
 sg13g2_decap_8 FILLER_104_264 ();
 sg13g2_fill_2 FILLER_104_271 ();
 sg13g2_decap_8 FILLER_104_277 ();
 sg13g2_decap_8 FILLER_104_284 ();
 sg13g2_decap_8 FILLER_104_291 ();
 sg13g2_decap_8 FILLER_104_298 ();
 sg13g2_decap_8 FILLER_104_305 ();
 sg13g2_decap_8 FILLER_104_312 ();
 sg13g2_fill_2 FILLER_104_319 ();
 sg13g2_decap_8 FILLER_104_331 ();
 sg13g2_decap_8 FILLER_104_338 ();
 sg13g2_decap_8 FILLER_104_345 ();
 sg13g2_decap_8 FILLER_104_352 ();
 sg13g2_decap_8 FILLER_104_359 ();
 sg13g2_decap_8 FILLER_104_366 ();
 sg13g2_decap_4 FILLER_104_373 ();
 sg13g2_fill_2 FILLER_104_377 ();
 sg13g2_decap_8 FILLER_104_387 ();
 sg13g2_fill_2 FILLER_104_394 ();
 sg13g2_fill_1 FILLER_104_396 ();
 sg13g2_decap_8 FILLER_104_402 ();
 sg13g2_decap_8 FILLER_104_409 ();
 sg13g2_decap_8 FILLER_104_416 ();
 sg13g2_fill_1 FILLER_104_423 ();
 sg13g2_decap_8 FILLER_104_436 ();
 sg13g2_decap_4 FILLER_104_458 ();
 sg13g2_fill_1 FILLER_104_462 ();
 sg13g2_decap_8 FILLER_104_482 ();
 sg13g2_decap_8 FILLER_104_489 ();
 sg13g2_decap_4 FILLER_104_496 ();
 sg13g2_fill_2 FILLER_104_500 ();
 sg13g2_decap_8 FILLER_104_507 ();
 sg13g2_decap_8 FILLER_104_514 ();
 sg13g2_decap_8 FILLER_104_521 ();
 sg13g2_decap_8 FILLER_104_528 ();
 sg13g2_decap_8 FILLER_104_535 ();
 sg13g2_decap_8 FILLER_104_542 ();
 sg13g2_decap_4 FILLER_104_549 ();
 sg13g2_decap_8 FILLER_104_557 ();
 sg13g2_decap_8 FILLER_104_564 ();
 sg13g2_decap_8 FILLER_104_571 ();
 sg13g2_decap_8 FILLER_104_578 ();
 sg13g2_decap_8 FILLER_104_585 ();
 sg13g2_fill_2 FILLER_104_592 ();
 sg13g2_decap_8 FILLER_104_605 ();
 sg13g2_decap_8 FILLER_104_612 ();
 sg13g2_decap_8 FILLER_104_619 ();
 sg13g2_decap_8 FILLER_104_626 ();
 sg13g2_decap_8 FILLER_104_633 ();
 sg13g2_decap_8 FILLER_104_640 ();
 sg13g2_decap_8 FILLER_104_647 ();
 sg13g2_decap_8 FILLER_104_654 ();
 sg13g2_decap_8 FILLER_104_661 ();
 sg13g2_decap_8 FILLER_104_668 ();
 sg13g2_decap_8 FILLER_104_675 ();
 sg13g2_decap_8 FILLER_104_682 ();
 sg13g2_decap_8 FILLER_104_689 ();
 sg13g2_decap_8 FILLER_104_696 ();
 sg13g2_decap_8 FILLER_104_703 ();
 sg13g2_decap_8 FILLER_104_710 ();
 sg13g2_decap_8 FILLER_104_717 ();
 sg13g2_decap_8 FILLER_104_724 ();
 sg13g2_decap_8 FILLER_104_731 ();
 sg13g2_decap_8 FILLER_104_738 ();
 sg13g2_decap_8 FILLER_104_745 ();
 sg13g2_decap_4 FILLER_104_752 ();
 sg13g2_fill_2 FILLER_104_756 ();
 sg13g2_decap_8 FILLER_104_768 ();
 sg13g2_decap_8 FILLER_104_775 ();
 sg13g2_decap_8 FILLER_104_782 ();
 sg13g2_decap_8 FILLER_104_789 ();
 sg13g2_decap_4 FILLER_104_796 ();
 sg13g2_decap_8 FILLER_104_809 ();
 sg13g2_fill_1 FILLER_104_816 ();
 sg13g2_decap_8 FILLER_104_822 ();
 sg13g2_decap_8 FILLER_104_829 ();
 sg13g2_decap_8 FILLER_104_836 ();
 sg13g2_decap_4 FILLER_104_843 ();
 sg13g2_decap_8 FILLER_104_850 ();
 sg13g2_decap_8 FILLER_104_857 ();
 sg13g2_decap_8 FILLER_104_864 ();
 sg13g2_decap_8 FILLER_104_871 ();
 sg13g2_decap_8 FILLER_104_878 ();
 sg13g2_decap_8 FILLER_104_885 ();
 sg13g2_decap_8 FILLER_104_892 ();
 sg13g2_fill_2 FILLER_104_899 ();
 sg13g2_decap_8 FILLER_104_904 ();
 sg13g2_decap_8 FILLER_104_911 ();
 sg13g2_decap_8 FILLER_104_918 ();
 sg13g2_decap_8 FILLER_104_925 ();
 sg13g2_decap_8 FILLER_104_932 ();
 sg13g2_decap_8 FILLER_104_939 ();
 sg13g2_decap_8 FILLER_104_946 ();
 sg13g2_decap_8 FILLER_104_953 ();
 sg13g2_decap_8 FILLER_104_960 ();
 sg13g2_decap_8 FILLER_104_967 ();
 sg13g2_decap_8 FILLER_104_974 ();
 sg13g2_decap_4 FILLER_104_981 ();
 sg13g2_fill_2 FILLER_104_990 ();
 sg13g2_fill_1 FILLER_104_992 ();
 sg13g2_decap_8 FILLER_104_997 ();
 sg13g2_fill_2 FILLER_104_1004 ();
 sg13g2_fill_1 FILLER_104_1006 ();
 sg13g2_fill_2 FILLER_104_1015 ();
 sg13g2_fill_2 FILLER_104_1025 ();
 sg13g2_fill_1 FILLER_104_1027 ();
 sg13g2_fill_2 FILLER_104_1054 ();
 sg13g2_fill_1 FILLER_104_1056 ();
 sg13g2_decap_8 FILLER_104_1083 ();
 sg13g2_decap_8 FILLER_104_1090 ();
 sg13g2_decap_8 FILLER_104_1100 ();
 sg13g2_fill_1 FILLER_104_1107 ();
 sg13g2_fill_1 FILLER_104_1125 ();
 sg13g2_decap_8 FILLER_104_1160 ();
 sg13g2_decap_8 FILLER_104_1167 ();
 sg13g2_decap_8 FILLER_104_1174 ();
 sg13g2_decap_8 FILLER_104_1181 ();
 sg13g2_decap_8 FILLER_104_1188 ();
 sg13g2_decap_8 FILLER_104_1195 ();
 sg13g2_decap_8 FILLER_104_1202 ();
 sg13g2_decap_8 FILLER_104_1209 ();
 sg13g2_decap_8 FILLER_104_1216 ();
 sg13g2_decap_8 FILLER_104_1223 ();
 sg13g2_decap_4 FILLER_104_1230 ();
 sg13g2_fill_2 FILLER_104_1234 ();
 sg13g2_decap_8 FILLER_104_1244 ();
 sg13g2_decap_8 FILLER_104_1251 ();
 sg13g2_decap_8 FILLER_104_1258 ();
 sg13g2_decap_8 FILLER_104_1265 ();
 sg13g2_decap_8 FILLER_104_1272 ();
 sg13g2_decap_4 FILLER_104_1279 ();
 sg13g2_decap_8 FILLER_104_1291 ();
 sg13g2_decap_8 FILLER_104_1298 ();
 sg13g2_decap_8 FILLER_104_1305 ();
 sg13g2_decap_8 FILLER_104_1312 ();
 sg13g2_fill_2 FILLER_104_1319 ();
 sg13g2_fill_1 FILLER_104_1321 ();
 sg13g2_decap_8 FILLER_104_1348 ();
 sg13g2_fill_2 FILLER_104_1355 ();
 sg13g2_fill_1 FILLER_104_1357 ();
 sg13g2_decap_4 FILLER_104_1362 ();
 sg13g2_decap_8 FILLER_104_1382 ();
 sg13g2_decap_8 FILLER_104_1389 ();
 sg13g2_fill_1 FILLER_104_1396 ();
 sg13g2_decap_8 FILLER_104_1425 ();
 sg13g2_decap_8 FILLER_104_1432 ();
 sg13g2_decap_8 FILLER_104_1439 ();
 sg13g2_decap_4 FILLER_104_1446 ();
 sg13g2_fill_2 FILLER_104_1450 ();
 sg13g2_fill_2 FILLER_104_1494 ();
 sg13g2_fill_1 FILLER_104_1496 ();
 sg13g2_decap_8 FILLER_104_1513 ();
 sg13g2_decap_8 FILLER_104_1520 ();
 sg13g2_decap_8 FILLER_104_1527 ();
 sg13g2_decap_4 FILLER_104_1534 ();
 sg13g2_decap_8 FILLER_104_1562 ();
 sg13g2_decap_4 FILLER_104_1569 ();
 sg13g2_fill_2 FILLER_104_1573 ();
 sg13g2_decap_8 FILLER_104_1583 ();
 sg13g2_decap_8 FILLER_104_1590 ();
 sg13g2_decap_8 FILLER_104_1597 ();
 sg13g2_decap_8 FILLER_104_1604 ();
 sg13g2_decap_8 FILLER_104_1611 ();
 sg13g2_decap_8 FILLER_104_1618 ();
 sg13g2_decap_8 FILLER_104_1625 ();
 sg13g2_decap_8 FILLER_104_1632 ();
 sg13g2_decap_4 FILLER_104_1639 ();
 sg13g2_fill_2 FILLER_104_1643 ();
 sg13g2_fill_1 FILLER_104_1655 ();
 sg13g2_fill_1 FILLER_104_1668 ();
 sg13g2_decap_8 FILLER_104_1686 ();
 sg13g2_decap_8 FILLER_104_1693 ();
 sg13g2_decap_8 FILLER_104_1700 ();
 sg13g2_fill_2 FILLER_104_1707 ();
 sg13g2_fill_2 FILLER_104_1719 ();
 sg13g2_fill_1 FILLER_104_1721 ();
 sg13g2_decap_8 FILLER_104_1730 ();
 sg13g2_decap_8 FILLER_104_1737 ();
 sg13g2_decap_8 FILLER_104_1744 ();
 sg13g2_decap_8 FILLER_104_1751 ();
 sg13g2_decap_8 FILLER_104_1758 ();
 sg13g2_fill_2 FILLER_104_1765 ();
 sg13g2_fill_1 FILLER_104_1767 ();
 sg13g2_decap_8 FILLER_105_0 ();
 sg13g2_decap_8 FILLER_105_7 ();
 sg13g2_decap_8 FILLER_105_14 ();
 sg13g2_decap_8 FILLER_105_21 ();
 sg13g2_decap_8 FILLER_105_28 ();
 sg13g2_decap_8 FILLER_105_35 ();
 sg13g2_decap_8 FILLER_105_42 ();
 sg13g2_decap_8 FILLER_105_49 ();
 sg13g2_decap_8 FILLER_105_56 ();
 sg13g2_decap_8 FILLER_105_63 ();
 sg13g2_decap_8 FILLER_105_70 ();
 sg13g2_decap_8 FILLER_105_77 ();
 sg13g2_decap_8 FILLER_105_84 ();
 sg13g2_decap_8 FILLER_105_91 ();
 sg13g2_decap_8 FILLER_105_98 ();
 sg13g2_decap_8 FILLER_105_105 ();
 sg13g2_decap_8 FILLER_105_112 ();
 sg13g2_decap_8 FILLER_105_119 ();
 sg13g2_decap_8 FILLER_105_126 ();
 sg13g2_decap_8 FILLER_105_133 ();
 sg13g2_decap_8 FILLER_105_140 ();
 sg13g2_fill_2 FILLER_105_147 ();
 sg13g2_fill_1 FILLER_105_149 ();
 sg13g2_decap_8 FILLER_105_154 ();
 sg13g2_decap_8 FILLER_105_161 ();
 sg13g2_decap_8 FILLER_105_168 ();
 sg13g2_decap_8 FILLER_105_175 ();
 sg13g2_decap_8 FILLER_105_182 ();
 sg13g2_fill_1 FILLER_105_197 ();
 sg13g2_decap_8 FILLER_105_203 ();
 sg13g2_decap_8 FILLER_105_210 ();
 sg13g2_decap_8 FILLER_105_217 ();
 sg13g2_decap_8 FILLER_105_224 ();
 sg13g2_decap_8 FILLER_105_231 ();
 sg13g2_decap_8 FILLER_105_238 ();
 sg13g2_decap_4 FILLER_105_245 ();
 sg13g2_fill_2 FILLER_105_257 ();
 sg13g2_fill_1 FILLER_105_259 ();
 sg13g2_decap_8 FILLER_105_288 ();
 sg13g2_decap_8 FILLER_105_295 ();
 sg13g2_decap_8 FILLER_105_302 ();
 sg13g2_decap_4 FILLER_105_309 ();
 sg13g2_decap_8 FILLER_105_334 ();
 sg13g2_decap_8 FILLER_105_341 ();
 sg13g2_decap_4 FILLER_105_348 ();
 sg13g2_decap_8 FILLER_105_357 ();
 sg13g2_decap_8 FILLER_105_364 ();
 sg13g2_decap_8 FILLER_105_371 ();
 sg13g2_decap_8 FILLER_105_378 ();
 sg13g2_decap_8 FILLER_105_385 ();
 sg13g2_decap_8 FILLER_105_392 ();
 sg13g2_decap_8 FILLER_105_399 ();
 sg13g2_decap_8 FILLER_105_406 ();
 sg13g2_decap_8 FILLER_105_413 ();
 sg13g2_decap_8 FILLER_105_420 ();
 sg13g2_decap_4 FILLER_105_427 ();
 sg13g2_fill_1 FILLER_105_431 ();
 sg13g2_decap_8 FILLER_105_451 ();
 sg13g2_fill_2 FILLER_105_458 ();
 sg13g2_fill_1 FILLER_105_460 ();
 sg13g2_decap_8 FILLER_105_473 ();
 sg13g2_decap_8 FILLER_105_480 ();
 sg13g2_decap_4 FILLER_105_487 ();
 sg13g2_fill_1 FILLER_105_491 ();
 sg13g2_decap_8 FILLER_105_505 ();
 sg13g2_decap_4 FILLER_105_512 ();
 sg13g2_fill_2 FILLER_105_522 ();
 sg13g2_decap_8 FILLER_105_532 ();
 sg13g2_decap_8 FILLER_105_539 ();
 sg13g2_decap_8 FILLER_105_546 ();
 sg13g2_decap_8 FILLER_105_553 ();
 sg13g2_fill_2 FILLER_105_560 ();
 sg13g2_decap_8 FILLER_105_570 ();
 sg13g2_decap_8 FILLER_105_577 ();
 sg13g2_fill_2 FILLER_105_584 ();
 sg13g2_decap_8 FILLER_105_599 ();
 sg13g2_decap_8 FILLER_105_606 ();
 sg13g2_decap_8 FILLER_105_613 ();
 sg13g2_decap_8 FILLER_105_633 ();
 sg13g2_fill_2 FILLER_105_640 ();
 sg13g2_fill_1 FILLER_105_642 ();
 sg13g2_decap_8 FILLER_105_651 ();
 sg13g2_fill_2 FILLER_105_658 ();
 sg13g2_decap_8 FILLER_105_668 ();
 sg13g2_decap_8 FILLER_105_675 ();
 sg13g2_decap_8 FILLER_105_682 ();
 sg13g2_decap_8 FILLER_105_689 ();
 sg13g2_decap_8 FILLER_105_696 ();
 sg13g2_decap_4 FILLER_105_703 ();
 sg13g2_fill_2 FILLER_105_707 ();
 sg13g2_decap_8 FILLER_105_724 ();
 sg13g2_decap_8 FILLER_105_731 ();
 sg13g2_decap_8 FILLER_105_738 ();
 sg13g2_decap_8 FILLER_105_745 ();
 sg13g2_decap_8 FILLER_105_752 ();
 sg13g2_fill_2 FILLER_105_759 ();
 sg13g2_fill_1 FILLER_105_761 ();
 sg13g2_decap_4 FILLER_105_779 ();
 sg13g2_fill_2 FILLER_105_783 ();
 sg13g2_decap_4 FILLER_105_798 ();
 sg13g2_fill_1 FILLER_105_802 ();
 sg13g2_decap_4 FILLER_105_806 ();
 sg13g2_fill_1 FILLER_105_810 ();
 sg13g2_decap_8 FILLER_105_824 ();
 sg13g2_decap_8 FILLER_105_831 ();
 sg13g2_decap_8 FILLER_105_838 ();
 sg13g2_decap_8 FILLER_105_845 ();
 sg13g2_decap_8 FILLER_105_852 ();
 sg13g2_decap_8 FILLER_105_859 ();
 sg13g2_decap_8 FILLER_105_866 ();
 sg13g2_decap_8 FILLER_105_873 ();
 sg13g2_decap_8 FILLER_105_880 ();
 sg13g2_decap_8 FILLER_105_887 ();
 sg13g2_fill_1 FILLER_105_894 ();
 sg13g2_fill_2 FILLER_105_934 ();
 sg13g2_decap_8 FILLER_105_949 ();
 sg13g2_fill_1 FILLER_105_956 ();
 sg13g2_decap_8 FILLER_105_965 ();
 sg13g2_fill_2 FILLER_105_972 ();
 sg13g2_fill_1 FILLER_105_974 ();
 sg13g2_decap_4 FILLER_105_1014 ();
 sg13g2_fill_1 FILLER_105_1018 ();
 sg13g2_decap_8 FILLER_105_1023 ();
 sg13g2_decap_8 FILLER_105_1030 ();
 sg13g2_fill_2 FILLER_105_1037 ();
 sg13g2_decap_8 FILLER_105_1043 ();
 sg13g2_decap_8 FILLER_105_1050 ();
 sg13g2_decap_8 FILLER_105_1057 ();
 sg13g2_decap_8 FILLER_105_1064 ();
 sg13g2_decap_8 FILLER_105_1071 ();
 sg13g2_decap_8 FILLER_105_1078 ();
 sg13g2_decap_8 FILLER_105_1085 ();
 sg13g2_fill_2 FILLER_105_1092 ();
 sg13g2_decap_8 FILLER_105_1105 ();
 sg13g2_decap_8 FILLER_105_1112 ();
 sg13g2_fill_2 FILLER_105_1119 ();
 sg13g2_fill_1 FILLER_105_1121 ();
 sg13g2_decap_8 FILLER_105_1126 ();
 sg13g2_fill_2 FILLER_105_1133 ();
 sg13g2_fill_1 FILLER_105_1135 ();
 sg13g2_fill_2 FILLER_105_1140 ();
 sg13g2_fill_1 FILLER_105_1142 ();
 sg13g2_decap_8 FILLER_105_1161 ();
 sg13g2_fill_2 FILLER_105_1168 ();
 sg13g2_fill_1 FILLER_105_1196 ();
 sg13g2_decap_8 FILLER_105_1206 ();
 sg13g2_decap_8 FILLER_105_1213 ();
 sg13g2_decap_8 FILLER_105_1220 ();
 sg13g2_decap_8 FILLER_105_1227 ();
 sg13g2_decap_8 FILLER_105_1234 ();
 sg13g2_decap_8 FILLER_105_1241 ();
 sg13g2_decap_8 FILLER_105_1248 ();
 sg13g2_fill_2 FILLER_105_1255 ();
 sg13g2_decap_8 FILLER_105_1261 ();
 sg13g2_decap_8 FILLER_105_1268 ();
 sg13g2_decap_8 FILLER_105_1275 ();
 sg13g2_decap_8 FILLER_105_1282 ();
 sg13g2_decap_4 FILLER_105_1289 ();
 sg13g2_fill_1 FILLER_105_1293 ();
 sg13g2_decap_8 FILLER_105_1302 ();
 sg13g2_decap_8 FILLER_105_1309 ();
 sg13g2_decap_8 FILLER_105_1316 ();
 sg13g2_decap_4 FILLER_105_1323 ();
 sg13g2_decap_8 FILLER_105_1340 ();
 sg13g2_decap_8 FILLER_105_1347 ();
 sg13g2_decap_8 FILLER_105_1354 ();
 sg13g2_decap_8 FILLER_105_1361 ();
 sg13g2_decap_8 FILLER_105_1368 ();
 sg13g2_decap_8 FILLER_105_1375 ();
 sg13g2_decap_8 FILLER_105_1382 ();
 sg13g2_fill_2 FILLER_105_1389 ();
 sg13g2_decap_8 FILLER_105_1399 ();
 sg13g2_decap_4 FILLER_105_1406 ();
 sg13g2_fill_1 FILLER_105_1410 ();
 sg13g2_decap_8 FILLER_105_1420 ();
 sg13g2_decap_8 FILLER_105_1435 ();
 sg13g2_decap_8 FILLER_105_1442 ();
 sg13g2_fill_1 FILLER_105_1449 ();
 sg13g2_decap_8 FILLER_105_1474 ();
 sg13g2_decap_8 FILLER_105_1481 ();
 sg13g2_decap_8 FILLER_105_1488 ();
 sg13g2_decap_8 FILLER_105_1495 ();
 sg13g2_decap_8 FILLER_105_1502 ();
 sg13g2_decap_8 FILLER_105_1509 ();
 sg13g2_decap_8 FILLER_105_1516 ();
 sg13g2_decap_8 FILLER_105_1523 ();
 sg13g2_fill_2 FILLER_105_1530 ();
 sg13g2_decap_8 FILLER_105_1557 ();
 sg13g2_decap_8 FILLER_105_1564 ();
 sg13g2_decap_8 FILLER_105_1571 ();
 sg13g2_decap_8 FILLER_105_1578 ();
 sg13g2_decap_8 FILLER_105_1585 ();
 sg13g2_decap_8 FILLER_105_1592 ();
 sg13g2_decap_8 FILLER_105_1599 ();
 sg13g2_decap_8 FILLER_105_1606 ();
 sg13g2_decap_8 FILLER_105_1613 ();
 sg13g2_decap_8 FILLER_105_1620 ();
 sg13g2_decap_4 FILLER_105_1631 ();
 sg13g2_decap_8 FILLER_105_1643 ();
 sg13g2_decap_8 FILLER_105_1650 ();
 sg13g2_fill_2 FILLER_105_1657 ();
 sg13g2_fill_1 FILLER_105_1659 ();
 sg13g2_fill_2 FILLER_105_1674 ();
 sg13g2_decap_8 FILLER_105_1690 ();
 sg13g2_decap_8 FILLER_105_1697 ();
 sg13g2_decap_8 FILLER_105_1704 ();
 sg13g2_fill_1 FILLER_105_1711 ();
 sg13g2_fill_2 FILLER_105_1720 ();
 sg13g2_fill_1 FILLER_105_1722 ();
 sg13g2_decap_8 FILLER_105_1731 ();
 sg13g2_decap_8 FILLER_105_1738 ();
 sg13g2_decap_8 FILLER_105_1745 ();
 sg13g2_decap_8 FILLER_105_1752 ();
 sg13g2_decap_8 FILLER_105_1759 ();
 sg13g2_fill_2 FILLER_105_1766 ();
 sg13g2_decap_8 FILLER_106_0 ();
 sg13g2_decap_4 FILLER_106_7 ();
 sg13g2_decap_4 FILLER_106_37 ();
 sg13g2_decap_4 FILLER_106_54 ();
 sg13g2_fill_1 FILLER_106_58 ();
 sg13g2_decap_8 FILLER_106_72 ();
 sg13g2_decap_8 FILLER_106_79 ();
 sg13g2_decap_8 FILLER_106_86 ();
 sg13g2_decap_8 FILLER_106_93 ();
 sg13g2_fill_2 FILLER_106_100 ();
 sg13g2_fill_1 FILLER_106_102 ();
 sg13g2_decap_8 FILLER_106_113 ();
 sg13g2_decap_8 FILLER_106_120 ();
 sg13g2_decap_8 FILLER_106_127 ();
 sg13g2_fill_2 FILLER_106_134 ();
 sg13g2_fill_1 FILLER_106_136 ();
 sg13g2_fill_2 FILLER_106_142 ();
 sg13g2_decap_8 FILLER_106_160 ();
 sg13g2_decap_4 FILLER_106_167 ();
 sg13g2_fill_1 FILLER_106_171 ();
 sg13g2_decap_8 FILLER_106_180 ();
 sg13g2_decap_8 FILLER_106_187 ();
 sg13g2_fill_1 FILLER_106_194 ();
 sg13g2_decap_8 FILLER_106_203 ();
 sg13g2_decap_8 FILLER_106_210 ();
 sg13g2_decap_8 FILLER_106_217 ();
 sg13g2_decap_8 FILLER_106_224 ();
 sg13g2_decap_8 FILLER_106_231 ();
 sg13g2_decap_8 FILLER_106_238 ();
 sg13g2_decap_8 FILLER_106_245 ();
 sg13g2_decap_8 FILLER_106_257 ();
 sg13g2_decap_8 FILLER_106_264 ();
 sg13g2_fill_2 FILLER_106_271 ();
 sg13g2_fill_1 FILLER_106_273 ();
 sg13g2_decap_8 FILLER_106_299 ();
 sg13g2_decap_8 FILLER_106_306 ();
 sg13g2_fill_2 FILLER_106_313 ();
 sg13g2_fill_1 FILLER_106_315 ();
 sg13g2_fill_1 FILLER_106_334 ();
 sg13g2_decap_8 FILLER_106_343 ();
 sg13g2_decap_8 FILLER_106_350 ();
 sg13g2_decap_8 FILLER_106_357 ();
 sg13g2_decap_8 FILLER_106_364 ();
 sg13g2_decap_8 FILLER_106_371 ();
 sg13g2_decap_8 FILLER_106_378 ();
 sg13g2_decap_8 FILLER_106_385 ();
 sg13g2_decap_8 FILLER_106_392 ();
 sg13g2_fill_1 FILLER_106_399 ();
 sg13g2_decap_4 FILLER_106_411 ();
 sg13g2_fill_1 FILLER_106_415 ();
 sg13g2_decap_8 FILLER_106_426 ();
 sg13g2_fill_2 FILLER_106_433 ();
 sg13g2_fill_2 FILLER_106_450 ();
 sg13g2_fill_1 FILLER_106_452 ();
 sg13g2_fill_2 FILLER_106_463 ();
 sg13g2_fill_1 FILLER_106_465 ();
 sg13g2_decap_8 FILLER_106_479 ();
 sg13g2_decap_8 FILLER_106_486 ();
 sg13g2_decap_8 FILLER_106_493 ();
 sg13g2_decap_4 FILLER_106_500 ();
 sg13g2_fill_2 FILLER_106_504 ();
 sg13g2_decap_4 FILLER_106_536 ();
 sg13g2_fill_1 FILLER_106_540 ();
 sg13g2_decap_8 FILLER_106_545 ();
 sg13g2_decap_8 FILLER_106_552 ();
 sg13g2_decap_8 FILLER_106_559 ();
 sg13g2_decap_8 FILLER_106_566 ();
 sg13g2_decap_8 FILLER_106_573 ();
 sg13g2_decap_8 FILLER_106_580 ();
 sg13g2_fill_2 FILLER_106_587 ();
 sg13g2_fill_1 FILLER_106_589 ();
 sg13g2_decap_8 FILLER_106_603 ();
 sg13g2_fill_1 FILLER_106_610 ();
 sg13g2_decap_8 FILLER_106_619 ();
 sg13g2_decap_8 FILLER_106_626 ();
 sg13g2_decap_8 FILLER_106_633 ();
 sg13g2_decap_8 FILLER_106_640 ();
 sg13g2_decap_8 FILLER_106_647 ();
 sg13g2_decap_8 FILLER_106_654 ();
 sg13g2_fill_2 FILLER_106_665 ();
 sg13g2_fill_1 FILLER_106_667 ();
 sg13g2_decap_8 FILLER_106_677 ();
 sg13g2_decap_8 FILLER_106_684 ();
 sg13g2_decap_8 FILLER_106_691 ();
 sg13g2_decap_8 FILLER_106_698 ();
 sg13g2_decap_4 FILLER_106_705 ();
 sg13g2_fill_2 FILLER_106_724 ();
 sg13g2_decap_8 FILLER_106_735 ();
 sg13g2_decap_8 FILLER_106_742 ();
 sg13g2_decap_4 FILLER_106_749 ();
 sg13g2_decap_8 FILLER_106_769 ();
 sg13g2_decap_8 FILLER_106_776 ();
 sg13g2_decap_8 FILLER_106_783 ();
 sg13g2_decap_8 FILLER_106_790 ();
 sg13g2_fill_1 FILLER_106_797 ();
 sg13g2_decap_8 FILLER_106_806 ();
 sg13g2_decap_8 FILLER_106_813 ();
 sg13g2_decap_8 FILLER_106_820 ();
 sg13g2_decap_8 FILLER_106_837 ();
 sg13g2_decap_8 FILLER_106_866 ();
 sg13g2_decap_8 FILLER_106_873 ();
 sg13g2_decap_8 FILLER_106_880 ();
 sg13g2_decap_8 FILLER_106_887 ();
 sg13g2_decap_8 FILLER_106_894 ();
 sg13g2_decap_8 FILLER_106_901 ();
 sg13g2_decap_8 FILLER_106_908 ();
 sg13g2_decap_4 FILLER_106_915 ();
 sg13g2_decap_8 FILLER_106_923 ();
 sg13g2_fill_2 FILLER_106_930 ();
 sg13g2_fill_1 FILLER_106_963 ();
 sg13g2_decap_4 FILLER_106_973 ();
 sg13g2_fill_2 FILLER_106_977 ();
 sg13g2_decap_8 FILLER_106_1002 ();
 sg13g2_fill_2 FILLER_106_1009 ();
 sg13g2_fill_1 FILLER_106_1011 ();
 sg13g2_decap_8 FILLER_106_1021 ();
 sg13g2_decap_8 FILLER_106_1028 ();
 sg13g2_decap_8 FILLER_106_1035 ();
 sg13g2_decap_8 FILLER_106_1042 ();
 sg13g2_decap_8 FILLER_106_1049 ();
 sg13g2_decap_4 FILLER_106_1056 ();
 sg13g2_fill_1 FILLER_106_1060 ();
 sg13g2_decap_8 FILLER_106_1069 ();
 sg13g2_decap_4 FILLER_106_1076 ();
 sg13g2_fill_2 FILLER_106_1080 ();
 sg13g2_fill_2 FILLER_106_1095 ();
 sg13g2_decap_8 FILLER_106_1110 ();
 sg13g2_decap_8 FILLER_106_1117 ();
 sg13g2_decap_8 FILLER_106_1124 ();
 sg13g2_decap_8 FILLER_106_1131 ();
 sg13g2_decap_8 FILLER_106_1138 ();
 sg13g2_decap_8 FILLER_106_1145 ();
 sg13g2_decap_8 FILLER_106_1152 ();
 sg13g2_decap_8 FILLER_106_1159 ();
 sg13g2_decap_8 FILLER_106_1166 ();
 sg13g2_decap_8 FILLER_106_1173 ();
 sg13g2_fill_1 FILLER_106_1180 ();
 sg13g2_decap_4 FILLER_106_1185 ();
 sg13g2_fill_1 FILLER_106_1189 ();
 sg13g2_decap_8 FILLER_106_1219 ();
 sg13g2_decap_8 FILLER_106_1226 ();
 sg13g2_decap_8 FILLER_106_1233 ();
 sg13g2_decap_4 FILLER_106_1240 ();
 sg13g2_fill_2 FILLER_106_1244 ();
 sg13g2_decap_8 FILLER_106_1272 ();
 sg13g2_decap_8 FILLER_106_1279 ();
 sg13g2_fill_1 FILLER_106_1286 ();
 sg13g2_decap_8 FILLER_106_1300 ();
 sg13g2_decap_8 FILLER_106_1307 ();
 sg13g2_decap_8 FILLER_106_1314 ();
 sg13g2_fill_2 FILLER_106_1321 ();
 sg13g2_fill_1 FILLER_106_1323 ();
 sg13g2_decap_8 FILLER_106_1335 ();
 sg13g2_decap_8 FILLER_106_1342 ();
 sg13g2_decap_8 FILLER_106_1349 ();
 sg13g2_decap_4 FILLER_106_1356 ();
 sg13g2_fill_1 FILLER_106_1360 ();
 sg13g2_decap_8 FILLER_106_1366 ();
 sg13g2_decap_8 FILLER_106_1373 ();
 sg13g2_decap_8 FILLER_106_1380 ();
 sg13g2_decap_8 FILLER_106_1387 ();
 sg13g2_decap_8 FILLER_106_1394 ();
 sg13g2_decap_8 FILLER_106_1401 ();
 sg13g2_decap_8 FILLER_106_1408 ();
 sg13g2_decap_8 FILLER_106_1415 ();
 sg13g2_decap_8 FILLER_106_1422 ();
 sg13g2_decap_8 FILLER_106_1429 ();
 sg13g2_fill_1 FILLER_106_1436 ();
 sg13g2_decap_8 FILLER_106_1445 ();
 sg13g2_decap_8 FILLER_106_1452 ();
 sg13g2_fill_1 FILLER_106_1459 ();
 sg13g2_decap_4 FILLER_106_1464 ();
 sg13g2_decap_8 FILLER_106_1473 ();
 sg13g2_decap_8 FILLER_106_1480 ();
 sg13g2_decap_8 FILLER_106_1487 ();
 sg13g2_decap_8 FILLER_106_1494 ();
 sg13g2_decap_8 FILLER_106_1501 ();
 sg13g2_decap_8 FILLER_106_1508 ();
 sg13g2_decap_8 FILLER_106_1515 ();
 sg13g2_decap_8 FILLER_106_1522 ();
 sg13g2_decap_8 FILLER_106_1529 ();
 sg13g2_decap_8 FILLER_106_1536 ();
 sg13g2_decap_8 FILLER_106_1548 ();
 sg13g2_decap_8 FILLER_106_1555 ();
 sg13g2_decap_8 FILLER_106_1562 ();
 sg13g2_decap_8 FILLER_106_1569 ();
 sg13g2_decap_4 FILLER_106_1576 ();
 sg13g2_fill_2 FILLER_106_1580 ();
 sg13g2_decap_8 FILLER_106_1590 ();
 sg13g2_fill_1 FILLER_106_1597 ();
 sg13g2_decap_8 FILLER_106_1603 ();
 sg13g2_decap_8 FILLER_106_1610 ();
 sg13g2_decap_4 FILLER_106_1617 ();
 sg13g2_fill_1 FILLER_106_1621 ();
 sg13g2_decap_8 FILLER_106_1642 ();
 sg13g2_decap_8 FILLER_106_1649 ();
 sg13g2_decap_8 FILLER_106_1656 ();
 sg13g2_decap_4 FILLER_106_1663 ();
 sg13g2_fill_2 FILLER_106_1667 ();
 sg13g2_decap_8 FILLER_106_1673 ();
 sg13g2_decap_8 FILLER_106_1680 ();
 sg13g2_decap_8 FILLER_106_1687 ();
 sg13g2_decap_8 FILLER_106_1694 ();
 sg13g2_decap_8 FILLER_106_1701 ();
 sg13g2_decap_8 FILLER_106_1708 ();
 sg13g2_fill_1 FILLER_106_1715 ();
 sg13g2_decap_8 FILLER_106_1721 ();
 sg13g2_fill_2 FILLER_106_1728 ();
 sg13g2_fill_1 FILLER_106_1730 ();
 sg13g2_decap_8 FILLER_106_1735 ();
 sg13g2_decap_8 FILLER_106_1742 ();
 sg13g2_decap_8 FILLER_106_1749 ();
 sg13g2_decap_8 FILLER_106_1756 ();
 sg13g2_decap_4 FILLER_106_1763 ();
 sg13g2_fill_1 FILLER_106_1767 ();
 sg13g2_decap_8 FILLER_107_0 ();
 sg13g2_fill_2 FILLER_107_7 ();
 sg13g2_fill_1 FILLER_107_9 ();
 sg13g2_fill_2 FILLER_107_36 ();
 sg13g2_fill_1 FILLER_107_38 ();
 sg13g2_decap_8 FILLER_107_64 ();
 sg13g2_decap_4 FILLER_107_71 ();
 sg13g2_fill_1 FILLER_107_83 ();
 sg13g2_decap_8 FILLER_107_94 ();
 sg13g2_decap_4 FILLER_107_101 ();
 sg13g2_fill_2 FILLER_107_109 ();
 sg13g2_fill_2 FILLER_107_131 ();
 sg13g2_fill_1 FILLER_107_133 ();
 sg13g2_fill_2 FILLER_107_141 ();
 sg13g2_fill_1 FILLER_107_143 ();
 sg13g2_decap_8 FILLER_107_152 ();
 sg13g2_decap_8 FILLER_107_159 ();
 sg13g2_decap_8 FILLER_107_166 ();
 sg13g2_decap_8 FILLER_107_173 ();
 sg13g2_decap_8 FILLER_107_180 ();
 sg13g2_decap_8 FILLER_107_187 ();
 sg13g2_decap_8 FILLER_107_194 ();
 sg13g2_decap_8 FILLER_107_201 ();
 sg13g2_decap_8 FILLER_107_208 ();
 sg13g2_decap_4 FILLER_107_215 ();
 sg13g2_fill_1 FILLER_107_219 ();
 sg13g2_decap_8 FILLER_107_233 ();
 sg13g2_decap_8 FILLER_107_240 ();
 sg13g2_decap_8 FILLER_107_247 ();
 sg13g2_decap_8 FILLER_107_254 ();
 sg13g2_decap_8 FILLER_107_261 ();
 sg13g2_fill_2 FILLER_107_268 ();
 sg13g2_fill_1 FILLER_107_270 ();
 sg13g2_fill_2 FILLER_107_279 ();
 sg13g2_fill_1 FILLER_107_281 ();
 sg13g2_decap_8 FILLER_107_294 ();
 sg13g2_decap_8 FILLER_107_301 ();
 sg13g2_decap_8 FILLER_107_308 ();
 sg13g2_fill_2 FILLER_107_333 ();
 sg13g2_fill_1 FILLER_107_335 ();
 sg13g2_fill_2 FILLER_107_352 ();
 sg13g2_decap_8 FILLER_107_363 ();
 sg13g2_decap_8 FILLER_107_370 ();
 sg13g2_decap_8 FILLER_107_377 ();
 sg13g2_fill_2 FILLER_107_397 ();
 sg13g2_fill_1 FILLER_107_399 ();
 sg13g2_decap_8 FILLER_107_413 ();
 sg13g2_decap_8 FILLER_107_420 ();
 sg13g2_decap_8 FILLER_107_427 ();
 sg13g2_decap_8 FILLER_107_434 ();
 sg13g2_decap_8 FILLER_107_441 ();
 sg13g2_decap_8 FILLER_107_448 ();
 sg13g2_decap_8 FILLER_107_455 ();
 sg13g2_decap_4 FILLER_107_462 ();
 sg13g2_decap_8 FILLER_107_477 ();
 sg13g2_fill_2 FILLER_107_484 ();
 sg13g2_decap_8 FILLER_107_499 ();
 sg13g2_decap_8 FILLER_107_506 ();
 sg13g2_decap_8 FILLER_107_513 ();
 sg13g2_decap_8 FILLER_107_520 ();
 sg13g2_decap_8 FILLER_107_527 ();
 sg13g2_fill_2 FILLER_107_534 ();
 sg13g2_decap_8 FILLER_107_557 ();
 sg13g2_decap_8 FILLER_107_564 ();
 sg13g2_decap_8 FILLER_107_579 ();
 sg13g2_decap_8 FILLER_107_586 ();
 sg13g2_decap_8 FILLER_107_593 ();
 sg13g2_decap_8 FILLER_107_600 ();
 sg13g2_fill_2 FILLER_107_607 ();
 sg13g2_fill_2 FILLER_107_612 ();
 sg13g2_fill_1 FILLER_107_614 ();
 sg13g2_decap_8 FILLER_107_619 ();
 sg13g2_decap_8 FILLER_107_626 ();
 sg13g2_decap_8 FILLER_107_633 ();
 sg13g2_decap_4 FILLER_107_640 ();
 sg13g2_fill_2 FILLER_107_644 ();
 sg13g2_fill_2 FILLER_107_688 ();
 sg13g2_fill_2 FILLER_107_699 ();
 sg13g2_fill_1 FILLER_107_701 ();
 sg13g2_fill_2 FILLER_107_707 ();
 sg13g2_fill_1 FILLER_107_719 ();
 sg13g2_fill_1 FILLER_107_746 ();
 sg13g2_decap_8 FILLER_107_764 ();
 sg13g2_decap_8 FILLER_107_771 ();
 sg13g2_decap_8 FILLER_107_778 ();
 sg13g2_decap_8 FILLER_107_785 ();
 sg13g2_decap_8 FILLER_107_792 ();
 sg13g2_decap_4 FILLER_107_799 ();
 sg13g2_fill_1 FILLER_107_803 ();
 sg13g2_decap_8 FILLER_107_817 ();
 sg13g2_decap_8 FILLER_107_824 ();
 sg13g2_fill_1 FILLER_107_831 ();
 sg13g2_decap_8 FILLER_107_867 ();
 sg13g2_fill_2 FILLER_107_874 ();
 sg13g2_fill_1 FILLER_107_876 ();
 sg13g2_decap_8 FILLER_107_890 ();
 sg13g2_decap_8 FILLER_107_897 ();
 sg13g2_fill_2 FILLER_107_904 ();
 sg13g2_fill_1 FILLER_107_906 ();
 sg13g2_decap_8 FILLER_107_912 ();
 sg13g2_decap_8 FILLER_107_919 ();
 sg13g2_fill_2 FILLER_107_926 ();
 sg13g2_fill_1 FILLER_107_928 ();
 sg13g2_decap_4 FILLER_107_935 ();
 sg13g2_decap_4 FILLER_107_943 ();
 sg13g2_fill_1 FILLER_107_947 ();
 sg13g2_decap_8 FILLER_107_952 ();
 sg13g2_decap_4 FILLER_107_959 ();
 sg13g2_fill_1 FILLER_107_963 ();
 sg13g2_decap_8 FILLER_107_977 ();
 sg13g2_decap_8 FILLER_107_984 ();
 sg13g2_decap_8 FILLER_107_991 ();
 sg13g2_decap_4 FILLER_107_998 ();
 sg13g2_decap_8 FILLER_107_1007 ();
 sg13g2_decap_8 FILLER_107_1045 ();
 sg13g2_fill_2 FILLER_107_1052 ();
 sg13g2_fill_1 FILLER_107_1054 ();
 sg13g2_decap_8 FILLER_107_1059 ();
 sg13g2_decap_8 FILLER_107_1066 ();
 sg13g2_decap_8 FILLER_107_1073 ();
 sg13g2_decap_8 FILLER_107_1080 ();
 sg13g2_decap_4 FILLER_107_1087 ();
 sg13g2_fill_2 FILLER_107_1091 ();
 sg13g2_decap_8 FILLER_107_1097 ();
 sg13g2_decap_8 FILLER_107_1104 ();
 sg13g2_decap_8 FILLER_107_1111 ();
 sg13g2_decap_8 FILLER_107_1118 ();
 sg13g2_decap_8 FILLER_107_1125 ();
 sg13g2_decap_8 FILLER_107_1132 ();
 sg13g2_decap_8 FILLER_107_1139 ();
 sg13g2_decap_8 FILLER_107_1146 ();
 sg13g2_decap_8 FILLER_107_1153 ();
 sg13g2_decap_8 FILLER_107_1160 ();
 sg13g2_decap_8 FILLER_107_1167 ();
 sg13g2_decap_8 FILLER_107_1174 ();
 sg13g2_decap_8 FILLER_107_1181 ();
 sg13g2_decap_8 FILLER_107_1188 ();
 sg13g2_decap_8 FILLER_107_1195 ();
 sg13g2_decap_8 FILLER_107_1202 ();
 sg13g2_fill_2 FILLER_107_1209 ();
 sg13g2_fill_1 FILLER_107_1211 ();
 sg13g2_decap_8 FILLER_107_1233 ();
 sg13g2_decap_8 FILLER_107_1240 ();
 sg13g2_decap_8 FILLER_107_1247 ();
 sg13g2_decap_4 FILLER_107_1254 ();
 sg13g2_fill_2 FILLER_107_1258 ();
 sg13g2_decap_8 FILLER_107_1273 ();
 sg13g2_decap_4 FILLER_107_1280 ();
 sg13g2_decap_8 FILLER_107_1297 ();
 sg13g2_decap_8 FILLER_107_1304 ();
 sg13g2_decap_4 FILLER_107_1311 ();
 sg13g2_fill_1 FILLER_107_1315 ();
 sg13g2_decap_8 FILLER_107_1381 ();
 sg13g2_decap_8 FILLER_107_1388 ();
 sg13g2_decap_8 FILLER_107_1395 ();
 sg13g2_decap_8 FILLER_107_1402 ();
 sg13g2_fill_2 FILLER_107_1409 ();
 sg13g2_fill_1 FILLER_107_1411 ();
 sg13g2_decap_8 FILLER_107_1420 ();
 sg13g2_decap_8 FILLER_107_1427 ();
 sg13g2_decap_8 FILLER_107_1434 ();
 sg13g2_decap_8 FILLER_107_1441 ();
 sg13g2_decap_8 FILLER_107_1448 ();
 sg13g2_decap_8 FILLER_107_1455 ();
 sg13g2_decap_8 FILLER_107_1462 ();
 sg13g2_decap_8 FILLER_107_1469 ();
 sg13g2_decap_4 FILLER_107_1476 ();
 sg13g2_fill_2 FILLER_107_1480 ();
 sg13g2_decap_8 FILLER_107_1490 ();
 sg13g2_decap_8 FILLER_107_1497 ();
 sg13g2_decap_8 FILLER_107_1504 ();
 sg13g2_decap_8 FILLER_107_1511 ();
 sg13g2_decap_4 FILLER_107_1518 ();
 sg13g2_decap_8 FILLER_107_1530 ();
 sg13g2_decap_8 FILLER_107_1537 ();
 sg13g2_decap_8 FILLER_107_1544 ();
 sg13g2_decap_8 FILLER_107_1551 ();
 sg13g2_fill_1 FILLER_107_1558 ();
 sg13g2_decap_8 FILLER_107_1562 ();
 sg13g2_decap_8 FILLER_107_1569 ();
 sg13g2_decap_8 FILLER_107_1576 ();
 sg13g2_decap_8 FILLER_107_1583 ();
 sg13g2_fill_1 FILLER_107_1590 ();
 sg13g2_decap_8 FILLER_107_1612 ();
 sg13g2_decap_8 FILLER_107_1619 ();
 sg13g2_decap_8 FILLER_107_1626 ();
 sg13g2_decap_8 FILLER_107_1633 ();
 sg13g2_decap_4 FILLER_107_1640 ();
 sg13g2_fill_2 FILLER_107_1644 ();
 sg13g2_decap_8 FILLER_107_1658 ();
 sg13g2_decap_8 FILLER_107_1665 ();
 sg13g2_decap_8 FILLER_107_1672 ();
 sg13g2_decap_8 FILLER_107_1679 ();
 sg13g2_decap_8 FILLER_107_1686 ();
 sg13g2_decap_8 FILLER_107_1693 ();
 sg13g2_decap_8 FILLER_107_1700 ();
 sg13g2_decap_8 FILLER_107_1707 ();
 sg13g2_fill_2 FILLER_107_1739 ();
 sg13g2_fill_1 FILLER_107_1741 ();
 sg13g2_decap_8 FILLER_107_1752 ();
 sg13g2_decap_8 FILLER_107_1759 ();
 sg13g2_fill_2 FILLER_107_1766 ();
 sg13g2_decap_8 FILLER_108_0 ();
 sg13g2_decap_8 FILLER_108_7 ();
 sg13g2_decap_4 FILLER_108_14 ();
 sg13g2_fill_1 FILLER_108_18 ();
 sg13g2_decap_8 FILLER_108_47 ();
 sg13g2_decap_8 FILLER_108_54 ();
 sg13g2_decap_8 FILLER_108_61 ();
 sg13g2_fill_1 FILLER_108_68 ();
 sg13g2_decap_8 FILLER_108_77 ();
 sg13g2_decap_8 FILLER_108_89 ();
 sg13g2_fill_1 FILLER_108_96 ();
 sg13g2_fill_1 FILLER_108_110 ();
 sg13g2_decap_4 FILLER_108_121 ();
 sg13g2_decap_4 FILLER_108_133 ();
 sg13g2_fill_2 FILLER_108_137 ();
 sg13g2_decap_8 FILLER_108_147 ();
 sg13g2_decap_8 FILLER_108_154 ();
 sg13g2_decap_8 FILLER_108_161 ();
 sg13g2_decap_8 FILLER_108_168 ();
 sg13g2_decap_8 FILLER_108_175 ();
 sg13g2_decap_8 FILLER_108_182 ();
 sg13g2_fill_1 FILLER_108_189 ();
 sg13g2_decap_8 FILLER_108_198 ();
 sg13g2_decap_8 FILLER_108_205 ();
 sg13g2_decap_8 FILLER_108_212 ();
 sg13g2_decap_4 FILLER_108_219 ();
 sg13g2_fill_1 FILLER_108_223 ();
 sg13g2_fill_1 FILLER_108_236 ();
 sg13g2_decap_8 FILLER_108_245 ();
 sg13g2_decap_8 FILLER_108_252 ();
 sg13g2_decap_8 FILLER_108_259 ();
 sg13g2_decap_8 FILLER_108_266 ();
 sg13g2_decap_8 FILLER_108_273 ();
 sg13g2_fill_2 FILLER_108_280 ();
 sg13g2_decap_4 FILLER_108_286 ();
 sg13g2_fill_1 FILLER_108_290 ();
 sg13g2_decap_8 FILLER_108_303 ();
 sg13g2_decap_8 FILLER_108_310 ();
 sg13g2_decap_8 FILLER_108_317 ();
 sg13g2_decap_8 FILLER_108_324 ();
 sg13g2_decap_4 FILLER_108_331 ();
 sg13g2_fill_2 FILLER_108_335 ();
 sg13g2_decap_4 FILLER_108_340 ();
 sg13g2_decap_8 FILLER_108_364 ();
 sg13g2_decap_8 FILLER_108_371 ();
 sg13g2_decap_8 FILLER_108_378 ();
 sg13g2_fill_2 FILLER_108_385 ();
 sg13g2_decap_8 FILLER_108_418 ();
 sg13g2_decap_8 FILLER_108_425 ();
 sg13g2_fill_2 FILLER_108_432 ();
 sg13g2_fill_1 FILLER_108_434 ();
 sg13g2_decap_8 FILLER_108_443 ();
 sg13g2_fill_1 FILLER_108_450 ();
 sg13g2_decap_8 FILLER_108_460 ();
 sg13g2_decap_8 FILLER_108_467 ();
 sg13g2_decap_8 FILLER_108_474 ();
 sg13g2_decap_8 FILLER_108_481 ();
 sg13g2_decap_8 FILLER_108_488 ();
 sg13g2_decap_8 FILLER_108_495 ();
 sg13g2_decap_8 FILLER_108_502 ();
 sg13g2_decap_8 FILLER_108_509 ();
 sg13g2_decap_8 FILLER_108_516 ();
 sg13g2_decap_4 FILLER_108_523 ();
 sg13g2_fill_1 FILLER_108_527 ();
 sg13g2_decap_8 FILLER_108_540 ();
 sg13g2_fill_2 FILLER_108_547 ();
 sg13g2_fill_1 FILLER_108_549 ();
 sg13g2_decap_8 FILLER_108_558 ();
 sg13g2_decap_4 FILLER_108_565 ();
 sg13g2_fill_1 FILLER_108_569 ();
 sg13g2_decap_8 FILLER_108_580 ();
 sg13g2_decap_8 FILLER_108_587 ();
 sg13g2_decap_8 FILLER_108_594 ();
 sg13g2_fill_2 FILLER_108_601 ();
 sg13g2_decap_8 FILLER_108_626 ();
 sg13g2_decap_8 FILLER_108_633 ();
 sg13g2_decap_8 FILLER_108_640 ();
 sg13g2_fill_1 FILLER_108_647 ();
 sg13g2_decap_8 FILLER_108_665 ();
 sg13g2_decap_8 FILLER_108_672 ();
 sg13g2_decap_8 FILLER_108_679 ();
 sg13g2_decap_8 FILLER_108_686 ();
 sg13g2_decap_8 FILLER_108_693 ();
 sg13g2_decap_8 FILLER_108_700 ();
 sg13g2_fill_1 FILLER_108_723 ();
 sg13g2_decap_8 FILLER_108_728 ();
 sg13g2_decap_4 FILLER_108_735 ();
 sg13g2_fill_2 FILLER_108_739 ();
 sg13g2_decap_4 FILLER_108_745 ();
 sg13g2_fill_2 FILLER_108_749 ();
 sg13g2_decap_8 FILLER_108_770 ();
 sg13g2_decap_8 FILLER_108_777 ();
 sg13g2_decap_8 FILLER_108_784 ();
 sg13g2_decap_8 FILLER_108_791 ();
 sg13g2_fill_2 FILLER_108_798 ();
 sg13g2_decap_8 FILLER_108_826 ();
 sg13g2_decap_4 FILLER_108_833 ();
 sg13g2_fill_2 FILLER_108_837 ();
 sg13g2_decap_8 FILLER_108_845 ();
 sg13g2_decap_8 FILLER_108_856 ();
 sg13g2_decap_8 FILLER_108_863 ();
 sg13g2_decap_8 FILLER_108_870 ();
 sg13g2_fill_1 FILLER_108_877 ();
 sg13g2_decap_8 FILLER_108_904 ();
 sg13g2_decap_8 FILLER_108_911 ();
 sg13g2_decap_8 FILLER_108_918 ();
 sg13g2_decap_8 FILLER_108_925 ();
 sg13g2_decap_8 FILLER_108_932 ();
 sg13g2_decap_8 FILLER_108_947 ();
 sg13g2_decap_8 FILLER_108_954 ();
 sg13g2_decap_8 FILLER_108_961 ();
 sg13g2_decap_8 FILLER_108_968 ();
 sg13g2_fill_2 FILLER_108_975 ();
 sg13g2_fill_1 FILLER_108_977 ();
 sg13g2_decap_8 FILLER_108_991 ();
 sg13g2_decap_8 FILLER_108_998 ();
 sg13g2_decap_8 FILLER_108_1005 ();
 sg13g2_decap_8 FILLER_108_1012 ();
 sg13g2_decap_8 FILLER_108_1019 ();
 sg13g2_decap_4 FILLER_108_1026 ();
 sg13g2_decap_8 FILLER_108_1034 ();
 sg13g2_decap_8 FILLER_108_1041 ();
 sg13g2_fill_2 FILLER_108_1061 ();
 sg13g2_fill_1 FILLER_108_1063 ();
 sg13g2_decap_8 FILLER_108_1072 ();
 sg13g2_decap_8 FILLER_108_1079 ();
 sg13g2_decap_8 FILLER_108_1086 ();
 sg13g2_decap_8 FILLER_108_1093 ();
 sg13g2_decap_8 FILLER_108_1100 ();
 sg13g2_decap_8 FILLER_108_1107 ();
 sg13g2_decap_8 FILLER_108_1114 ();
 sg13g2_decap_8 FILLER_108_1121 ();
 sg13g2_fill_2 FILLER_108_1128 ();
 sg13g2_fill_1 FILLER_108_1134 ();
 sg13g2_decap_8 FILLER_108_1140 ();
 sg13g2_decap_8 FILLER_108_1147 ();
 sg13g2_fill_2 FILLER_108_1154 ();
 sg13g2_decap_8 FILLER_108_1169 ();
 sg13g2_decap_8 FILLER_108_1176 ();
 sg13g2_decap_8 FILLER_108_1183 ();
 sg13g2_fill_2 FILLER_108_1190 ();
 sg13g2_fill_1 FILLER_108_1192 ();
 sg13g2_decap_4 FILLER_108_1201 ();
 sg13g2_fill_2 FILLER_108_1205 ();
 sg13g2_decap_8 FILLER_108_1213 ();
 sg13g2_decap_4 FILLER_108_1220 ();
 sg13g2_fill_2 FILLER_108_1224 ();
 sg13g2_decap_8 FILLER_108_1239 ();
 sg13g2_decap_8 FILLER_108_1246 ();
 sg13g2_decap_4 FILLER_108_1264 ();
 sg13g2_fill_2 FILLER_108_1268 ();
 sg13g2_decap_8 FILLER_108_1299 ();
 sg13g2_fill_1 FILLER_108_1306 ();
 sg13g2_decap_4 FILLER_108_1315 ();
 sg13g2_decap_8 FILLER_108_1335 ();
 sg13g2_decap_8 FILLER_108_1342 ();
 sg13g2_decap_4 FILLER_108_1349 ();
 sg13g2_decap_8 FILLER_108_1357 ();
 sg13g2_decap_4 FILLER_108_1364 ();
 sg13g2_decap_8 FILLER_108_1377 ();
 sg13g2_decap_4 FILLER_108_1384 ();
 sg13g2_fill_1 FILLER_108_1388 ();
 sg13g2_decap_8 FILLER_108_1405 ();
 sg13g2_fill_2 FILLER_108_1412 ();
 sg13g2_decap_8 FILLER_108_1422 ();
 sg13g2_decap_8 FILLER_108_1429 ();
 sg13g2_decap_8 FILLER_108_1436 ();
 sg13g2_decap_8 FILLER_108_1443 ();
 sg13g2_decap_8 FILLER_108_1450 ();
 sg13g2_decap_8 FILLER_108_1457 ();
 sg13g2_decap_8 FILLER_108_1464 ();
 sg13g2_decap_4 FILLER_108_1471 ();
 sg13g2_decap_8 FILLER_108_1488 ();
 sg13g2_decap_4 FILLER_108_1495 ();
 sg13g2_fill_1 FILLER_108_1499 ();
 sg13g2_decap_8 FILLER_108_1508 ();
 sg13g2_decap_8 FILLER_108_1515 ();
 sg13g2_decap_8 FILLER_108_1522 ();
 sg13g2_decap_8 FILLER_108_1529 ();
 sg13g2_decap_8 FILLER_108_1536 ();
 sg13g2_decap_4 FILLER_108_1543 ();
 sg13g2_fill_1 FILLER_108_1547 ();
 sg13g2_fill_1 FILLER_108_1568 ();
 sg13g2_decap_8 FILLER_108_1578 ();
 sg13g2_decap_4 FILLER_108_1585 ();
 sg13g2_fill_1 FILLER_108_1589 ();
 sg13g2_decap_4 FILLER_108_1598 ();
 sg13g2_fill_1 FILLER_108_1602 ();
 sg13g2_decap_8 FILLER_108_1611 ();
 sg13g2_decap_8 FILLER_108_1618 ();
 sg13g2_decap_8 FILLER_108_1625 ();
 sg13g2_fill_2 FILLER_108_1642 ();
 sg13g2_decap_8 FILLER_108_1652 ();
 sg13g2_decap_8 FILLER_108_1659 ();
 sg13g2_decap_8 FILLER_108_1666 ();
 sg13g2_decap_8 FILLER_108_1673 ();
 sg13g2_decap_8 FILLER_108_1680 ();
 sg13g2_decap_8 FILLER_108_1687 ();
 sg13g2_decap_8 FILLER_108_1694 ();
 sg13g2_decap_8 FILLER_108_1701 ();
 sg13g2_decap_4 FILLER_108_1708 ();
 sg13g2_fill_1 FILLER_108_1712 ();
 sg13g2_fill_1 FILLER_108_1717 ();
 sg13g2_fill_2 FILLER_108_1739 ();
 sg13g2_decap_8 FILLER_108_1759 ();
 sg13g2_fill_2 FILLER_108_1766 ();
 sg13g2_decap_8 FILLER_109_0 ();
 sg13g2_decap_8 FILLER_109_7 ();
 sg13g2_decap_8 FILLER_109_14 ();
 sg13g2_decap_8 FILLER_109_21 ();
 sg13g2_decap_8 FILLER_109_28 ();
 sg13g2_decap_8 FILLER_109_35 ();
 sg13g2_decap_8 FILLER_109_42 ();
 sg13g2_fill_1 FILLER_109_49 ();
 sg13g2_fill_2 FILLER_109_58 ();
 sg13g2_decap_8 FILLER_109_64 ();
 sg13g2_decap_8 FILLER_109_71 ();
 sg13g2_decap_8 FILLER_109_78 ();
 sg13g2_decap_8 FILLER_109_85 ();
 sg13g2_decap_8 FILLER_109_92 ();
 sg13g2_decap_4 FILLER_109_99 ();
 sg13g2_fill_2 FILLER_109_103 ();
 sg13g2_decap_8 FILLER_109_109 ();
 sg13g2_decap_8 FILLER_109_116 ();
 sg13g2_decap_8 FILLER_109_123 ();
 sg13g2_decap_8 FILLER_109_130 ();
 sg13g2_fill_1 FILLER_109_137 ();
 sg13g2_decap_4 FILLER_109_141 ();
 sg13g2_fill_2 FILLER_109_145 ();
 sg13g2_decap_8 FILLER_109_156 ();
 sg13g2_decap_8 FILLER_109_163 ();
 sg13g2_decap_8 FILLER_109_170 ();
 sg13g2_decap_8 FILLER_109_177 ();
 sg13g2_decap_4 FILLER_109_184 ();
 sg13g2_fill_1 FILLER_109_188 ();
 sg13g2_fill_1 FILLER_109_205 ();
 sg13g2_decap_4 FILLER_109_214 ();
 sg13g2_fill_2 FILLER_109_218 ();
 sg13g2_decap_8 FILLER_109_228 ();
 sg13g2_decap_8 FILLER_109_240 ();
 sg13g2_decap_8 FILLER_109_247 ();
 sg13g2_decap_8 FILLER_109_262 ();
 sg13g2_decap_4 FILLER_109_269 ();
 sg13g2_fill_2 FILLER_109_277 ();
 sg13g2_decap_8 FILLER_109_287 ();
 sg13g2_decap_8 FILLER_109_294 ();
 sg13g2_decap_8 FILLER_109_301 ();
 sg13g2_decap_8 FILLER_109_308 ();
 sg13g2_decap_8 FILLER_109_315 ();
 sg13g2_decap_8 FILLER_109_322 ();
 sg13g2_decap_8 FILLER_109_329 ();
 sg13g2_fill_1 FILLER_109_336 ();
 sg13g2_decap_8 FILLER_109_342 ();
 sg13g2_decap_8 FILLER_109_349 ();
 sg13g2_decap_8 FILLER_109_356 ();
 sg13g2_decap_8 FILLER_109_363 ();
 sg13g2_decap_8 FILLER_109_370 ();
 sg13g2_fill_2 FILLER_109_377 ();
 sg13g2_fill_1 FILLER_109_379 ();
 sg13g2_decap_8 FILLER_109_397 ();
 sg13g2_decap_8 FILLER_109_404 ();
 sg13g2_decap_8 FILLER_109_411 ();
 sg13g2_decap_8 FILLER_109_418 ();
 sg13g2_decap_8 FILLER_109_425 ();
 sg13g2_decap_8 FILLER_109_432 ();
 sg13g2_decap_8 FILLER_109_447 ();
 sg13g2_decap_8 FILLER_109_454 ();
 sg13g2_decap_8 FILLER_109_461 ();
 sg13g2_decap_8 FILLER_109_468 ();
 sg13g2_decap_8 FILLER_109_475 ();
 sg13g2_fill_1 FILLER_109_482 ();
 sg13g2_decap_8 FILLER_109_508 ();
 sg13g2_decap_8 FILLER_109_515 ();
 sg13g2_decap_4 FILLER_109_522 ();
 sg13g2_fill_2 FILLER_109_526 ();
 sg13g2_decap_8 FILLER_109_541 ();
 sg13g2_decap_4 FILLER_109_548 ();
 sg13g2_fill_2 FILLER_109_552 ();
 sg13g2_decap_8 FILLER_109_583 ();
 sg13g2_decap_8 FILLER_109_590 ();
 sg13g2_fill_2 FILLER_109_597 ();
 sg13g2_fill_1 FILLER_109_599 ();
 sg13g2_decap_8 FILLER_109_647 ();
 sg13g2_decap_4 FILLER_109_654 ();
 sg13g2_decap_8 FILLER_109_676 ();
 sg13g2_decap_8 FILLER_109_683 ();
 sg13g2_fill_1 FILLER_109_690 ();
 sg13g2_decap_8 FILLER_109_696 ();
 sg13g2_decap_8 FILLER_109_703 ();
 sg13g2_decap_8 FILLER_109_710 ();
 sg13g2_decap_8 FILLER_109_717 ();
 sg13g2_decap_8 FILLER_109_724 ();
 sg13g2_decap_8 FILLER_109_731 ();
 sg13g2_decap_8 FILLER_109_738 ();
 sg13g2_decap_8 FILLER_109_745 ();
 sg13g2_decap_8 FILLER_109_752 ();
 sg13g2_decap_8 FILLER_109_759 ();
 sg13g2_decap_8 FILLER_109_766 ();
 sg13g2_decap_8 FILLER_109_773 ();
 sg13g2_decap_8 FILLER_109_780 ();
 sg13g2_decap_8 FILLER_109_787 ();
 sg13g2_decap_8 FILLER_109_794 ();
 sg13g2_decap_8 FILLER_109_801 ();
 sg13g2_fill_2 FILLER_109_808 ();
 sg13g2_fill_1 FILLER_109_810 ();
 sg13g2_decap_8 FILLER_109_815 ();
 sg13g2_decap_8 FILLER_109_822 ();
 sg13g2_decap_8 FILLER_109_829 ();
 sg13g2_decap_4 FILLER_109_836 ();
 sg13g2_fill_1 FILLER_109_840 ();
 sg13g2_decap_8 FILLER_109_850 ();
 sg13g2_decap_8 FILLER_109_857 ();
 sg13g2_decap_8 FILLER_109_864 ();
 sg13g2_decap_8 FILLER_109_871 ();
 sg13g2_decap_8 FILLER_109_878 ();
 sg13g2_decap_4 FILLER_109_885 ();
 sg13g2_fill_1 FILLER_109_893 ();
 sg13g2_decap_8 FILLER_109_898 ();
 sg13g2_decap_8 FILLER_109_905 ();
 sg13g2_decap_8 FILLER_109_912 ();
 sg13g2_decap_8 FILLER_109_919 ();
 sg13g2_decap_8 FILLER_109_926 ();
 sg13g2_decap_4 FILLER_109_933 ();
 sg13g2_fill_1 FILLER_109_937 ();
 sg13g2_decap_8 FILLER_109_951 ();
 sg13g2_decap_8 FILLER_109_958 ();
 sg13g2_decap_8 FILLER_109_965 ();
 sg13g2_decap_8 FILLER_109_972 ();
 sg13g2_decap_8 FILLER_109_979 ();
 sg13g2_decap_8 FILLER_109_986 ();
 sg13g2_decap_8 FILLER_109_993 ();
 sg13g2_decap_8 FILLER_109_1000 ();
 sg13g2_decap_8 FILLER_109_1007 ();
 sg13g2_decap_8 FILLER_109_1014 ();
 sg13g2_decap_8 FILLER_109_1021 ();
 sg13g2_decap_8 FILLER_109_1028 ();
 sg13g2_decap_8 FILLER_109_1035 ();
 sg13g2_decap_8 FILLER_109_1042 ();
 sg13g2_decap_8 FILLER_109_1049 ();
 sg13g2_decap_8 FILLER_109_1056 ();
 sg13g2_decap_8 FILLER_109_1063 ();
 sg13g2_decap_8 FILLER_109_1070 ();
 sg13g2_decap_8 FILLER_109_1077 ();
 sg13g2_decap_4 FILLER_109_1084 ();
 sg13g2_fill_2 FILLER_109_1088 ();
 sg13g2_decap_8 FILLER_109_1094 ();
 sg13g2_decap_4 FILLER_109_1101 ();
 sg13g2_fill_1 FILLER_109_1105 ();
 sg13g2_decap_8 FILLER_109_1145 ();
 sg13g2_decap_8 FILLER_109_1177 ();
 sg13g2_decap_8 FILLER_109_1184 ();
 sg13g2_decap_8 FILLER_109_1191 ();
 sg13g2_fill_2 FILLER_109_1198 ();
 sg13g2_fill_1 FILLER_109_1200 ();
 sg13g2_decap_8 FILLER_109_1215 ();
 sg13g2_decap_4 FILLER_109_1222 ();
 sg13g2_fill_1 FILLER_109_1252 ();
 sg13g2_decap_8 FILLER_109_1258 ();
 sg13g2_decap_8 FILLER_109_1265 ();
 sg13g2_fill_2 FILLER_109_1272 ();
 sg13g2_decap_8 FILLER_109_1287 ();
 sg13g2_decap_8 FILLER_109_1294 ();
 sg13g2_decap_8 FILLER_109_1301 ();
 sg13g2_decap_8 FILLER_109_1308 ();
 sg13g2_decap_8 FILLER_109_1315 ();
 sg13g2_decap_8 FILLER_109_1322 ();
 sg13g2_decap_8 FILLER_109_1329 ();
 sg13g2_decap_8 FILLER_109_1336 ();
 sg13g2_decap_8 FILLER_109_1343 ();
 sg13g2_decap_8 FILLER_109_1350 ();
 sg13g2_decap_8 FILLER_109_1357 ();
 sg13g2_decap_4 FILLER_109_1364 ();
 sg13g2_fill_2 FILLER_109_1368 ();
 sg13g2_decap_8 FILLER_109_1380 ();
 sg13g2_fill_2 FILLER_109_1387 ();
 sg13g2_decap_8 FILLER_109_1394 ();
 sg13g2_decap_8 FILLER_109_1401 ();
 sg13g2_decap_8 FILLER_109_1408 ();
 sg13g2_decap_4 FILLER_109_1415 ();
 sg13g2_fill_1 FILLER_109_1419 ();
 sg13g2_fill_2 FILLER_109_1425 ();
 sg13g2_fill_1 FILLER_109_1427 ();
 sg13g2_decap_8 FILLER_109_1433 ();
 sg13g2_fill_2 FILLER_109_1440 ();
 sg13g2_decap_8 FILLER_109_1450 ();
 sg13g2_decap_8 FILLER_109_1457 ();
 sg13g2_fill_2 FILLER_109_1464 ();
 sg13g2_fill_1 FILLER_109_1466 ();
 sg13g2_fill_1 FILLER_109_1472 ();
 sg13g2_fill_1 FILLER_109_1483 ();
 sg13g2_decap_8 FILLER_109_1490 ();
 sg13g2_decap_8 FILLER_109_1497 ();
 sg13g2_decap_8 FILLER_109_1504 ();
 sg13g2_fill_2 FILLER_109_1511 ();
 sg13g2_decap_4 FILLER_109_1529 ();
 sg13g2_decap_4 FILLER_109_1541 ();
 sg13g2_fill_2 FILLER_109_1545 ();
 sg13g2_decap_4 FILLER_109_1555 ();
 sg13g2_decap_8 FILLER_109_1590 ();
 sg13g2_decap_8 FILLER_109_1597 ();
 sg13g2_decap_8 FILLER_109_1604 ();
 sg13g2_decap_8 FILLER_109_1611 ();
 sg13g2_decap_8 FILLER_109_1618 ();
 sg13g2_decap_8 FILLER_109_1645 ();
 sg13g2_decap_8 FILLER_109_1652 ();
 sg13g2_decap_8 FILLER_109_1659 ();
 sg13g2_fill_2 FILLER_109_1666 ();
 sg13g2_fill_1 FILLER_109_1668 ();
 sg13g2_decap_4 FILLER_109_1677 ();
 sg13g2_decap_8 FILLER_109_1694 ();
 sg13g2_decap_8 FILLER_109_1701 ();
 sg13g2_decap_8 FILLER_109_1708 ();
 sg13g2_decap_8 FILLER_109_1715 ();
 sg13g2_decap_4 FILLER_109_1722 ();
 sg13g2_fill_2 FILLER_109_1726 ();
 sg13g2_decap_8 FILLER_109_1740 ();
 sg13g2_decap_8 FILLER_109_1747 ();
 sg13g2_decap_8 FILLER_109_1754 ();
 sg13g2_decap_8 FILLER_109_1761 ();
 sg13g2_decap_8 FILLER_110_0 ();
 sg13g2_decap_8 FILLER_110_7 ();
 sg13g2_decap_8 FILLER_110_14 ();
 sg13g2_decap_8 FILLER_110_21 ();
 sg13g2_decap_8 FILLER_110_28 ();
 sg13g2_decap_8 FILLER_110_35 ();
 sg13g2_decap_8 FILLER_110_42 ();
 sg13g2_decap_8 FILLER_110_49 ();
 sg13g2_fill_2 FILLER_110_56 ();
 sg13g2_fill_1 FILLER_110_58 ();
 sg13g2_decap_8 FILLER_110_68 ();
 sg13g2_decap_8 FILLER_110_75 ();
 sg13g2_decap_4 FILLER_110_82 ();
 sg13g2_decap_8 FILLER_110_93 ();
 sg13g2_decap_8 FILLER_110_100 ();
 sg13g2_decap_8 FILLER_110_107 ();
 sg13g2_decap_8 FILLER_110_114 ();
 sg13g2_decap_8 FILLER_110_121 ();
 sg13g2_decap_8 FILLER_110_128 ();
 sg13g2_decap_8 FILLER_110_155 ();
 sg13g2_decap_8 FILLER_110_162 ();
 sg13g2_decap_8 FILLER_110_169 ();
 sg13g2_decap_4 FILLER_110_176 ();
 sg13g2_fill_1 FILLER_110_180 ();
 sg13g2_fill_1 FILLER_110_202 ();
 sg13g2_decap_8 FILLER_110_208 ();
 sg13g2_decap_8 FILLER_110_215 ();
 sg13g2_decap_8 FILLER_110_222 ();
 sg13g2_decap_8 FILLER_110_229 ();
 sg13g2_decap_8 FILLER_110_236 ();
 sg13g2_decap_8 FILLER_110_243 ();
 sg13g2_decap_8 FILLER_110_250 ();
 sg13g2_decap_8 FILLER_110_257 ();
 sg13g2_decap_8 FILLER_110_264 ();
 sg13g2_fill_2 FILLER_110_271 ();
 sg13g2_decap_4 FILLER_110_284 ();
 sg13g2_fill_1 FILLER_110_288 ();
 sg13g2_decap_8 FILLER_110_293 ();
 sg13g2_decap_8 FILLER_110_300 ();
 sg13g2_decap_8 FILLER_110_307 ();
 sg13g2_decap_8 FILLER_110_314 ();
 sg13g2_decap_8 FILLER_110_321 ();
 sg13g2_decap_8 FILLER_110_328 ();
 sg13g2_decap_8 FILLER_110_335 ();
 sg13g2_decap_8 FILLER_110_342 ();
 sg13g2_decap_8 FILLER_110_349 ();
 sg13g2_decap_8 FILLER_110_356 ();
 sg13g2_fill_2 FILLER_110_363 ();
 sg13g2_fill_1 FILLER_110_365 ();
 sg13g2_decap_4 FILLER_110_379 ();
 sg13g2_decap_8 FILLER_110_394 ();
 sg13g2_decap_8 FILLER_110_401 ();
 sg13g2_decap_8 FILLER_110_408 ();
 sg13g2_decap_8 FILLER_110_415 ();
 sg13g2_decap_8 FILLER_110_422 ();
 sg13g2_decap_8 FILLER_110_429 ();
 sg13g2_decap_8 FILLER_110_436 ();
 sg13g2_fill_2 FILLER_110_443 ();
 sg13g2_fill_1 FILLER_110_445 ();
 sg13g2_decap_8 FILLER_110_451 ();
 sg13g2_decap_8 FILLER_110_458 ();
 sg13g2_decap_8 FILLER_110_465 ();
 sg13g2_decap_8 FILLER_110_472 ();
 sg13g2_decap_8 FILLER_110_479 ();
 sg13g2_fill_2 FILLER_110_486 ();
 sg13g2_decap_8 FILLER_110_513 ();
 sg13g2_decap_8 FILLER_110_520 ();
 sg13g2_decap_8 FILLER_110_527 ();
 sg13g2_decap_8 FILLER_110_534 ();
 sg13g2_decap_8 FILLER_110_541 ();
 sg13g2_decap_8 FILLER_110_548 ();
 sg13g2_decap_8 FILLER_110_555 ();
 sg13g2_decap_8 FILLER_110_562 ();
 sg13g2_decap_8 FILLER_110_569 ();
 sg13g2_decap_8 FILLER_110_576 ();
 sg13g2_decap_8 FILLER_110_583 ();
 sg13g2_decap_8 FILLER_110_590 ();
 sg13g2_decap_4 FILLER_110_597 ();
 sg13g2_fill_1 FILLER_110_601 ();
 sg13g2_decap_8 FILLER_110_635 ();
 sg13g2_decap_8 FILLER_110_642 ();
 sg13g2_decap_4 FILLER_110_649 ();
 sg13g2_fill_2 FILLER_110_653 ();
 sg13g2_decap_8 FILLER_110_660 ();
 sg13g2_decap_8 FILLER_110_667 ();
 sg13g2_decap_8 FILLER_110_674 ();
 sg13g2_decap_8 FILLER_110_681 ();
 sg13g2_decap_8 FILLER_110_688 ();
 sg13g2_decap_8 FILLER_110_695 ();
 sg13g2_fill_1 FILLER_110_702 ();
 sg13g2_decap_8 FILLER_110_707 ();
 sg13g2_decap_8 FILLER_110_714 ();
 sg13g2_decap_8 FILLER_110_721 ();
 sg13g2_decap_8 FILLER_110_728 ();
 sg13g2_decap_8 FILLER_110_735 ();
 sg13g2_decap_8 FILLER_110_742 ();
 sg13g2_decap_8 FILLER_110_749 ();
 sg13g2_decap_8 FILLER_110_756 ();
 sg13g2_decap_8 FILLER_110_763 ();
 sg13g2_decap_8 FILLER_110_770 ();
 sg13g2_fill_2 FILLER_110_777 ();
 sg13g2_fill_1 FILLER_110_779 ();
 sg13g2_decap_8 FILLER_110_784 ();
 sg13g2_decap_8 FILLER_110_791 ();
 sg13g2_decap_8 FILLER_110_798 ();
 sg13g2_decap_8 FILLER_110_805 ();
 sg13g2_decap_4 FILLER_110_838 ();
 sg13g2_fill_2 FILLER_110_842 ();
 sg13g2_decap_8 FILLER_110_857 ();
 sg13g2_decap_8 FILLER_110_864 ();
 sg13g2_decap_8 FILLER_110_871 ();
 sg13g2_decap_4 FILLER_110_878 ();
 sg13g2_fill_2 FILLER_110_882 ();
 sg13g2_decap_8 FILLER_110_923 ();
 sg13g2_decap_8 FILLER_110_930 ();
 sg13g2_decap_8 FILLER_110_937 ();
 sg13g2_decap_8 FILLER_110_944 ();
 sg13g2_decap_8 FILLER_110_951 ();
 sg13g2_decap_8 FILLER_110_958 ();
 sg13g2_decap_8 FILLER_110_965 ();
 sg13g2_decap_8 FILLER_110_972 ();
 sg13g2_decap_8 FILLER_110_979 ();
 sg13g2_decap_8 FILLER_110_986 ();
 sg13g2_decap_4 FILLER_110_993 ();
 sg13g2_fill_1 FILLER_110_997 ();
 sg13g2_decap_8 FILLER_110_1013 ();
 sg13g2_decap_8 FILLER_110_1020 ();
 sg13g2_decap_8 FILLER_110_1027 ();
 sg13g2_fill_2 FILLER_110_1034 ();
 sg13g2_fill_1 FILLER_110_1036 ();
 sg13g2_fill_2 FILLER_110_1042 ();
 sg13g2_decap_8 FILLER_110_1053 ();
 sg13g2_decap_8 FILLER_110_1060 ();
 sg13g2_fill_1 FILLER_110_1067 ();
 sg13g2_decap_8 FILLER_110_1102 ();
 sg13g2_decap_4 FILLER_110_1109 ();
 sg13g2_fill_2 FILLER_110_1113 ();
 sg13g2_decap_8 FILLER_110_1124 ();
 sg13g2_decap_4 FILLER_110_1131 ();
 sg13g2_decap_4 FILLER_110_1144 ();
 sg13g2_fill_1 FILLER_110_1148 ();
 sg13g2_decap_8 FILLER_110_1175 ();
 sg13g2_decap_8 FILLER_110_1182 ();
 sg13g2_decap_8 FILLER_110_1189 ();
 sg13g2_decap_8 FILLER_110_1196 ();
 sg13g2_fill_1 FILLER_110_1203 ();
 sg13g2_fill_2 FILLER_110_1210 ();
 sg13g2_decap_8 FILLER_110_1222 ();
 sg13g2_decap_8 FILLER_110_1229 ();
 sg13g2_fill_2 FILLER_110_1236 ();
 sg13g2_fill_1 FILLER_110_1238 ();
 sg13g2_decap_8 FILLER_110_1252 ();
 sg13g2_decap_8 FILLER_110_1259 ();
 sg13g2_decap_8 FILLER_110_1266 ();
 sg13g2_decap_8 FILLER_110_1273 ();
 sg13g2_decap_8 FILLER_110_1280 ();
 sg13g2_decap_8 FILLER_110_1287 ();
 sg13g2_decap_8 FILLER_110_1294 ();
 sg13g2_decap_8 FILLER_110_1301 ();
 sg13g2_decap_8 FILLER_110_1308 ();
 sg13g2_decap_8 FILLER_110_1315 ();
 sg13g2_decap_8 FILLER_110_1322 ();
 sg13g2_decap_8 FILLER_110_1329 ();
 sg13g2_fill_1 FILLER_110_1336 ();
 sg13g2_decap_8 FILLER_110_1345 ();
 sg13g2_decap_8 FILLER_110_1352 ();
 sg13g2_fill_2 FILLER_110_1359 ();
 sg13g2_fill_1 FILLER_110_1361 ();
 sg13g2_decap_8 FILLER_110_1374 ();
 sg13g2_decap_8 FILLER_110_1381 ();
 sg13g2_decap_8 FILLER_110_1388 ();
 sg13g2_decap_8 FILLER_110_1395 ();
 sg13g2_decap_4 FILLER_110_1402 ();
 sg13g2_fill_1 FILLER_110_1406 ();
 sg13g2_fill_2 FILLER_110_1415 ();
 sg13g2_decap_4 FILLER_110_1422 ();
 sg13g2_decap_8 FILLER_110_1438 ();
 sg13g2_decap_8 FILLER_110_1445 ();
 sg13g2_decap_4 FILLER_110_1452 ();
 sg13g2_fill_2 FILLER_110_1456 ();
 sg13g2_fill_2 FILLER_110_1467 ();
 sg13g2_fill_1 FILLER_110_1469 ();
 sg13g2_decap_8 FILLER_110_1483 ();
 sg13g2_decap_8 FILLER_110_1490 ();
 sg13g2_decap_8 FILLER_110_1497 ();
 sg13g2_decap_4 FILLER_110_1504 ();
 sg13g2_fill_1 FILLER_110_1508 ();
 sg13g2_decap_8 FILLER_110_1523 ();
 sg13g2_decap_8 FILLER_110_1530 ();
 sg13g2_decap_8 FILLER_110_1537 ();
 sg13g2_decap_8 FILLER_110_1544 ();
 sg13g2_decap_8 FILLER_110_1551 ();
 sg13g2_fill_2 FILLER_110_1558 ();
 sg13g2_decap_8 FILLER_110_1565 ();
 sg13g2_decap_4 FILLER_110_1572 ();
 sg13g2_fill_1 FILLER_110_1576 ();
 sg13g2_fill_2 FILLER_110_1581 ();
 sg13g2_fill_2 FILLER_110_1592 ();
 sg13g2_fill_1 FILLER_110_1594 ();
 sg13g2_decap_8 FILLER_110_1603 ();
 sg13g2_decap_8 FILLER_110_1610 ();
 sg13g2_decap_8 FILLER_110_1617 ();
 sg13g2_decap_8 FILLER_110_1624 ();
 sg13g2_decap_8 FILLER_110_1631 ();
 sg13g2_decap_8 FILLER_110_1638 ();
 sg13g2_decap_8 FILLER_110_1645 ();
 sg13g2_decap_8 FILLER_110_1652 ();
 sg13g2_decap_8 FILLER_110_1659 ();
 sg13g2_decap_8 FILLER_110_1666 ();
 sg13g2_decap_8 FILLER_110_1673 ();
 sg13g2_fill_2 FILLER_110_1680 ();
 sg13g2_fill_1 FILLER_110_1682 ();
 sg13g2_decap_8 FILLER_110_1691 ();
 sg13g2_decap_8 FILLER_110_1698 ();
 sg13g2_decap_8 FILLER_110_1705 ();
 sg13g2_fill_2 FILLER_110_1712 ();
 sg13g2_fill_1 FILLER_110_1714 ();
 sg13g2_decap_8 FILLER_110_1731 ();
 sg13g2_decap_8 FILLER_110_1738 ();
 sg13g2_decap_8 FILLER_110_1745 ();
 sg13g2_decap_8 FILLER_110_1752 ();
 sg13g2_decap_8 FILLER_110_1759 ();
 sg13g2_fill_2 FILLER_110_1766 ();
 sg13g2_decap_8 FILLER_111_0 ();
 sg13g2_decap_8 FILLER_111_7 ();
 sg13g2_fill_2 FILLER_111_14 ();
 sg13g2_fill_1 FILLER_111_16 ();
 sg13g2_decap_4 FILLER_111_37 ();
 sg13g2_fill_1 FILLER_111_41 ();
 sg13g2_decap_8 FILLER_111_50 ();
 sg13g2_decap_8 FILLER_111_57 ();
 sg13g2_decap_8 FILLER_111_64 ();
 sg13g2_fill_2 FILLER_111_71 ();
 sg13g2_fill_1 FILLER_111_73 ();
 sg13g2_decap_8 FILLER_111_103 ();
 sg13g2_decap_8 FILLER_111_110 ();
 sg13g2_decap_8 FILLER_111_117 ();
 sg13g2_decap_4 FILLER_111_124 ();
 sg13g2_fill_1 FILLER_111_128 ();
 sg13g2_decap_8 FILLER_111_166 ();
 sg13g2_decap_8 FILLER_111_200 ();
 sg13g2_decap_8 FILLER_111_207 ();
 sg13g2_decap_8 FILLER_111_214 ();
 sg13g2_decap_8 FILLER_111_221 ();
 sg13g2_decap_8 FILLER_111_228 ();
 sg13g2_decap_8 FILLER_111_235 ();
 sg13g2_decap_8 FILLER_111_242 ();
 sg13g2_decap_8 FILLER_111_249 ();
 sg13g2_decap_8 FILLER_111_256 ();
 sg13g2_decap_4 FILLER_111_263 ();
 sg13g2_fill_2 FILLER_111_288 ();
 sg13g2_decap_8 FILLER_111_303 ();
 sg13g2_decap_8 FILLER_111_310 ();
 sg13g2_decap_8 FILLER_111_317 ();
 sg13g2_decap_8 FILLER_111_324 ();
 sg13g2_decap_8 FILLER_111_331 ();
 sg13g2_fill_1 FILLER_111_338 ();
 sg13g2_decap_8 FILLER_111_352 ();
 sg13g2_decap_8 FILLER_111_359 ();
 sg13g2_decap_8 FILLER_111_366 ();
 sg13g2_decap_4 FILLER_111_386 ();
 sg13g2_fill_2 FILLER_111_390 ();
 sg13g2_decap_4 FILLER_111_413 ();
 sg13g2_fill_1 FILLER_111_417 ();
 sg13g2_decap_8 FILLER_111_426 ();
 sg13g2_fill_1 FILLER_111_446 ();
 sg13g2_decap_8 FILLER_111_455 ();
 sg13g2_fill_2 FILLER_111_462 ();
 sg13g2_fill_1 FILLER_111_464 ();
 sg13g2_decap_8 FILLER_111_475 ();
 sg13g2_decap_4 FILLER_111_482 ();
 sg13g2_fill_1 FILLER_111_486 ();
 sg13g2_fill_2 FILLER_111_492 ();
 sg13g2_fill_1 FILLER_111_494 ();
 sg13g2_decap_8 FILLER_111_506 ();
 sg13g2_decap_8 FILLER_111_513 ();
 sg13g2_decap_8 FILLER_111_520 ();
 sg13g2_decap_8 FILLER_111_527 ();
 sg13g2_decap_8 FILLER_111_534 ();
 sg13g2_decap_8 FILLER_111_541 ();
 sg13g2_decap_8 FILLER_111_548 ();
 sg13g2_decap_8 FILLER_111_555 ();
 sg13g2_fill_2 FILLER_111_562 ();
 sg13g2_fill_1 FILLER_111_564 ();
 sg13g2_decap_8 FILLER_111_583 ();
 sg13g2_decap_8 FILLER_111_590 ();
 sg13g2_decap_8 FILLER_111_597 ();
 sg13g2_decap_8 FILLER_111_604 ();
 sg13g2_decap_8 FILLER_111_611 ();
 sg13g2_decap_8 FILLER_111_618 ();
 sg13g2_decap_8 FILLER_111_625 ();
 sg13g2_decap_8 FILLER_111_632 ();
 sg13g2_decap_8 FILLER_111_639 ();
 sg13g2_decap_8 FILLER_111_646 ();
 sg13g2_decap_8 FILLER_111_653 ();
 sg13g2_decap_8 FILLER_111_660 ();
 sg13g2_decap_8 FILLER_111_667 ();
 sg13g2_decap_8 FILLER_111_674 ();
 sg13g2_fill_2 FILLER_111_681 ();
 sg13g2_fill_2 FILLER_111_699 ();
 sg13g2_decap_8 FILLER_111_713 ();
 sg13g2_decap_8 FILLER_111_720 ();
 sg13g2_decap_8 FILLER_111_727 ();
 sg13g2_decap_8 FILLER_111_734 ();
 sg13g2_decap_8 FILLER_111_741 ();
 sg13g2_decap_8 FILLER_111_748 ();
 sg13g2_fill_2 FILLER_111_755 ();
 sg13g2_fill_2 FILLER_111_767 ();
 sg13g2_fill_2 FILLER_111_795 ();
 sg13g2_fill_1 FILLER_111_797 ();
 sg13g2_fill_1 FILLER_111_822 ();
 sg13g2_decap_8 FILLER_111_827 ();
 sg13g2_decap_8 FILLER_111_834 ();
 sg13g2_decap_8 FILLER_111_841 ();
 sg13g2_decap_8 FILLER_111_848 ();
 sg13g2_decap_8 FILLER_111_855 ();
 sg13g2_decap_8 FILLER_111_862 ();
 sg13g2_decap_8 FILLER_111_869 ();
 sg13g2_decap_4 FILLER_111_876 ();
 sg13g2_decap_4 FILLER_111_885 ();
 sg13g2_fill_1 FILLER_111_889 ();
 sg13g2_decap_8 FILLER_111_899 ();
 sg13g2_decap_8 FILLER_111_906 ();
 sg13g2_decap_8 FILLER_111_913 ();
 sg13g2_decap_8 FILLER_111_920 ();
 sg13g2_decap_8 FILLER_111_927 ();
 sg13g2_decap_4 FILLER_111_934 ();
 sg13g2_fill_1 FILLER_111_938 ();
 sg13g2_decap_8 FILLER_111_952 ();
 sg13g2_decap_4 FILLER_111_967 ();
 sg13g2_decap_8 FILLER_111_988 ();
 sg13g2_fill_1 FILLER_111_995 ();
 sg13g2_fill_2 FILLER_111_1002 ();
 sg13g2_fill_1 FILLER_111_1030 ();
 sg13g2_decap_8 FILLER_111_1073 ();
 sg13g2_decap_8 FILLER_111_1080 ();
 sg13g2_decap_8 FILLER_111_1087 ();
 sg13g2_decap_8 FILLER_111_1094 ();
 sg13g2_decap_8 FILLER_111_1114 ();
 sg13g2_decap_8 FILLER_111_1121 ();
 sg13g2_fill_2 FILLER_111_1134 ();
 sg13g2_decap_8 FILLER_111_1143 ();
 sg13g2_decap_8 FILLER_111_1150 ();
 sg13g2_fill_2 FILLER_111_1157 ();
 sg13g2_fill_1 FILLER_111_1159 ();
 sg13g2_decap_4 FILLER_111_1164 ();
 sg13g2_fill_2 FILLER_111_1168 ();
 sg13g2_decap_8 FILLER_111_1179 ();
 sg13g2_decap_8 FILLER_111_1186 ();
 sg13g2_decap_8 FILLER_111_1193 ();
 sg13g2_decap_8 FILLER_111_1200 ();
 sg13g2_decap_4 FILLER_111_1207 ();
 sg13g2_decap_8 FILLER_111_1219 ();
 sg13g2_fill_2 FILLER_111_1226 ();
 sg13g2_decap_8 FILLER_111_1241 ();
 sg13g2_decap_8 FILLER_111_1248 ();
 sg13g2_decap_8 FILLER_111_1255 ();
 sg13g2_decap_8 FILLER_111_1262 ();
 sg13g2_decap_8 FILLER_111_1269 ();
 sg13g2_decap_4 FILLER_111_1276 ();
 sg13g2_decap_8 FILLER_111_1288 ();
 sg13g2_decap_8 FILLER_111_1295 ();
 sg13g2_decap_8 FILLER_111_1302 ();
 sg13g2_decap_8 FILLER_111_1309 ();
 sg13g2_decap_8 FILLER_111_1316 ();
 sg13g2_decap_8 FILLER_111_1323 ();
 sg13g2_decap_8 FILLER_111_1330 ();
 sg13g2_decap_8 FILLER_111_1345 ();
 sg13g2_decap_8 FILLER_111_1352 ();
 sg13g2_decap_8 FILLER_111_1359 ();
 sg13g2_decap_8 FILLER_111_1366 ();
 sg13g2_decap_8 FILLER_111_1373 ();
 sg13g2_decap_8 FILLER_111_1380 ();
 sg13g2_decap_8 FILLER_111_1395 ();
 sg13g2_decap_8 FILLER_111_1402 ();
 sg13g2_decap_8 FILLER_111_1409 ();
 sg13g2_decap_8 FILLER_111_1416 ();
 sg13g2_fill_2 FILLER_111_1423 ();
 sg13g2_decap_8 FILLER_111_1430 ();
 sg13g2_decap_8 FILLER_111_1437 ();
 sg13g2_fill_2 FILLER_111_1444 ();
 sg13g2_fill_2 FILLER_111_1458 ();
 sg13g2_fill_2 FILLER_111_1473 ();
 sg13g2_fill_1 FILLER_111_1475 ();
 sg13g2_decap_8 FILLER_111_1486 ();
 sg13g2_fill_2 FILLER_111_1493 ();
 sg13g2_decap_8 FILLER_111_1500 ();
 sg13g2_decap_4 FILLER_111_1507 ();
 sg13g2_decap_8 FILLER_111_1519 ();
 sg13g2_fill_2 FILLER_111_1526 ();
 sg13g2_decap_4 FILLER_111_1536 ();
 sg13g2_fill_1 FILLER_111_1540 ();
 sg13g2_decap_8 FILLER_111_1545 ();
 sg13g2_decap_8 FILLER_111_1552 ();
 sg13g2_decap_4 FILLER_111_1559 ();
 sg13g2_decap_4 FILLER_111_1571 ();
 sg13g2_decap_8 FILLER_111_1591 ();
 sg13g2_decap_8 FILLER_111_1598 ();
 sg13g2_decap_8 FILLER_111_1605 ();
 sg13g2_decap_8 FILLER_111_1612 ();
 sg13g2_decap_4 FILLER_111_1619 ();
 sg13g2_fill_1 FILLER_111_1631 ();
 sg13g2_decap_4 FILLER_111_1637 ();
 sg13g2_fill_1 FILLER_111_1665 ();
 sg13g2_decap_8 FILLER_111_1695 ();
 sg13g2_decap_8 FILLER_111_1702 ();
 sg13g2_decap_8 FILLER_111_1709 ();
 sg13g2_decap_4 FILLER_111_1716 ();
 sg13g2_fill_1 FILLER_111_1720 ();
 sg13g2_decap_8 FILLER_111_1729 ();
 sg13g2_decap_8 FILLER_111_1736 ();
 sg13g2_decap_8 FILLER_111_1743 ();
 sg13g2_decap_8 FILLER_111_1750 ();
 sg13g2_decap_8 FILLER_111_1757 ();
 sg13g2_decap_4 FILLER_111_1764 ();
 sg13g2_decap_8 FILLER_112_0 ();
 sg13g2_decap_8 FILLER_112_7 ();
 sg13g2_decap_8 FILLER_112_14 ();
 sg13g2_fill_2 FILLER_112_21 ();
 sg13g2_decap_8 FILLER_112_40 ();
 sg13g2_decap_8 FILLER_112_47 ();
 sg13g2_fill_2 FILLER_112_54 ();
 sg13g2_fill_1 FILLER_112_56 ();
 sg13g2_fill_2 FILLER_112_65 ();
 sg13g2_fill_1 FILLER_112_67 ();
 sg13g2_decap_8 FILLER_112_103 ();
 sg13g2_decap_8 FILLER_112_110 ();
 sg13g2_decap_8 FILLER_112_117 ();
 sg13g2_decap_4 FILLER_112_124 ();
 sg13g2_fill_2 FILLER_112_128 ();
 sg13g2_fill_2 FILLER_112_146 ();
 sg13g2_decap_8 FILLER_112_153 ();
 sg13g2_decap_8 FILLER_112_160 ();
 sg13g2_decap_8 FILLER_112_167 ();
 sg13g2_decap_4 FILLER_112_174 ();
 sg13g2_decap_8 FILLER_112_196 ();
 sg13g2_decap_8 FILLER_112_203 ();
 sg13g2_decap_8 FILLER_112_210 ();
 sg13g2_decap_4 FILLER_112_217 ();
 sg13g2_fill_1 FILLER_112_221 ();
 sg13g2_fill_2 FILLER_112_227 ();
 sg13g2_decap_8 FILLER_112_233 ();
 sg13g2_decap_8 FILLER_112_240 ();
 sg13g2_decap_8 FILLER_112_247 ();
 sg13g2_decap_8 FILLER_112_254 ();
 sg13g2_decap_8 FILLER_112_261 ();
 sg13g2_fill_1 FILLER_112_268 ();
 sg13g2_decap_8 FILLER_112_282 ();
 sg13g2_decap_8 FILLER_112_289 ();
 sg13g2_decap_8 FILLER_112_296 ();
 sg13g2_decap_8 FILLER_112_303 ();
 sg13g2_decap_8 FILLER_112_310 ();
 sg13g2_decap_8 FILLER_112_317 ();
 sg13g2_fill_2 FILLER_112_324 ();
 sg13g2_decap_8 FILLER_112_339 ();
 sg13g2_decap_8 FILLER_112_346 ();
 sg13g2_decap_8 FILLER_112_362 ();
 sg13g2_decap_8 FILLER_112_369 ();
 sg13g2_decap_8 FILLER_112_376 ();
 sg13g2_decap_8 FILLER_112_383 ();
 sg13g2_decap_4 FILLER_112_390 ();
 sg13g2_fill_2 FILLER_112_394 ();
 sg13g2_decap_8 FILLER_112_409 ();
 sg13g2_decap_8 FILLER_112_416 ();
 sg13g2_decap_8 FILLER_112_423 ();
 sg13g2_decap_8 FILLER_112_430 ();
 sg13g2_decap_4 FILLER_112_437 ();
 sg13g2_decap_8 FILLER_112_454 ();
 sg13g2_decap_8 FILLER_112_461 ();
 sg13g2_decap_8 FILLER_112_468 ();
 sg13g2_decap_8 FILLER_112_475 ();
 sg13g2_decap_4 FILLER_112_482 ();
 sg13g2_fill_1 FILLER_112_486 ();
 sg13g2_decap_8 FILLER_112_495 ();
 sg13g2_decap_8 FILLER_112_502 ();
 sg13g2_decap_8 FILLER_112_509 ();
 sg13g2_decap_8 FILLER_112_516 ();
 sg13g2_decap_8 FILLER_112_523 ();
 sg13g2_decap_8 FILLER_112_530 ();
 sg13g2_decap_8 FILLER_112_537 ();
 sg13g2_decap_8 FILLER_112_544 ();
 sg13g2_decap_8 FILLER_112_551 ();
 sg13g2_decap_4 FILLER_112_558 ();
 sg13g2_fill_1 FILLER_112_562 ();
 sg13g2_decap_8 FILLER_112_579 ();
 sg13g2_decap_8 FILLER_112_586 ();
 sg13g2_decap_8 FILLER_112_593 ();
 sg13g2_decap_8 FILLER_112_600 ();
 sg13g2_decap_8 FILLER_112_607 ();
 sg13g2_decap_8 FILLER_112_614 ();
 sg13g2_decap_8 FILLER_112_621 ();
 sg13g2_decap_4 FILLER_112_628 ();
 sg13g2_fill_2 FILLER_112_632 ();
 sg13g2_decap_4 FILLER_112_650 ();
 sg13g2_fill_1 FILLER_112_654 ();
 sg13g2_decap_8 FILLER_112_664 ();
 sg13g2_decap_8 FILLER_112_671 ();
 sg13g2_decap_4 FILLER_112_678 ();
 sg13g2_fill_1 FILLER_112_682 ();
 sg13g2_decap_8 FILLER_112_687 ();
 sg13g2_decap_8 FILLER_112_694 ();
 sg13g2_fill_1 FILLER_112_701 ();
 sg13g2_decap_8 FILLER_112_718 ();
 sg13g2_decap_8 FILLER_112_725 ();
 sg13g2_decap_4 FILLER_112_732 ();
 sg13g2_decap_8 FILLER_112_740 ();
 sg13g2_fill_1 FILLER_112_747 ();
 sg13g2_decap_8 FILLER_112_753 ();
 sg13g2_decap_8 FILLER_112_760 ();
 sg13g2_decap_8 FILLER_112_767 ();
 sg13g2_decap_8 FILLER_112_774 ();
 sg13g2_decap_4 FILLER_112_781 ();
 sg13g2_fill_2 FILLER_112_785 ();
 sg13g2_fill_1 FILLER_112_818 ();
 sg13g2_decap_8 FILLER_112_834 ();
 sg13g2_decap_8 FILLER_112_841 ();
 sg13g2_decap_8 FILLER_112_848 ();
 sg13g2_decap_8 FILLER_112_855 ();
 sg13g2_decap_8 FILLER_112_862 ();
 sg13g2_decap_4 FILLER_112_869 ();
 sg13g2_decap_8 FILLER_112_908 ();
 sg13g2_decap_8 FILLER_112_915 ();
 sg13g2_decap_8 FILLER_112_922 ();
 sg13g2_decap_8 FILLER_112_929 ();
 sg13g2_fill_2 FILLER_112_936 ();
 sg13g2_decap_8 FILLER_112_951 ();
 sg13g2_fill_2 FILLER_112_958 ();
 sg13g2_decap_4 FILLER_112_964 ();
 sg13g2_fill_1 FILLER_112_968 ();
 sg13g2_decap_8 FILLER_112_995 ();
 sg13g2_fill_2 FILLER_112_1002 ();
 sg13g2_decap_8 FILLER_112_1010 ();
 sg13g2_decap_8 FILLER_112_1017 ();
 sg13g2_decap_8 FILLER_112_1024 ();
 sg13g2_decap_8 FILLER_112_1031 ();
 sg13g2_fill_1 FILLER_112_1038 ();
 sg13g2_fill_1 FILLER_112_1044 ();
 sg13g2_decap_8 FILLER_112_1052 ();
 sg13g2_fill_1 FILLER_112_1059 ();
 sg13g2_decap_8 FILLER_112_1069 ();
 sg13g2_decap_8 FILLER_112_1076 ();
 sg13g2_decap_8 FILLER_112_1083 ();
 sg13g2_decap_8 FILLER_112_1090 ();
 sg13g2_decap_8 FILLER_112_1097 ();
 sg13g2_decap_4 FILLER_112_1104 ();
 sg13g2_fill_2 FILLER_112_1117 ();
 sg13g2_decap_8 FILLER_112_1143 ();
 sg13g2_decap_8 FILLER_112_1150 ();
 sg13g2_decap_8 FILLER_112_1157 ();
 sg13g2_decap_8 FILLER_112_1164 ();
 sg13g2_fill_2 FILLER_112_1171 ();
 sg13g2_decap_8 FILLER_112_1204 ();
 sg13g2_decap_8 FILLER_112_1211 ();
 sg13g2_decap_8 FILLER_112_1218 ();
 sg13g2_decap_8 FILLER_112_1225 ();
 sg13g2_decap_8 FILLER_112_1245 ();
 sg13g2_decap_4 FILLER_112_1252 ();
 sg13g2_fill_2 FILLER_112_1256 ();
 sg13g2_decap_8 FILLER_112_1266 ();
 sg13g2_decap_8 FILLER_112_1273 ();
 sg13g2_decap_8 FILLER_112_1280 ();
 sg13g2_decap_8 FILLER_112_1287 ();
 sg13g2_decap_8 FILLER_112_1294 ();
 sg13g2_fill_2 FILLER_112_1311 ();
 sg13g2_decap_8 FILLER_112_1327 ();
 sg13g2_decap_8 FILLER_112_1334 ();
 sg13g2_decap_8 FILLER_112_1341 ();
 sg13g2_fill_2 FILLER_112_1348 ();
 sg13g2_fill_1 FILLER_112_1350 ();
 sg13g2_decap_4 FILLER_112_1359 ();
 sg13g2_decap_4 FILLER_112_1379 ();
 sg13g2_fill_1 FILLER_112_1383 ();
 sg13g2_decap_8 FILLER_112_1392 ();
 sg13g2_decap_4 FILLER_112_1399 ();
 sg13g2_fill_1 FILLER_112_1411 ();
 sg13g2_decap_8 FILLER_112_1420 ();
 sg13g2_decap_8 FILLER_112_1427 ();
 sg13g2_decap_8 FILLER_112_1434 ();
 sg13g2_decap_8 FILLER_112_1441 ();
 sg13g2_decap_4 FILLER_112_1448 ();
 sg13g2_decap_8 FILLER_112_1474 ();
 sg13g2_decap_8 FILLER_112_1481 ();
 sg13g2_decap_8 FILLER_112_1488 ();
 sg13g2_fill_2 FILLER_112_1495 ();
 sg13g2_decap_8 FILLER_112_1513 ();
 sg13g2_decap_8 FILLER_112_1520 ();
 sg13g2_decap_8 FILLER_112_1527 ();
 sg13g2_decap_8 FILLER_112_1534 ();
 sg13g2_decap_8 FILLER_112_1541 ();
 sg13g2_decap_8 FILLER_112_1548 ();
 sg13g2_decap_8 FILLER_112_1555 ();
 sg13g2_decap_8 FILLER_112_1562 ();
 sg13g2_decap_4 FILLER_112_1569 ();
 sg13g2_fill_1 FILLER_112_1573 ();
 sg13g2_fill_1 FILLER_112_1582 ();
 sg13g2_decap_8 FILLER_112_1591 ();
 sg13g2_decap_8 FILLER_112_1598 ();
 sg13g2_decap_8 FILLER_112_1605 ();
 sg13g2_decap_8 FILLER_112_1612 ();
 sg13g2_decap_4 FILLER_112_1619 ();
 sg13g2_decap_8 FILLER_112_1644 ();
 sg13g2_decap_8 FILLER_112_1659 ();
 sg13g2_decap_8 FILLER_112_1666 ();
 sg13g2_decap_8 FILLER_112_1673 ();
 sg13g2_fill_1 FILLER_112_1680 ();
 sg13g2_decap_8 FILLER_112_1685 ();
 sg13g2_decap_8 FILLER_112_1692 ();
 sg13g2_decap_8 FILLER_112_1699 ();
 sg13g2_fill_2 FILLER_112_1710 ();
 sg13g2_fill_1 FILLER_112_1712 ();
 sg13g2_decap_8 FILLER_112_1720 ();
 sg13g2_decap_8 FILLER_112_1727 ();
 sg13g2_decap_4 FILLER_112_1734 ();
 sg13g2_fill_2 FILLER_112_1738 ();
 sg13g2_decap_8 FILLER_112_1751 ();
 sg13g2_decap_8 FILLER_112_1758 ();
 sg13g2_fill_2 FILLER_112_1765 ();
 sg13g2_fill_1 FILLER_112_1767 ();
 sg13g2_decap_8 FILLER_113_0 ();
 sg13g2_decap_8 FILLER_113_7 ();
 sg13g2_decap_8 FILLER_113_14 ();
 sg13g2_fill_2 FILLER_113_21 ();
 sg13g2_fill_1 FILLER_113_23 ();
 sg13g2_decap_8 FILLER_113_28 ();
 sg13g2_decap_8 FILLER_113_35 ();
 sg13g2_decap_8 FILLER_113_42 ();
 sg13g2_decap_4 FILLER_113_49 ();
 sg13g2_decap_8 FILLER_113_77 ();
 sg13g2_decap_8 FILLER_113_84 ();
 sg13g2_fill_1 FILLER_113_91 ();
 sg13g2_decap_8 FILLER_113_96 ();
 sg13g2_decap_8 FILLER_113_103 ();
 sg13g2_decap_8 FILLER_113_110 ();
 sg13g2_decap_4 FILLER_113_117 ();
 sg13g2_fill_1 FILLER_113_121 ();
 sg13g2_decap_8 FILLER_113_126 ();
 sg13g2_decap_4 FILLER_113_133 ();
 sg13g2_fill_1 FILLER_113_137 ();
 sg13g2_decap_8 FILLER_113_149 ();
 sg13g2_decap_8 FILLER_113_156 ();
 sg13g2_decap_8 FILLER_113_163 ();
 sg13g2_decap_8 FILLER_113_170 ();
 sg13g2_decap_8 FILLER_113_177 ();
 sg13g2_decap_8 FILLER_113_184 ();
 sg13g2_decap_8 FILLER_113_191 ();
 sg13g2_decap_8 FILLER_113_198 ();
 sg13g2_decap_8 FILLER_113_205 ();
 sg13g2_decap_8 FILLER_113_212 ();
 sg13g2_fill_2 FILLER_113_219 ();
 sg13g2_decap_8 FILLER_113_241 ();
 sg13g2_decap_8 FILLER_113_248 ();
 sg13g2_decap_4 FILLER_113_255 ();
 sg13g2_fill_1 FILLER_113_259 ();
 sg13g2_decap_8 FILLER_113_268 ();
 sg13g2_decap_8 FILLER_113_275 ();
 sg13g2_decap_8 FILLER_113_282 ();
 sg13g2_decap_8 FILLER_113_289 ();
 sg13g2_decap_8 FILLER_113_296 ();
 sg13g2_decap_8 FILLER_113_303 ();
 sg13g2_decap_8 FILLER_113_310 ();
 sg13g2_fill_2 FILLER_113_317 ();
 sg13g2_fill_1 FILLER_113_319 ();
 sg13g2_fill_1 FILLER_113_333 ();
 sg13g2_decap_8 FILLER_113_360 ();
 sg13g2_decap_8 FILLER_113_367 ();
 sg13g2_decap_8 FILLER_113_374 ();
 sg13g2_decap_8 FILLER_113_381 ();
 sg13g2_decap_8 FILLER_113_388 ();
 sg13g2_decap_8 FILLER_113_395 ();
 sg13g2_decap_8 FILLER_113_402 ();
 sg13g2_decap_4 FILLER_113_409 ();
 sg13g2_decap_8 FILLER_113_421 ();
 sg13g2_decap_4 FILLER_113_428 ();
 sg13g2_decap_8 FILLER_113_447 ();
 sg13g2_decap_4 FILLER_113_454 ();
 sg13g2_fill_2 FILLER_113_458 ();
 sg13g2_decap_8 FILLER_113_463 ();
 sg13g2_decap_8 FILLER_113_470 ();
 sg13g2_decap_8 FILLER_113_477 ();
 sg13g2_decap_8 FILLER_113_484 ();
 sg13g2_decap_8 FILLER_113_491 ();
 sg13g2_decap_8 FILLER_113_498 ();
 sg13g2_fill_1 FILLER_113_505 ();
 sg13g2_decap_8 FILLER_113_516 ();
 sg13g2_decap_8 FILLER_113_523 ();
 sg13g2_decap_4 FILLER_113_530 ();
 sg13g2_fill_2 FILLER_113_534 ();
 sg13g2_decap_8 FILLER_113_556 ();
 sg13g2_decap_8 FILLER_113_563 ();
 sg13g2_decap_8 FILLER_113_570 ();
 sg13g2_decap_8 FILLER_113_577 ();
 sg13g2_decap_8 FILLER_113_584 ();
 sg13g2_decap_8 FILLER_113_591 ();
 sg13g2_decap_8 FILLER_113_598 ();
 sg13g2_decap_8 FILLER_113_605 ();
 sg13g2_fill_2 FILLER_113_612 ();
 sg13g2_fill_1 FILLER_113_614 ();
 sg13g2_decap_8 FILLER_113_619 ();
 sg13g2_decap_8 FILLER_113_626 ();
 sg13g2_decap_8 FILLER_113_642 ();
 sg13g2_fill_2 FILLER_113_649 ();
 sg13g2_decap_8 FILLER_113_669 ();
 sg13g2_decap_8 FILLER_113_676 ();
 sg13g2_decap_8 FILLER_113_683 ();
 sg13g2_decap_4 FILLER_113_690 ();
 sg13g2_fill_2 FILLER_113_694 ();
 sg13g2_decap_8 FILLER_113_728 ();
 sg13g2_fill_1 FILLER_113_735 ();
 sg13g2_decap_8 FILLER_113_767 ();
 sg13g2_decap_8 FILLER_113_774 ();
 sg13g2_decap_8 FILLER_113_781 ();
 sg13g2_fill_2 FILLER_113_788 ();
 sg13g2_fill_1 FILLER_113_790 ();
 sg13g2_fill_1 FILLER_113_800 ();
 sg13g2_decap_8 FILLER_113_805 ();
 sg13g2_decap_8 FILLER_113_812 ();
 sg13g2_decap_8 FILLER_113_819 ();
 sg13g2_decap_4 FILLER_113_826 ();
 sg13g2_decap_8 FILLER_113_851 ();
 sg13g2_decap_8 FILLER_113_858 ();
 sg13g2_decap_4 FILLER_113_865 ();
 sg13g2_fill_1 FILLER_113_882 ();
 sg13g2_decap_8 FILLER_113_891 ();
 sg13g2_fill_1 FILLER_113_898 ();
 sg13g2_decap_8 FILLER_113_912 ();
 sg13g2_decap_8 FILLER_113_919 ();
 sg13g2_decap_8 FILLER_113_926 ();
 sg13g2_decap_8 FILLER_113_933 ();
 sg13g2_decap_8 FILLER_113_940 ();
 sg13g2_decap_8 FILLER_113_947 ();
 sg13g2_decap_8 FILLER_113_954 ();
 sg13g2_decap_8 FILLER_113_965 ();
 sg13g2_decap_4 FILLER_113_972 ();
 sg13g2_fill_2 FILLER_113_976 ();
 sg13g2_fill_2 FILLER_113_986 ();
 sg13g2_fill_1 FILLER_113_988 ();
 sg13g2_decap_8 FILLER_113_1024 ();
 sg13g2_decap_8 FILLER_113_1031 ();
 sg13g2_decap_4 FILLER_113_1038 ();
 sg13g2_fill_1 FILLER_113_1042 ();
 sg13g2_decap_8 FILLER_113_1064 ();
 sg13g2_decap_8 FILLER_113_1071 ();
 sg13g2_decap_8 FILLER_113_1078 ();
 sg13g2_decap_8 FILLER_113_1085 ();
 sg13g2_fill_2 FILLER_113_1092 ();
 sg13g2_fill_1 FILLER_113_1094 ();
 sg13g2_decap_8 FILLER_113_1101 ();
 sg13g2_decap_8 FILLER_113_1116 ();
 sg13g2_decap_4 FILLER_113_1123 ();
 sg13g2_fill_1 FILLER_113_1127 ();
 sg13g2_decap_4 FILLER_113_1137 ();
 sg13g2_fill_1 FILLER_113_1141 ();
 sg13g2_decap_8 FILLER_113_1148 ();
 sg13g2_decap_8 FILLER_113_1155 ();
 sg13g2_decap_8 FILLER_113_1162 ();
 sg13g2_decap_8 FILLER_113_1169 ();
 sg13g2_decap_8 FILLER_113_1176 ();
 sg13g2_fill_1 FILLER_113_1183 ();
 sg13g2_decap_8 FILLER_113_1188 ();
 sg13g2_decap_8 FILLER_113_1208 ();
 sg13g2_decap_8 FILLER_113_1215 ();
 sg13g2_fill_2 FILLER_113_1222 ();
 sg13g2_fill_1 FILLER_113_1224 ();
 sg13g2_decap_8 FILLER_113_1233 ();
 sg13g2_decap_8 FILLER_113_1240 ();
 sg13g2_fill_1 FILLER_113_1247 ();
 sg13g2_fill_2 FILLER_113_1277 ();
 sg13g2_fill_1 FILLER_113_1279 ();
 sg13g2_decap_8 FILLER_113_1329 ();
 sg13g2_decap_8 FILLER_113_1336 ();
 sg13g2_decap_8 FILLER_113_1343 ();
 sg13g2_decap_8 FILLER_113_1350 ();
 sg13g2_decap_8 FILLER_113_1357 ();
 sg13g2_decap_8 FILLER_113_1364 ();
 sg13g2_fill_2 FILLER_113_1371 ();
 sg13g2_fill_1 FILLER_113_1373 ();
 sg13g2_fill_2 FILLER_113_1396 ();
 sg13g2_fill_1 FILLER_113_1398 ();
 sg13g2_decap_8 FILLER_113_1403 ();
 sg13g2_decap_8 FILLER_113_1410 ();
 sg13g2_decap_8 FILLER_113_1417 ();
 sg13g2_decap_8 FILLER_113_1424 ();
 sg13g2_decap_8 FILLER_113_1431 ();
 sg13g2_decap_8 FILLER_113_1438 ();
 sg13g2_decap_8 FILLER_113_1445 ();
 sg13g2_decap_8 FILLER_113_1452 ();
 sg13g2_decap_8 FILLER_113_1459 ();
 sg13g2_decap_8 FILLER_113_1466 ();
 sg13g2_decap_8 FILLER_113_1473 ();
 sg13g2_decap_8 FILLER_113_1480 ();
 sg13g2_decap_8 FILLER_113_1487 ();
 sg13g2_decap_4 FILLER_113_1494 ();
 sg13g2_fill_1 FILLER_113_1498 ();
 sg13g2_decap_8 FILLER_113_1512 ();
 sg13g2_decap_8 FILLER_113_1519 ();
 sg13g2_decap_8 FILLER_113_1526 ();
 sg13g2_decap_4 FILLER_113_1533 ();
 sg13g2_fill_2 FILLER_113_1537 ();
 sg13g2_fill_2 FILLER_113_1543 ();
 sg13g2_decap_8 FILLER_113_1551 ();
 sg13g2_decap_8 FILLER_113_1558 ();
 sg13g2_decap_8 FILLER_113_1565 ();
 sg13g2_decap_8 FILLER_113_1572 ();
 sg13g2_decap_8 FILLER_113_1579 ();
 sg13g2_decap_8 FILLER_113_1586 ();
 sg13g2_decap_4 FILLER_113_1593 ();
 sg13g2_decap_8 FILLER_113_1604 ();
 sg13g2_decap_8 FILLER_113_1611 ();
 sg13g2_decap_8 FILLER_113_1618 ();
 sg13g2_decap_4 FILLER_113_1625 ();
 sg13g2_fill_1 FILLER_113_1629 ();
 sg13g2_fill_2 FILLER_113_1634 ();
 sg13g2_decap_8 FILLER_113_1648 ();
 sg13g2_decap_8 FILLER_113_1655 ();
 sg13g2_decap_8 FILLER_113_1662 ();
 sg13g2_decap_8 FILLER_113_1669 ();
 sg13g2_decap_8 FILLER_113_1676 ();
 sg13g2_decap_8 FILLER_113_1683 ();
 sg13g2_decap_4 FILLER_113_1690 ();
 sg13g2_fill_2 FILLER_113_1694 ();
 sg13g2_decap_8 FILLER_113_1713 ();
 sg13g2_fill_1 FILLER_113_1720 ();
 sg13g2_fill_1 FILLER_113_1734 ();
 sg13g2_decap_8 FILLER_113_1759 ();
 sg13g2_fill_2 FILLER_113_1766 ();
 sg13g2_decap_8 FILLER_114_0 ();
 sg13g2_decap_8 FILLER_114_7 ();
 sg13g2_decap_4 FILLER_114_14 ();
 sg13g2_fill_2 FILLER_114_18 ();
 sg13g2_decap_8 FILLER_114_36 ();
 sg13g2_decap_4 FILLER_114_43 ();
 sg13g2_fill_1 FILLER_114_47 ();
 sg13g2_decap_8 FILLER_114_56 ();
 sg13g2_decap_8 FILLER_114_63 ();
 sg13g2_decap_8 FILLER_114_78 ();
 sg13g2_decap_8 FILLER_114_85 ();
 sg13g2_decap_8 FILLER_114_92 ();
 sg13g2_decap_8 FILLER_114_99 ();
 sg13g2_decap_8 FILLER_114_106 ();
 sg13g2_fill_2 FILLER_114_113 ();
 sg13g2_fill_1 FILLER_114_115 ();
 sg13g2_fill_1 FILLER_114_128 ();
 sg13g2_decap_8 FILLER_114_134 ();
 sg13g2_decap_8 FILLER_114_141 ();
 sg13g2_decap_8 FILLER_114_148 ();
 sg13g2_decap_8 FILLER_114_155 ();
 sg13g2_fill_1 FILLER_114_167 ();
 sg13g2_decap_8 FILLER_114_172 ();
 sg13g2_fill_2 FILLER_114_179 ();
 sg13g2_fill_1 FILLER_114_181 ();
 sg13g2_decap_8 FILLER_114_187 ();
 sg13g2_decap_8 FILLER_114_194 ();
 sg13g2_decap_8 FILLER_114_201 ();
 sg13g2_decap_4 FILLER_114_208 ();
 sg13g2_fill_1 FILLER_114_212 ();
 sg13g2_decap_8 FILLER_114_231 ();
 sg13g2_decap_8 FILLER_114_238 ();
 sg13g2_decap_8 FILLER_114_245 ();
 sg13g2_decap_8 FILLER_114_252 ();
 sg13g2_decap_8 FILLER_114_259 ();
 sg13g2_decap_8 FILLER_114_266 ();
 sg13g2_decap_4 FILLER_114_273 ();
 sg13g2_fill_2 FILLER_114_277 ();
 sg13g2_decap_8 FILLER_114_287 ();
 sg13g2_decap_8 FILLER_114_294 ();
 sg13g2_decap_8 FILLER_114_301 ();
 sg13g2_decap_8 FILLER_114_308 ();
 sg13g2_decap_8 FILLER_114_315 ();
 sg13g2_decap_8 FILLER_114_322 ();
 sg13g2_fill_2 FILLER_114_337 ();
 sg13g2_fill_1 FILLER_114_339 ();
 sg13g2_decap_8 FILLER_114_359 ();
 sg13g2_decap_8 FILLER_114_366 ();
 sg13g2_decap_8 FILLER_114_373 ();
 sg13g2_decap_8 FILLER_114_380 ();
 sg13g2_decap_8 FILLER_114_387 ();
 sg13g2_fill_1 FILLER_114_394 ();
 sg13g2_decap_8 FILLER_114_404 ();
 sg13g2_decap_8 FILLER_114_411 ();
 sg13g2_decap_8 FILLER_114_418 ();
 sg13g2_decap_8 FILLER_114_425 ();
 sg13g2_decap_8 FILLER_114_432 ();
 sg13g2_decap_8 FILLER_114_439 ();
 sg13g2_decap_8 FILLER_114_446 ();
 sg13g2_decap_8 FILLER_114_453 ();
 sg13g2_decap_8 FILLER_114_465 ();
 sg13g2_decap_8 FILLER_114_472 ();
 sg13g2_decap_8 FILLER_114_479 ();
 sg13g2_decap_8 FILLER_114_486 ();
 sg13g2_fill_2 FILLER_114_493 ();
 sg13g2_fill_1 FILLER_114_495 ();
 sg13g2_decap_8 FILLER_114_514 ();
 sg13g2_decap_8 FILLER_114_521 ();
 sg13g2_decap_4 FILLER_114_528 ();
 sg13g2_decap_8 FILLER_114_558 ();
 sg13g2_decap_8 FILLER_114_565 ();
 sg13g2_decap_8 FILLER_114_572 ();
 sg13g2_decap_8 FILLER_114_579 ();
 sg13g2_decap_8 FILLER_114_586 ();
 sg13g2_decap_8 FILLER_114_593 ();
 sg13g2_decap_4 FILLER_114_600 ();
 sg13g2_decap_4 FILLER_114_630 ();
 sg13g2_fill_2 FILLER_114_634 ();
 sg13g2_decap_4 FILLER_114_649 ();
 sg13g2_fill_1 FILLER_114_653 ();
 sg13g2_decap_8 FILLER_114_659 ();
 sg13g2_decap_8 FILLER_114_674 ();
 sg13g2_decap_8 FILLER_114_681 ();
 sg13g2_decap_8 FILLER_114_688 ();
 sg13g2_decap_8 FILLER_114_695 ();
 sg13g2_fill_2 FILLER_114_702 ();
 sg13g2_fill_1 FILLER_114_704 ();
 sg13g2_fill_2 FILLER_114_710 ();
 sg13g2_fill_1 FILLER_114_712 ();
 sg13g2_decap_8 FILLER_114_721 ();
 sg13g2_decap_8 FILLER_114_728 ();
 sg13g2_decap_8 FILLER_114_735 ();
 sg13g2_decap_8 FILLER_114_742 ();
 sg13g2_decap_4 FILLER_114_749 ();
 sg13g2_fill_1 FILLER_114_753 ();
 sg13g2_decap_8 FILLER_114_772 ();
 sg13g2_decap_8 FILLER_114_779 ();
 sg13g2_decap_4 FILLER_114_786 ();
 sg13g2_fill_2 FILLER_114_790 ();
 sg13g2_decap_8 FILLER_114_818 ();
 sg13g2_decap_8 FILLER_114_825 ();
 sg13g2_decap_8 FILLER_114_832 ();
 sg13g2_decap_4 FILLER_114_839 ();
 sg13g2_fill_2 FILLER_114_843 ();
 sg13g2_decap_8 FILLER_114_858 ();
 sg13g2_decap_8 FILLER_114_865 ();
 sg13g2_decap_8 FILLER_114_872 ();
 sg13g2_decap_8 FILLER_114_879 ();
 sg13g2_decap_8 FILLER_114_886 ();
 sg13g2_decap_8 FILLER_114_893 ();
 sg13g2_decap_8 FILLER_114_900 ();
 sg13g2_fill_1 FILLER_114_907 ();
 sg13g2_decap_8 FILLER_114_923 ();
 sg13g2_decap_8 FILLER_114_930 ();
 sg13g2_decap_8 FILLER_114_937 ();
 sg13g2_decap_4 FILLER_114_944 ();
 sg13g2_fill_1 FILLER_114_948 ();
 sg13g2_decap_8 FILLER_114_960 ();
 sg13g2_decap_8 FILLER_114_967 ();
 sg13g2_decap_8 FILLER_114_974 ();
 sg13g2_decap_8 FILLER_114_981 ();
 sg13g2_decap_8 FILLER_114_988 ();
 sg13g2_decap_8 FILLER_114_995 ();
 sg13g2_fill_1 FILLER_114_1002 ();
 sg13g2_fill_1 FILLER_114_1008 ();
 sg13g2_decap_8 FILLER_114_1013 ();
 sg13g2_decap_8 FILLER_114_1020 ();
 sg13g2_decap_8 FILLER_114_1027 ();
 sg13g2_decap_8 FILLER_114_1034 ();
 sg13g2_decap_8 FILLER_114_1041 ();
 sg13g2_decap_8 FILLER_114_1048 ();
 sg13g2_decap_8 FILLER_114_1055 ();
 sg13g2_decap_8 FILLER_114_1062 ();
 sg13g2_fill_2 FILLER_114_1069 ();
 sg13g2_decap_8 FILLER_114_1075 ();
 sg13g2_decap_4 FILLER_114_1082 ();
 sg13g2_decap_8 FILLER_114_1112 ();
 sg13g2_decap_8 FILLER_114_1119 ();
 sg13g2_fill_2 FILLER_114_1126 ();
 sg13g2_fill_1 FILLER_114_1128 ();
 sg13g2_decap_8 FILLER_114_1155 ();
 sg13g2_decap_8 FILLER_114_1162 ();
 sg13g2_decap_8 FILLER_114_1169 ();
 sg13g2_decap_8 FILLER_114_1176 ();
 sg13g2_decap_4 FILLER_114_1195 ();
 sg13g2_decap_8 FILLER_114_1207 ();
 sg13g2_decap_8 FILLER_114_1214 ();
 sg13g2_decap_8 FILLER_114_1221 ();
 sg13g2_decap_8 FILLER_114_1228 ();
 sg13g2_decap_8 FILLER_114_1235 ();
 sg13g2_decap_4 FILLER_114_1242 ();
 sg13g2_fill_1 FILLER_114_1246 ();
 sg13g2_fill_1 FILLER_114_1255 ();
 sg13g2_decap_8 FILLER_114_1260 ();
 sg13g2_decap_4 FILLER_114_1267 ();
 sg13g2_decap_8 FILLER_114_1284 ();
 sg13g2_fill_1 FILLER_114_1291 ();
 sg13g2_decap_8 FILLER_114_1322 ();
 sg13g2_decap_8 FILLER_114_1329 ();
 sg13g2_decap_8 FILLER_114_1336 ();
 sg13g2_decap_4 FILLER_114_1343 ();
 sg13g2_fill_1 FILLER_114_1347 ();
 sg13g2_decap_8 FILLER_114_1356 ();
 sg13g2_decap_8 FILLER_114_1363 ();
 sg13g2_decap_8 FILLER_114_1370 ();
 sg13g2_fill_2 FILLER_114_1377 ();
 sg13g2_fill_1 FILLER_114_1387 ();
 sg13g2_decap_4 FILLER_114_1401 ();
 sg13g2_fill_1 FILLER_114_1405 ();
 sg13g2_decap_8 FILLER_114_1412 ();
 sg13g2_fill_1 FILLER_114_1419 ();
 sg13g2_decap_8 FILLER_114_1445 ();
 sg13g2_decap_8 FILLER_114_1452 ();
 sg13g2_decap_8 FILLER_114_1459 ();
 sg13g2_decap_8 FILLER_114_1466 ();
 sg13g2_decap_8 FILLER_114_1473 ();
 sg13g2_decap_4 FILLER_114_1480 ();
 sg13g2_fill_2 FILLER_114_1484 ();
 sg13g2_decap_8 FILLER_114_1503 ();
 sg13g2_decap_8 FILLER_114_1510 ();
 sg13g2_decap_4 FILLER_114_1517 ();
 sg13g2_fill_2 FILLER_114_1521 ();
 sg13g2_decap_4 FILLER_114_1529 ();
 sg13g2_decap_8 FILLER_114_1554 ();
 sg13g2_decap_8 FILLER_114_1561 ();
 sg13g2_decap_8 FILLER_114_1568 ();
 sg13g2_decap_8 FILLER_114_1575 ();
 sg13g2_decap_8 FILLER_114_1582 ();
 sg13g2_fill_2 FILLER_114_1589 ();
 sg13g2_decap_8 FILLER_114_1610 ();
 sg13g2_decap_8 FILLER_114_1617 ();
 sg13g2_decap_8 FILLER_114_1624 ();
 sg13g2_decap_8 FILLER_114_1631 ();
 sg13g2_decap_8 FILLER_114_1638 ();
 sg13g2_decap_8 FILLER_114_1645 ();
 sg13g2_decap_8 FILLER_114_1652 ();
 sg13g2_decap_4 FILLER_114_1659 ();
 sg13g2_fill_1 FILLER_114_1663 ();
 sg13g2_decap_8 FILLER_114_1669 ();
 sg13g2_decap_4 FILLER_114_1676 ();
 sg13g2_fill_1 FILLER_114_1680 ();
 sg13g2_decap_8 FILLER_114_1689 ();
 sg13g2_decap_8 FILLER_114_1696 ();
 sg13g2_decap_4 FILLER_114_1703 ();
 sg13g2_fill_1 FILLER_114_1707 ();
 sg13g2_decap_8 FILLER_114_1716 ();
 sg13g2_decap_4 FILLER_114_1723 ();
 sg13g2_decap_8 FILLER_114_1739 ();
 sg13g2_decap_8 FILLER_114_1746 ();
 sg13g2_decap_8 FILLER_114_1753 ();
 sg13g2_decap_8 FILLER_114_1760 ();
 sg13g2_fill_1 FILLER_114_1767 ();
 sg13g2_decap_8 FILLER_115_0 ();
 sg13g2_decap_8 FILLER_115_7 ();
 sg13g2_decap_4 FILLER_115_14 ();
 sg13g2_fill_2 FILLER_115_18 ();
 sg13g2_decap_8 FILLER_115_37 ();
 sg13g2_decap_8 FILLER_115_44 ();
 sg13g2_decap_8 FILLER_115_51 ();
 sg13g2_decap_8 FILLER_115_58 ();
 sg13g2_decap_8 FILLER_115_65 ();
 sg13g2_decap_8 FILLER_115_72 ();
 sg13g2_decap_4 FILLER_115_79 ();
 sg13g2_fill_2 FILLER_115_83 ();
 sg13g2_decap_8 FILLER_115_102 ();
 sg13g2_fill_2 FILLER_115_109 ();
 sg13g2_fill_1 FILLER_115_111 ();
 sg13g2_decap_8 FILLER_115_136 ();
 sg13g2_decap_8 FILLER_115_143 ();
 sg13g2_decap_8 FILLER_115_150 ();
 sg13g2_fill_2 FILLER_115_157 ();
 sg13g2_fill_2 FILLER_115_168 ();
 sg13g2_fill_1 FILLER_115_170 ();
 sg13g2_fill_1 FILLER_115_187 ();
 sg13g2_decap_4 FILLER_115_196 ();
 sg13g2_fill_2 FILLER_115_200 ();
 sg13g2_decap_8 FILLER_115_228 ();
 sg13g2_decap_8 FILLER_115_235 ();
 sg13g2_decap_4 FILLER_115_242 ();
 sg13g2_fill_2 FILLER_115_246 ();
 sg13g2_fill_2 FILLER_115_256 ();
 sg13g2_decap_4 FILLER_115_270 ();
 sg13g2_fill_1 FILLER_115_274 ();
 sg13g2_decap_4 FILLER_115_286 ();
 sg13g2_fill_2 FILLER_115_290 ();
 sg13g2_decap_8 FILLER_115_300 ();
 sg13g2_decap_8 FILLER_115_307 ();
 sg13g2_decap_4 FILLER_115_322 ();
 sg13g2_fill_1 FILLER_115_326 ();
 sg13g2_decap_8 FILLER_115_340 ();
 sg13g2_decap_8 FILLER_115_347 ();
 sg13g2_decap_8 FILLER_115_354 ();
 sg13g2_fill_2 FILLER_115_361 ();
 sg13g2_fill_1 FILLER_115_363 ();
 sg13g2_fill_2 FILLER_115_390 ();
 sg13g2_fill_1 FILLER_115_392 ();
 sg13g2_decap_4 FILLER_115_406 ();
 sg13g2_decap_8 FILLER_115_426 ();
 sg13g2_decap_8 FILLER_115_433 ();
 sg13g2_decap_8 FILLER_115_440 ();
 sg13g2_decap_8 FILLER_115_447 ();
 sg13g2_decap_8 FILLER_115_454 ();
 sg13g2_fill_2 FILLER_115_461 ();
 sg13g2_fill_1 FILLER_115_463 ();
 sg13g2_fill_1 FILLER_115_474 ();
 sg13g2_decap_4 FILLER_115_509 ();
 sg13g2_decap_8 FILLER_115_518 ();
 sg13g2_decap_4 FILLER_115_525 ();
 sg13g2_decap_8 FILLER_115_558 ();
 sg13g2_decap_8 FILLER_115_565 ();
 sg13g2_decap_8 FILLER_115_572 ();
 sg13g2_decap_8 FILLER_115_579 ();
 sg13g2_decap_8 FILLER_115_586 ();
 sg13g2_decap_8 FILLER_115_606 ();
 sg13g2_decap_8 FILLER_115_613 ();
 sg13g2_decap_8 FILLER_115_620 ();
 sg13g2_decap_8 FILLER_115_627 ();
 sg13g2_decap_8 FILLER_115_634 ();
 sg13g2_decap_8 FILLER_115_641 ();
 sg13g2_decap_8 FILLER_115_648 ();
 sg13g2_fill_1 FILLER_115_655 ();
 sg13g2_decap_8 FILLER_115_664 ();
 sg13g2_decap_4 FILLER_115_671 ();
 sg13g2_decap_8 FILLER_115_680 ();
 sg13g2_decap_8 FILLER_115_687 ();
 sg13g2_decap_8 FILLER_115_694 ();
 sg13g2_decap_8 FILLER_115_701 ();
 sg13g2_decap_8 FILLER_115_708 ();
 sg13g2_decap_8 FILLER_115_715 ();
 sg13g2_decap_8 FILLER_115_722 ();
 sg13g2_decap_8 FILLER_115_729 ();
 sg13g2_decap_8 FILLER_115_736 ();
 sg13g2_decap_8 FILLER_115_743 ();
 sg13g2_decap_8 FILLER_115_750 ();
 sg13g2_decap_8 FILLER_115_757 ();
 sg13g2_decap_8 FILLER_115_764 ();
 sg13g2_decap_8 FILLER_115_771 ();
 sg13g2_decap_8 FILLER_115_778 ();
 sg13g2_decap_8 FILLER_115_785 ();
 sg13g2_decap_8 FILLER_115_792 ();
 sg13g2_decap_4 FILLER_115_799 ();
 sg13g2_decap_8 FILLER_115_807 ();
 sg13g2_decap_8 FILLER_115_814 ();
 sg13g2_fill_1 FILLER_115_821 ();
 sg13g2_decap_8 FILLER_115_835 ();
 sg13g2_decap_4 FILLER_115_842 ();
 sg13g2_fill_2 FILLER_115_846 ();
 sg13g2_decap_8 FILLER_115_859 ();
 sg13g2_decap_4 FILLER_115_866 ();
 sg13g2_decap_8 FILLER_115_879 ();
 sg13g2_decap_8 FILLER_115_886 ();
 sg13g2_fill_1 FILLER_115_893 ();
 sg13g2_fill_2 FILLER_115_902 ();
 sg13g2_fill_2 FILLER_115_930 ();
 sg13g2_fill_1 FILLER_115_932 ();
 sg13g2_decap_8 FILLER_115_940 ();
 sg13g2_fill_2 FILLER_115_947 ();
 sg13g2_fill_1 FILLER_115_949 ();
 sg13g2_decap_8 FILLER_115_960 ();
 sg13g2_decap_8 FILLER_115_967 ();
 sg13g2_fill_2 FILLER_115_974 ();
 sg13g2_fill_1 FILLER_115_976 ();
 sg13g2_decap_8 FILLER_115_992 ();
 sg13g2_decap_8 FILLER_115_999 ();
 sg13g2_decap_8 FILLER_115_1006 ();
 sg13g2_decap_8 FILLER_115_1013 ();
 sg13g2_decap_8 FILLER_115_1020 ();
 sg13g2_decap_8 FILLER_115_1027 ();
 sg13g2_decap_8 FILLER_115_1034 ();
 sg13g2_decap_8 FILLER_115_1041 ();
 sg13g2_decap_8 FILLER_115_1048 ();
 sg13g2_decap_8 FILLER_115_1055 ();
 sg13g2_decap_8 FILLER_115_1062 ();
 sg13g2_decap_8 FILLER_115_1069 ();
 sg13g2_fill_1 FILLER_115_1076 ();
 sg13g2_fill_2 FILLER_115_1090 ();
 sg13g2_decap_8 FILLER_115_1111 ();
 sg13g2_decap_8 FILLER_115_1118 ();
 sg13g2_decap_8 FILLER_115_1125 ();
 sg13g2_decap_8 FILLER_115_1132 ();
 sg13g2_fill_1 FILLER_115_1139 ();
 sg13g2_decap_8 FILLER_115_1152 ();
 sg13g2_decap_8 FILLER_115_1159 ();
 sg13g2_fill_2 FILLER_115_1166 ();
 sg13g2_decap_8 FILLER_115_1174 ();
 sg13g2_decap_8 FILLER_115_1181 ();
 sg13g2_decap_8 FILLER_115_1188 ();
 sg13g2_decap_8 FILLER_115_1195 ();
 sg13g2_decap_8 FILLER_115_1202 ();
 sg13g2_decap_8 FILLER_115_1209 ();
 sg13g2_fill_2 FILLER_115_1216 ();
 sg13g2_fill_1 FILLER_115_1218 ();
 sg13g2_decap_8 FILLER_115_1229 ();
 sg13g2_fill_1 FILLER_115_1236 ();
 sg13g2_decap_8 FILLER_115_1241 ();
 sg13g2_decap_8 FILLER_115_1248 ();
 sg13g2_decap_4 FILLER_115_1255 ();
 sg13g2_fill_1 FILLER_115_1259 ();
 sg13g2_decap_8 FILLER_115_1265 ();
 sg13g2_decap_8 FILLER_115_1272 ();
 sg13g2_decap_8 FILLER_115_1279 ();
 sg13g2_decap_8 FILLER_115_1286 ();
 sg13g2_decap_8 FILLER_115_1293 ();
 sg13g2_decap_8 FILLER_115_1300 ();
 sg13g2_decap_8 FILLER_115_1307 ();
 sg13g2_decap_8 FILLER_115_1314 ();
 sg13g2_fill_2 FILLER_115_1321 ();
 sg13g2_fill_2 FILLER_115_1331 ();
 sg13g2_fill_1 FILLER_115_1333 ();
 sg13g2_decap_8 FILLER_115_1337 ();
 sg13g2_decap_8 FILLER_115_1344 ();
 sg13g2_fill_1 FILLER_115_1351 ();
 sg13g2_decap_8 FILLER_115_1370 ();
 sg13g2_decap_8 FILLER_115_1377 ();
 sg13g2_decap_8 FILLER_115_1384 ();
 sg13g2_decap_8 FILLER_115_1391 ();
 sg13g2_decap_8 FILLER_115_1398 ();
 sg13g2_decap_8 FILLER_115_1405 ();
 sg13g2_decap_4 FILLER_115_1412 ();
 sg13g2_decap_8 FILLER_115_1424 ();
 sg13g2_decap_8 FILLER_115_1431 ();
 sg13g2_decap_8 FILLER_115_1438 ();
 sg13g2_decap_8 FILLER_115_1445 ();
 sg13g2_decap_8 FILLER_115_1452 ();
 sg13g2_decap_8 FILLER_115_1459 ();
 sg13g2_decap_8 FILLER_115_1466 ();
 sg13g2_decap_8 FILLER_115_1478 ();
 sg13g2_decap_8 FILLER_115_1485 ();
 sg13g2_decap_4 FILLER_115_1492 ();
 sg13g2_fill_2 FILLER_115_1496 ();
 sg13g2_decap_8 FILLER_115_1506 ();
 sg13g2_fill_2 FILLER_115_1513 ();
 sg13g2_fill_1 FILLER_115_1515 ();
 sg13g2_decap_8 FILLER_115_1537 ();
 sg13g2_decap_8 FILLER_115_1544 ();
 sg13g2_decap_4 FILLER_115_1551 ();
 sg13g2_decap_8 FILLER_115_1563 ();
 sg13g2_decap_8 FILLER_115_1570 ();
 sg13g2_fill_1 FILLER_115_1577 ();
 sg13g2_decap_8 FILLER_115_1591 ();
 sg13g2_fill_1 FILLER_115_1598 ();
 sg13g2_decap_8 FILLER_115_1604 ();
 sg13g2_decap_8 FILLER_115_1611 ();
 sg13g2_decap_8 FILLER_115_1618 ();
 sg13g2_decap_8 FILLER_115_1625 ();
 sg13g2_decap_8 FILLER_115_1632 ();
 sg13g2_decap_4 FILLER_115_1639 ();
 sg13g2_decap_8 FILLER_115_1670 ();
 sg13g2_decap_8 FILLER_115_1690 ();
 sg13g2_decap_8 FILLER_115_1697 ();
 sg13g2_decap_8 FILLER_115_1704 ();
 sg13g2_decap_8 FILLER_115_1711 ();
 sg13g2_decap_8 FILLER_115_1718 ();
 sg13g2_decap_8 FILLER_115_1725 ();
 sg13g2_decap_8 FILLER_115_1732 ();
 sg13g2_decap_8 FILLER_115_1739 ();
 sg13g2_decap_8 FILLER_115_1746 ();
 sg13g2_decap_8 FILLER_115_1753 ();
 sg13g2_decap_8 FILLER_115_1760 ();
 sg13g2_fill_1 FILLER_115_1767 ();
 sg13g2_decap_8 FILLER_116_0 ();
 sg13g2_decap_8 FILLER_116_7 ();
 sg13g2_decap_4 FILLER_116_14 ();
 sg13g2_fill_2 FILLER_116_21 ();
 sg13g2_fill_1 FILLER_116_23 ();
 sg13g2_decap_8 FILLER_116_28 ();
 sg13g2_decap_8 FILLER_116_35 ();
 sg13g2_decap_8 FILLER_116_42 ();
 sg13g2_decap_8 FILLER_116_49 ();
 sg13g2_decap_8 FILLER_116_56 ();
 sg13g2_decap_8 FILLER_116_63 ();
 sg13g2_decap_8 FILLER_116_70 ();
 sg13g2_decap_4 FILLER_116_77 ();
 sg13g2_decap_8 FILLER_116_89 ();
 sg13g2_fill_1 FILLER_116_96 ();
 sg13g2_decap_8 FILLER_116_103 ();
 sg13g2_decap_4 FILLER_116_110 ();
 sg13g2_fill_1 FILLER_116_114 ();
 sg13g2_decap_8 FILLER_116_123 ();
 sg13g2_fill_2 FILLER_116_130 ();
 sg13g2_decap_8 FILLER_116_142 ();
 sg13g2_decap_8 FILLER_116_149 ();
 sg13g2_decap_4 FILLER_116_156 ();
 sg13g2_fill_2 FILLER_116_160 ();
 sg13g2_decap_4 FILLER_116_167 ();
 sg13g2_fill_2 FILLER_116_171 ();
 sg13g2_decap_8 FILLER_116_179 ();
 sg13g2_decap_8 FILLER_116_186 ();
 sg13g2_decap_8 FILLER_116_193 ();
 sg13g2_decap_4 FILLER_116_200 ();
 sg13g2_fill_1 FILLER_116_204 ();
 sg13g2_decap_8 FILLER_116_213 ();
 sg13g2_decap_8 FILLER_116_220 ();
 sg13g2_decap_8 FILLER_116_227 ();
 sg13g2_decap_8 FILLER_116_234 ();
 sg13g2_decap_4 FILLER_116_241 ();
 sg13g2_fill_2 FILLER_116_250 ();
 sg13g2_decap_8 FILLER_116_279 ();
 sg13g2_decap_8 FILLER_116_286 ();
 sg13g2_decap_8 FILLER_116_293 ();
 sg13g2_decap_8 FILLER_116_300 ();
 sg13g2_decap_8 FILLER_116_307 ();
 sg13g2_decap_4 FILLER_116_314 ();
 sg13g2_fill_1 FILLER_116_318 ();
 sg13g2_fill_2 FILLER_116_327 ();
 sg13g2_fill_1 FILLER_116_329 ();
 sg13g2_decap_8 FILLER_116_334 ();
 sg13g2_decap_8 FILLER_116_341 ();
 sg13g2_decap_8 FILLER_116_348 ();
 sg13g2_decap_8 FILLER_116_355 ();
 sg13g2_decap_8 FILLER_116_362 ();
 sg13g2_decap_4 FILLER_116_369 ();
 sg13g2_fill_2 FILLER_116_373 ();
 sg13g2_decap_8 FILLER_116_405 ();
 sg13g2_fill_2 FILLER_116_412 ();
 sg13g2_fill_2 FILLER_116_426 ();
 sg13g2_decap_8 FILLER_116_441 ();
 sg13g2_decap_8 FILLER_116_461 ();
 sg13g2_decap_4 FILLER_116_468 ();
 sg13g2_fill_1 FILLER_116_472 ();
 sg13g2_decap_4 FILLER_116_479 ();
 sg13g2_fill_2 FILLER_116_483 ();
 sg13g2_decap_8 FILLER_116_498 ();
 sg13g2_decap_8 FILLER_116_505 ();
 sg13g2_fill_2 FILLER_116_512 ();
 sg13g2_decap_8 FILLER_116_527 ();
 sg13g2_fill_2 FILLER_116_534 ();
 sg13g2_fill_1 FILLER_116_536 ();
 sg13g2_decap_8 FILLER_116_547 ();
 sg13g2_decap_8 FILLER_116_554 ();
 sg13g2_decap_8 FILLER_116_561 ();
 sg13g2_decap_8 FILLER_116_568 ();
 sg13g2_fill_2 FILLER_116_575 ();
 sg13g2_fill_1 FILLER_116_577 ();
 sg13g2_decap_8 FILLER_116_604 ();
 sg13g2_decap_8 FILLER_116_611 ();
 sg13g2_decap_8 FILLER_116_618 ();
 sg13g2_fill_2 FILLER_116_625 ();
 sg13g2_decap_8 FILLER_116_638 ();
 sg13g2_decap_8 FILLER_116_645 ();
 sg13g2_decap_8 FILLER_116_652 ();
 sg13g2_fill_2 FILLER_116_659 ();
 sg13g2_fill_1 FILLER_116_669 ();
 sg13g2_decap_8 FILLER_116_691 ();
 sg13g2_decap_8 FILLER_116_698 ();
 sg13g2_decap_8 FILLER_116_705 ();
 sg13g2_decap_8 FILLER_116_712 ();
 sg13g2_decap_8 FILLER_116_719 ();
 sg13g2_decap_8 FILLER_116_726 ();
 sg13g2_decap_4 FILLER_116_733 ();
 sg13g2_fill_2 FILLER_116_737 ();
 sg13g2_decap_8 FILLER_116_749 ();
 sg13g2_fill_2 FILLER_116_756 ();
 sg13g2_decap_8 FILLER_116_763 ();
 sg13g2_decap_4 FILLER_116_770 ();
 sg13g2_fill_2 FILLER_116_774 ();
 sg13g2_decap_8 FILLER_116_798 ();
 sg13g2_decap_4 FILLER_116_805 ();
 sg13g2_fill_1 FILLER_116_809 ();
 sg13g2_decap_8 FILLER_116_813 ();
 sg13g2_decap_4 FILLER_116_820 ();
 sg13g2_decap_8 FILLER_116_829 ();
 sg13g2_decap_8 FILLER_116_845 ();
 sg13g2_decap_8 FILLER_116_852 ();
 sg13g2_decap_4 FILLER_116_859 ();
 sg13g2_fill_1 FILLER_116_863 ();
 sg13g2_decap_8 FILLER_116_878 ();
 sg13g2_decap_8 FILLER_116_885 ();
 sg13g2_decap_8 FILLER_116_892 ();
 sg13g2_decap_8 FILLER_116_899 ();
 sg13g2_decap_8 FILLER_116_906 ();
 sg13g2_fill_2 FILLER_116_913 ();
 sg13g2_decap_8 FILLER_116_923 ();
 sg13g2_fill_2 FILLER_116_930 ();
 sg13g2_fill_1 FILLER_116_932 ();
 sg13g2_decap_8 FILLER_116_941 ();
 sg13g2_fill_2 FILLER_116_948 ();
 sg13g2_fill_2 FILLER_116_976 ();
 sg13g2_decap_8 FILLER_116_991 ();
 sg13g2_fill_1 FILLER_116_998 ();
 sg13g2_decap_4 FILLER_116_1012 ();
 sg13g2_fill_2 FILLER_116_1016 ();
 sg13g2_fill_1 FILLER_116_1026 ();
 sg13g2_decap_8 FILLER_116_1036 ();
 sg13g2_decap_8 FILLER_116_1043 ();
 sg13g2_decap_8 FILLER_116_1050 ();
 sg13g2_fill_1 FILLER_116_1057 ();
 sg13g2_decap_8 FILLER_116_1071 ();
 sg13g2_decap_8 FILLER_116_1078 ();
 sg13g2_decap_8 FILLER_116_1085 ();
 sg13g2_decap_4 FILLER_116_1092 ();
 sg13g2_fill_1 FILLER_116_1096 ();
 sg13g2_decap_8 FILLER_116_1101 ();
 sg13g2_decap_8 FILLER_116_1108 ();
 sg13g2_decap_8 FILLER_116_1115 ();
 sg13g2_decap_8 FILLER_116_1122 ();
 sg13g2_decap_8 FILLER_116_1129 ();
 sg13g2_fill_2 FILLER_116_1136 ();
 sg13g2_decap_8 FILLER_116_1146 ();
 sg13g2_decap_8 FILLER_116_1153 ();
 sg13g2_decap_8 FILLER_116_1160 ();
 sg13g2_decap_8 FILLER_116_1167 ();
 sg13g2_decap_8 FILLER_116_1174 ();
 sg13g2_decap_8 FILLER_116_1181 ();
 sg13g2_decap_8 FILLER_116_1188 ();
 sg13g2_fill_2 FILLER_116_1195 ();
 sg13g2_decap_8 FILLER_116_1205 ();
 sg13g2_decap_4 FILLER_116_1212 ();
 sg13g2_fill_2 FILLER_116_1216 ();
 sg13g2_decap_8 FILLER_116_1231 ();
 sg13g2_decap_8 FILLER_116_1238 ();
 sg13g2_decap_8 FILLER_116_1245 ();
 sg13g2_decap_8 FILLER_116_1252 ();
 sg13g2_decap_8 FILLER_116_1259 ();
 sg13g2_decap_8 FILLER_116_1266 ();
 sg13g2_decap_8 FILLER_116_1273 ();
 sg13g2_decap_8 FILLER_116_1280 ();
 sg13g2_decap_8 FILLER_116_1287 ();
 sg13g2_decap_4 FILLER_116_1294 ();
 sg13g2_fill_2 FILLER_116_1298 ();
 sg13g2_decap_8 FILLER_116_1306 ();
 sg13g2_decap_8 FILLER_116_1313 ();
 sg13g2_fill_2 FILLER_116_1320 ();
 sg13g2_fill_1 FILLER_116_1322 ();
 sg13g2_decap_4 FILLER_116_1326 ();
 sg13g2_fill_1 FILLER_116_1330 ();
 sg13g2_decap_4 FILLER_116_1339 ();
 sg13g2_fill_1 FILLER_116_1353 ();
 sg13g2_decap_8 FILLER_116_1358 ();
 sg13g2_decap_8 FILLER_116_1365 ();
 sg13g2_decap_8 FILLER_116_1372 ();
 sg13g2_decap_8 FILLER_116_1387 ();
 sg13g2_decap_8 FILLER_116_1394 ();
 sg13g2_decap_8 FILLER_116_1401 ();
 sg13g2_decap_8 FILLER_116_1408 ();
 sg13g2_decap_8 FILLER_116_1415 ();
 sg13g2_decap_8 FILLER_116_1422 ();
 sg13g2_decap_8 FILLER_116_1429 ();
 sg13g2_decap_8 FILLER_116_1436 ();
 sg13g2_decap_8 FILLER_116_1443 ();
 sg13g2_decap_8 FILLER_116_1450 ();
 sg13g2_decap_8 FILLER_116_1457 ();
 sg13g2_fill_2 FILLER_116_1464 ();
 sg13g2_decap_4 FILLER_116_1474 ();
 sg13g2_fill_2 FILLER_116_1478 ();
 sg13g2_decap_8 FILLER_116_1499 ();
 sg13g2_decap_8 FILLER_116_1506 ();
 sg13g2_fill_2 FILLER_116_1513 ();
 sg13g2_decap_8 FILLER_116_1523 ();
 sg13g2_decap_8 FILLER_116_1530 ();
 sg13g2_decap_8 FILLER_116_1537 ();
 sg13g2_decap_8 FILLER_116_1544 ();
 sg13g2_decap_8 FILLER_116_1551 ();
 sg13g2_decap_8 FILLER_116_1558 ();
 sg13g2_decap_8 FILLER_116_1565 ();
 sg13g2_decap_8 FILLER_116_1572 ();
 sg13g2_decap_8 FILLER_116_1579 ();
 sg13g2_decap_8 FILLER_116_1586 ();
 sg13g2_decap_8 FILLER_116_1593 ();
 sg13g2_decap_8 FILLER_116_1600 ();
 sg13g2_fill_2 FILLER_116_1607 ();
 sg13g2_decap_8 FILLER_116_1621 ();
 sg13g2_decap_8 FILLER_116_1628 ();
 sg13g2_decap_8 FILLER_116_1635 ();
 sg13g2_decap_8 FILLER_116_1642 ();
 sg13g2_decap_8 FILLER_116_1649 ();
 sg13g2_decap_8 FILLER_116_1656 ();
 sg13g2_decap_8 FILLER_116_1663 ();
 sg13g2_decap_8 FILLER_116_1670 ();
 sg13g2_decap_8 FILLER_116_1677 ();
 sg13g2_decap_8 FILLER_116_1684 ();
 sg13g2_decap_8 FILLER_116_1691 ();
 sg13g2_decap_8 FILLER_116_1698 ();
 sg13g2_decap_8 FILLER_116_1705 ();
 sg13g2_decap_8 FILLER_116_1712 ();
 sg13g2_decap_4 FILLER_116_1719 ();
 sg13g2_fill_2 FILLER_116_1723 ();
 sg13g2_fill_2 FILLER_116_1743 ();
 sg13g2_fill_1 FILLER_116_1745 ();
 sg13g2_decap_8 FILLER_116_1752 ();
 sg13g2_decap_8 FILLER_116_1759 ();
 sg13g2_fill_2 FILLER_116_1766 ();
 sg13g2_decap_8 FILLER_117_0 ();
 sg13g2_decap_4 FILLER_117_7 ();
 sg13g2_fill_2 FILLER_117_11 ();
 sg13g2_fill_2 FILLER_117_25 ();
 sg13g2_decap_4 FILLER_117_35 ();
 sg13g2_decap_8 FILLER_117_44 ();
 sg13g2_decap_8 FILLER_117_51 ();
 sg13g2_decap_8 FILLER_117_58 ();
 sg13g2_decap_8 FILLER_117_65 ();
 sg13g2_decap_8 FILLER_117_72 ();
 sg13g2_decap_4 FILLER_117_79 ();
 sg13g2_decap_8 FILLER_117_96 ();
 sg13g2_decap_8 FILLER_117_103 ();
 sg13g2_decap_8 FILLER_117_110 ();
 sg13g2_decap_8 FILLER_117_117 ();
 sg13g2_decap_8 FILLER_117_124 ();
 sg13g2_decap_8 FILLER_117_131 ();
 sg13g2_decap_8 FILLER_117_138 ();
 sg13g2_decap_8 FILLER_117_145 ();
 sg13g2_decap_8 FILLER_117_152 ();
 sg13g2_decap_8 FILLER_117_159 ();
 sg13g2_decap_8 FILLER_117_166 ();
 sg13g2_decap_8 FILLER_117_173 ();
 sg13g2_decap_8 FILLER_117_180 ();
 sg13g2_decap_8 FILLER_117_187 ();
 sg13g2_decap_8 FILLER_117_194 ();
 sg13g2_decap_8 FILLER_117_205 ();
 sg13g2_decap_8 FILLER_117_212 ();
 sg13g2_decap_8 FILLER_117_219 ();
 sg13g2_decap_8 FILLER_117_226 ();
 sg13g2_decap_8 FILLER_117_233 ();
 sg13g2_fill_2 FILLER_117_240 ();
 sg13g2_fill_2 FILLER_117_249 ();
 sg13g2_fill_1 FILLER_117_251 ();
 sg13g2_decap_4 FILLER_117_257 ();
 sg13g2_fill_1 FILLER_117_261 ();
 sg13g2_decap_8 FILLER_117_267 ();
 sg13g2_fill_1 FILLER_117_274 ();
 sg13g2_decap_8 FILLER_117_278 ();
 sg13g2_decap_8 FILLER_117_285 ();
 sg13g2_decap_8 FILLER_117_292 ();
 sg13g2_decap_8 FILLER_117_299 ();
 sg13g2_decap_8 FILLER_117_306 ();
 sg13g2_decap_8 FILLER_117_313 ();
 sg13g2_fill_2 FILLER_117_320 ();
 sg13g2_fill_1 FILLER_117_322 ();
 sg13g2_decap_8 FILLER_117_329 ();
 sg13g2_decap_8 FILLER_117_336 ();
 sg13g2_decap_8 FILLER_117_343 ();
 sg13g2_decap_8 FILLER_117_350 ();
 sg13g2_fill_2 FILLER_117_357 ();
 sg13g2_fill_1 FILLER_117_359 ();
 sg13g2_decap_8 FILLER_117_364 ();
 sg13g2_decap_4 FILLER_117_371 ();
 sg13g2_fill_1 FILLER_117_375 ();
 sg13g2_decap_8 FILLER_117_381 ();
 sg13g2_fill_2 FILLER_117_388 ();
 sg13g2_decap_8 FILLER_117_394 ();
 sg13g2_decap_8 FILLER_117_401 ();
 sg13g2_decap_8 FILLER_117_408 ();
 sg13g2_fill_2 FILLER_117_415 ();
 sg13g2_decap_8 FILLER_117_432 ();
 sg13g2_decap_8 FILLER_117_439 ();
 sg13g2_decap_8 FILLER_117_446 ();
 sg13g2_decap_8 FILLER_117_453 ();
 sg13g2_decap_8 FILLER_117_460 ();
 sg13g2_decap_8 FILLER_117_467 ();
 sg13g2_fill_2 FILLER_117_474 ();
 sg13g2_decap_8 FILLER_117_495 ();
 sg13g2_decap_8 FILLER_117_502 ();
 sg13g2_decap_8 FILLER_117_509 ();
 sg13g2_decap_8 FILLER_117_516 ();
 sg13g2_decap_8 FILLER_117_523 ();
 sg13g2_decap_8 FILLER_117_530 ();
 sg13g2_decap_8 FILLER_117_537 ();
 sg13g2_decap_8 FILLER_117_544 ();
 sg13g2_decap_8 FILLER_117_551 ();
 sg13g2_fill_2 FILLER_117_558 ();
 sg13g2_decap_8 FILLER_117_573 ();
 sg13g2_decap_8 FILLER_117_580 ();
 sg13g2_decap_8 FILLER_117_587 ();
 sg13g2_decap_8 FILLER_117_594 ();
 sg13g2_decap_8 FILLER_117_601 ();
 sg13g2_decap_8 FILLER_117_608 ();
 sg13g2_decap_4 FILLER_117_615 ();
 sg13g2_decap_8 FILLER_117_632 ();
 sg13g2_decap_8 FILLER_117_639 ();
 sg13g2_decap_8 FILLER_117_646 ();
 sg13g2_fill_2 FILLER_117_653 ();
 sg13g2_fill_1 FILLER_117_677 ();
 sg13g2_decap_8 FILLER_117_686 ();
 sg13g2_decap_8 FILLER_117_693 ();
 sg13g2_decap_8 FILLER_117_700 ();
 sg13g2_decap_8 FILLER_117_707 ();
 sg13g2_decap_4 FILLER_117_714 ();
 sg13g2_fill_1 FILLER_117_718 ();
 sg13g2_decap_8 FILLER_117_731 ();
 sg13g2_decap_8 FILLER_117_738 ();
 sg13g2_decap_8 FILLER_117_745 ();
 sg13g2_fill_2 FILLER_117_752 ();
 sg13g2_decap_8 FILLER_117_759 ();
 sg13g2_fill_1 FILLER_117_766 ();
 sg13g2_decap_8 FILLER_117_775 ();
 sg13g2_decap_8 FILLER_117_782 ();
 sg13g2_decap_8 FILLER_117_789 ();
 sg13g2_decap_8 FILLER_117_796 ();
 sg13g2_decap_8 FILLER_117_803 ();
 sg13g2_decap_4 FILLER_117_826 ();
 sg13g2_fill_2 FILLER_117_834 ();
 sg13g2_decap_4 FILLER_117_859 ();
 sg13g2_fill_1 FILLER_117_863 ();
 sg13g2_decap_8 FILLER_117_877 ();
 sg13g2_decap_8 FILLER_117_884 ();
 sg13g2_decap_8 FILLER_117_891 ();
 sg13g2_decap_8 FILLER_117_898 ();
 sg13g2_decap_8 FILLER_117_905 ();
 sg13g2_decap_4 FILLER_117_912 ();
 sg13g2_fill_1 FILLER_117_916 ();
 sg13g2_decap_8 FILLER_117_930 ();
 sg13g2_decap_8 FILLER_117_937 ();
 sg13g2_decap_8 FILLER_117_944 ();
 sg13g2_decap_4 FILLER_117_951 ();
 sg13g2_fill_1 FILLER_117_955 ();
 sg13g2_decap_8 FILLER_117_969 ();
 sg13g2_decap_8 FILLER_117_976 ();
 sg13g2_decap_8 FILLER_117_983 ();
 sg13g2_decap_8 FILLER_117_990 ();
 sg13g2_decap_8 FILLER_117_997 ();
 sg13g2_decap_8 FILLER_117_1004 ();
 sg13g2_decap_8 FILLER_117_1011 ();
 sg13g2_decap_8 FILLER_117_1018 ();
 sg13g2_decap_8 FILLER_117_1025 ();
 sg13g2_decap_8 FILLER_117_1032 ();
 sg13g2_decap_4 FILLER_117_1039 ();
 sg13g2_decap_8 FILLER_117_1069 ();
 sg13g2_decap_8 FILLER_117_1076 ();
 sg13g2_decap_8 FILLER_117_1083 ();
 sg13g2_decap_8 FILLER_117_1090 ();
 sg13g2_decap_8 FILLER_117_1097 ();
 sg13g2_decap_8 FILLER_117_1104 ();
 sg13g2_decap_8 FILLER_117_1111 ();
 sg13g2_fill_1 FILLER_117_1118 ();
 sg13g2_decap_8 FILLER_117_1123 ();
 sg13g2_decap_8 FILLER_117_1130 ();
 sg13g2_decap_8 FILLER_117_1137 ();
 sg13g2_decap_8 FILLER_117_1144 ();
 sg13g2_decap_8 FILLER_117_1151 ();
 sg13g2_decap_8 FILLER_117_1158 ();
 sg13g2_decap_4 FILLER_117_1165 ();
 sg13g2_decap_8 FILLER_117_1174 ();
 sg13g2_decap_8 FILLER_117_1181 ();
 sg13g2_decap_8 FILLER_117_1188 ();
 sg13g2_decap_8 FILLER_117_1195 ();
 sg13g2_decap_8 FILLER_117_1208 ();
 sg13g2_decap_8 FILLER_117_1215 ();
 sg13g2_decap_4 FILLER_117_1222 ();
 sg13g2_decap_8 FILLER_117_1239 ();
 sg13g2_decap_8 FILLER_117_1246 ();
 sg13g2_decap_4 FILLER_117_1253 ();
 sg13g2_decap_8 FILLER_117_1268 ();
 sg13g2_decap_8 FILLER_117_1275 ();
 sg13g2_decap_8 FILLER_117_1282 ();
 sg13g2_fill_1 FILLER_117_1294 ();
 sg13g2_decap_8 FILLER_117_1311 ();
 sg13g2_fill_2 FILLER_117_1318 ();
 sg13g2_fill_2 FILLER_117_1332 ();
 sg13g2_decap_8 FILLER_117_1365 ();
 sg13g2_decap_8 FILLER_117_1372 ();
 sg13g2_decap_8 FILLER_117_1379 ();
 sg13g2_fill_2 FILLER_117_1386 ();
 sg13g2_fill_1 FILLER_117_1388 ();
 sg13g2_decap_8 FILLER_117_1405 ();
 sg13g2_decap_8 FILLER_117_1412 ();
 sg13g2_decap_8 FILLER_117_1432 ();
 sg13g2_decap_8 FILLER_117_1439 ();
 sg13g2_decap_8 FILLER_117_1446 ();
 sg13g2_fill_1 FILLER_117_1453 ();
 sg13g2_fill_2 FILLER_117_1462 ();
 sg13g2_fill_2 FILLER_117_1484 ();
 sg13g2_fill_2 FILLER_117_1501 ();
 sg13g2_fill_1 FILLER_117_1503 ();
 sg13g2_decap_8 FILLER_117_1512 ();
 sg13g2_decap_8 FILLER_117_1519 ();
 sg13g2_decap_8 FILLER_117_1526 ();
 sg13g2_decap_8 FILLER_117_1533 ();
 sg13g2_decap_8 FILLER_117_1549 ();
 sg13g2_decap_8 FILLER_117_1556 ();
 sg13g2_decap_8 FILLER_117_1563 ();
 sg13g2_decap_8 FILLER_117_1570 ();
 sg13g2_decap_8 FILLER_117_1577 ();
 sg13g2_decap_8 FILLER_117_1584 ();
 sg13g2_decap_4 FILLER_117_1591 ();
 sg13g2_decap_4 FILLER_117_1615 ();
 sg13g2_fill_1 FILLER_117_1619 ();
 sg13g2_decap_8 FILLER_117_1625 ();
 sg13g2_decap_8 FILLER_117_1632 ();
 sg13g2_decap_4 FILLER_117_1639 ();
 sg13g2_decap_8 FILLER_117_1648 ();
 sg13g2_decap_8 FILLER_117_1655 ();
 sg13g2_decap_8 FILLER_117_1662 ();
 sg13g2_decap_8 FILLER_117_1669 ();
 sg13g2_decap_8 FILLER_117_1676 ();
 sg13g2_decap_8 FILLER_117_1683 ();
 sg13g2_decap_8 FILLER_117_1690 ();
 sg13g2_decap_8 FILLER_117_1697 ();
 sg13g2_decap_8 FILLER_117_1704 ();
 sg13g2_decap_8 FILLER_117_1711 ();
 sg13g2_decap_8 FILLER_117_1718 ();
 sg13g2_decap_8 FILLER_117_1750 ();
 sg13g2_decap_8 FILLER_117_1757 ();
 sg13g2_decap_4 FILLER_117_1764 ();
 sg13g2_decap_8 FILLER_118_0 ();
 sg13g2_decap_8 FILLER_118_7 ();
 sg13g2_decap_8 FILLER_118_14 ();
 sg13g2_fill_2 FILLER_118_36 ();
 sg13g2_decap_8 FILLER_118_54 ();
 sg13g2_decap_8 FILLER_118_61 ();
 sg13g2_decap_8 FILLER_118_68 ();
 sg13g2_decap_8 FILLER_118_101 ();
 sg13g2_decap_8 FILLER_118_108 ();
 sg13g2_fill_2 FILLER_118_115 ();
 sg13g2_fill_1 FILLER_118_117 ();
 sg13g2_decap_8 FILLER_118_127 ();
 sg13g2_decap_8 FILLER_118_134 ();
 sg13g2_decap_4 FILLER_118_141 ();
 sg13g2_decap_8 FILLER_118_153 ();
 sg13g2_decap_8 FILLER_118_160 ();
 sg13g2_decap_8 FILLER_118_167 ();
 sg13g2_decap_8 FILLER_118_182 ();
 sg13g2_decap_8 FILLER_118_189 ();
 sg13g2_decap_4 FILLER_118_196 ();
 sg13g2_decap_8 FILLER_118_208 ();
 sg13g2_decap_8 FILLER_118_215 ();
 sg13g2_decap_4 FILLER_118_222 ();
 sg13g2_fill_1 FILLER_118_226 ();
 sg13g2_decap_8 FILLER_118_234 ();
 sg13g2_decap_8 FILLER_118_241 ();
 sg13g2_fill_2 FILLER_118_248 ();
 sg13g2_decap_8 FILLER_118_281 ();
 sg13g2_decap_8 FILLER_118_288 ();
 sg13g2_decap_8 FILLER_118_295 ();
 sg13g2_decap_8 FILLER_118_302 ();
 sg13g2_decap_8 FILLER_118_309 ();
 sg13g2_fill_2 FILLER_118_316 ();
 sg13g2_fill_1 FILLER_118_318 ();
 sg13g2_decap_8 FILLER_118_338 ();
 sg13g2_decap_8 FILLER_118_345 ();
 sg13g2_decap_8 FILLER_118_352 ();
 sg13g2_fill_2 FILLER_118_359 ();
 sg13g2_decap_8 FILLER_118_378 ();
 sg13g2_decap_8 FILLER_118_385 ();
 sg13g2_decap_8 FILLER_118_392 ();
 sg13g2_decap_4 FILLER_118_399 ();
 sg13g2_fill_2 FILLER_118_420 ();
 sg13g2_decap_8 FILLER_118_437 ();
 sg13g2_decap_8 FILLER_118_444 ();
 sg13g2_decap_8 FILLER_118_451 ();
 sg13g2_decap_8 FILLER_118_458 ();
 sg13g2_fill_1 FILLER_118_465 ();
 sg13g2_decap_8 FILLER_118_474 ();
 sg13g2_decap_8 FILLER_118_481 ();
 sg13g2_decap_8 FILLER_118_488 ();
 sg13g2_decap_8 FILLER_118_495 ();
 sg13g2_decap_8 FILLER_118_502 ();
 sg13g2_decap_8 FILLER_118_509 ();
 sg13g2_decap_8 FILLER_118_516 ();
 sg13g2_fill_2 FILLER_118_523 ();
 sg13g2_fill_1 FILLER_118_525 ();
 sg13g2_decap_8 FILLER_118_530 ();
 sg13g2_decap_8 FILLER_118_537 ();
 sg13g2_decap_8 FILLER_118_544 ();
 sg13g2_decap_8 FILLER_118_551 ();
 sg13g2_decap_8 FILLER_118_558 ();
 sg13g2_fill_2 FILLER_118_565 ();
 sg13g2_decap_8 FILLER_118_605 ();
 sg13g2_fill_2 FILLER_118_612 ();
 sg13g2_decap_8 FILLER_118_622 ();
 sg13g2_decap_8 FILLER_118_629 ();
 sg13g2_decap_8 FILLER_118_636 ();
 sg13g2_decap_8 FILLER_118_643 ();
 sg13g2_decap_8 FILLER_118_650 ();
 sg13g2_decap_4 FILLER_118_657 ();
 sg13g2_fill_1 FILLER_118_661 ();
 sg13g2_decap_8 FILLER_118_678 ();
 sg13g2_decap_8 FILLER_118_685 ();
 sg13g2_decap_4 FILLER_118_696 ();
 sg13g2_decap_8 FILLER_118_708 ();
 sg13g2_fill_2 FILLER_118_715 ();
 sg13g2_fill_1 FILLER_118_717 ();
 sg13g2_decap_8 FILLER_118_737 ();
 sg13g2_decap_8 FILLER_118_744 ();
 sg13g2_decap_8 FILLER_118_751 ();
 sg13g2_decap_4 FILLER_118_758 ();
 sg13g2_fill_1 FILLER_118_762 ();
 sg13g2_decap_4 FILLER_118_779 ();
 sg13g2_fill_1 FILLER_118_783 ();
 sg13g2_decap_8 FILLER_118_794 ();
 sg13g2_decap_4 FILLER_118_801 ();
 sg13g2_fill_2 FILLER_118_805 ();
 sg13g2_decap_4 FILLER_118_832 ();
 sg13g2_fill_1 FILLER_118_836 ();
 sg13g2_decap_8 FILLER_118_845 ();
 sg13g2_decap_8 FILLER_118_852 ();
 sg13g2_decap_8 FILLER_118_859 ();
 sg13g2_decap_8 FILLER_118_866 ();
 sg13g2_decap_4 FILLER_118_873 ();
 sg13g2_fill_1 FILLER_118_877 ();
 sg13g2_decap_8 FILLER_118_891 ();
 sg13g2_decap_8 FILLER_118_898 ();
 sg13g2_decap_8 FILLER_118_905 ();
 sg13g2_decap_8 FILLER_118_912 ();
 sg13g2_decap_8 FILLER_118_919 ();
 sg13g2_decap_8 FILLER_118_926 ();
 sg13g2_decap_8 FILLER_118_933 ();
 sg13g2_decap_8 FILLER_118_940 ();
 sg13g2_decap_8 FILLER_118_947 ();
 sg13g2_decap_8 FILLER_118_980 ();
 sg13g2_decap_8 FILLER_118_987 ();
 sg13g2_decap_8 FILLER_118_994 ();
 sg13g2_decap_8 FILLER_118_1001 ();
 sg13g2_decap_8 FILLER_118_1008 ();
 sg13g2_fill_2 FILLER_118_1015 ();
 sg13g2_fill_1 FILLER_118_1017 ();
 sg13g2_decap_8 FILLER_118_1021 ();
 sg13g2_decap_8 FILLER_118_1028 ();
 sg13g2_decap_8 FILLER_118_1035 ();
 sg13g2_decap_8 FILLER_118_1042 ();
 sg13g2_decap_4 FILLER_118_1049 ();
 sg13g2_fill_1 FILLER_118_1053 ();
 sg13g2_decap_8 FILLER_118_1058 ();
 sg13g2_decap_8 FILLER_118_1065 ();
 sg13g2_decap_8 FILLER_118_1072 ();
 sg13g2_fill_1 FILLER_118_1088 ();
 sg13g2_decap_8 FILLER_118_1107 ();
 sg13g2_fill_1 FILLER_118_1114 ();
 sg13g2_decap_8 FILLER_118_1163 ();
 sg13g2_decap_8 FILLER_118_1183 ();
 sg13g2_decap_8 FILLER_118_1190 ();
 sg13g2_decap_8 FILLER_118_1197 ();
 sg13g2_decap_8 FILLER_118_1204 ();
 sg13g2_decap_8 FILLER_118_1211 ();
 sg13g2_decap_8 FILLER_118_1218 ();
 sg13g2_fill_2 FILLER_118_1225 ();
 sg13g2_decap_8 FILLER_118_1243 ();
 sg13g2_decap_4 FILLER_118_1250 ();
 sg13g2_fill_1 FILLER_118_1254 ();
 sg13g2_decap_8 FILLER_118_1279 ();
 sg13g2_decap_4 FILLER_118_1286 ();
 sg13g2_fill_1 FILLER_118_1290 ();
 sg13g2_decap_8 FILLER_118_1304 ();
 sg13g2_decap_8 FILLER_118_1311 ();
 sg13g2_decap_4 FILLER_118_1318 ();
 sg13g2_fill_1 FILLER_118_1322 ();
 sg13g2_fill_1 FILLER_118_1326 ();
 sg13g2_fill_2 FILLER_118_1349 ();
 sg13g2_fill_1 FILLER_118_1351 ();
 sg13g2_decap_8 FILLER_118_1358 ();
 sg13g2_decap_8 FILLER_118_1365 ();
 sg13g2_decap_8 FILLER_118_1372 ();
 sg13g2_decap_8 FILLER_118_1379 ();
 sg13g2_decap_8 FILLER_118_1386 ();
 sg13g2_decap_8 FILLER_118_1393 ();
 sg13g2_decap_8 FILLER_118_1400 ();
 sg13g2_decap_8 FILLER_118_1407 ();
 sg13g2_decap_4 FILLER_118_1414 ();
 sg13g2_decap_8 FILLER_118_1446 ();
 sg13g2_decap_8 FILLER_118_1453 ();
 sg13g2_decap_8 FILLER_118_1460 ();
 sg13g2_decap_8 FILLER_118_1479 ();
 sg13g2_decap_8 FILLER_118_1486 ();
 sg13g2_decap_8 FILLER_118_1493 ();
 sg13g2_decap_8 FILLER_118_1500 ();
 sg13g2_decap_8 FILLER_118_1520 ();
 sg13g2_decap_8 FILLER_118_1527 ();
 sg13g2_decap_8 FILLER_118_1543 ();
 sg13g2_decap_4 FILLER_118_1550 ();
 sg13g2_fill_1 FILLER_118_1554 ();
 sg13g2_decap_8 FILLER_118_1567 ();
 sg13g2_decap_8 FILLER_118_1574 ();
 sg13g2_decap_4 FILLER_118_1581 ();
 sg13g2_fill_1 FILLER_118_1585 ();
 sg13g2_fill_2 FILLER_118_1594 ();
 sg13g2_fill_2 FILLER_118_1604 ();
 sg13g2_decap_4 FILLER_118_1638 ();
 sg13g2_fill_2 FILLER_118_1642 ();
 sg13g2_fill_2 FILLER_118_1649 ();
 sg13g2_decap_8 FILLER_118_1659 ();
 sg13g2_decap_4 FILLER_118_1666 ();
 sg13g2_fill_2 FILLER_118_1670 ();
 sg13g2_decap_4 FILLER_118_1679 ();
 sg13g2_decap_4 FILLER_118_1705 ();
 sg13g2_fill_1 FILLER_118_1709 ();
 sg13g2_decap_8 FILLER_118_1713 ();
 sg13g2_fill_2 FILLER_118_1720 ();
 sg13g2_fill_1 FILLER_118_1722 ();
 sg13g2_fill_1 FILLER_118_1727 ();
 sg13g2_decap_8 FILLER_118_1752 ();
 sg13g2_decap_8 FILLER_118_1759 ();
 sg13g2_fill_2 FILLER_118_1766 ();
 sg13g2_decap_8 FILLER_119_0 ();
 sg13g2_decap_8 FILLER_119_7 ();
 sg13g2_decap_8 FILLER_119_14 ();
 sg13g2_decap_4 FILLER_119_21 ();
 sg13g2_decap_4 FILLER_119_30 ();
 sg13g2_fill_1 FILLER_119_34 ();
 sg13g2_decap_8 FILLER_119_43 ();
 sg13g2_decap_8 FILLER_119_50 ();
 sg13g2_decap_8 FILLER_119_57 ();
 sg13g2_decap_8 FILLER_119_64 ();
 sg13g2_decap_4 FILLER_119_71 ();
 sg13g2_fill_1 FILLER_119_75 ();
 sg13g2_decap_8 FILLER_119_94 ();
 sg13g2_decap_8 FILLER_119_101 ();
 sg13g2_fill_2 FILLER_119_108 ();
 sg13g2_fill_1 FILLER_119_110 ();
 sg13g2_fill_2 FILLER_119_127 ();
 sg13g2_fill_1 FILLER_119_129 ();
 sg13g2_decap_4 FILLER_119_137 ();
 sg13g2_fill_2 FILLER_119_141 ();
 sg13g2_decap_8 FILLER_119_147 ();
 sg13g2_fill_1 FILLER_119_154 ();
 sg13g2_decap_8 FILLER_119_159 ();
 sg13g2_decap_8 FILLER_119_174 ();
 sg13g2_decap_8 FILLER_119_181 ();
 sg13g2_decap_8 FILLER_119_188 ();
 sg13g2_fill_2 FILLER_119_195 ();
 sg13g2_decap_4 FILLER_119_221 ();
 sg13g2_fill_2 FILLER_119_225 ();
 sg13g2_decap_8 FILLER_119_235 ();
 sg13g2_decap_8 FILLER_119_242 ();
 sg13g2_decap_8 FILLER_119_249 ();
 sg13g2_decap_8 FILLER_119_264 ();
 sg13g2_decap_8 FILLER_119_271 ();
 sg13g2_decap_8 FILLER_119_278 ();
 sg13g2_decap_8 FILLER_119_290 ();
 sg13g2_decap_4 FILLER_119_305 ();
 sg13g2_decap_8 FILLER_119_334 ();
 sg13g2_decap_8 FILLER_119_341 ();
 sg13g2_decap_8 FILLER_119_352 ();
 sg13g2_fill_1 FILLER_119_359 ();
 sg13g2_decap_8 FILLER_119_364 ();
 sg13g2_decap_8 FILLER_119_371 ();
 sg13g2_decap_8 FILLER_119_378 ();
 sg13g2_decap_8 FILLER_119_385 ();
 sg13g2_decap_4 FILLER_119_392 ();
 sg13g2_fill_1 FILLER_119_396 ();
 sg13g2_decap_4 FILLER_119_410 ();
 sg13g2_decap_4 FILLER_119_422 ();
 sg13g2_decap_8 FILLER_119_435 ();
 sg13g2_decap_8 FILLER_119_442 ();
 sg13g2_decap_8 FILLER_119_449 ();
 sg13g2_decap_8 FILLER_119_456 ();
 sg13g2_decap_4 FILLER_119_463 ();
 sg13g2_fill_2 FILLER_119_467 ();
 sg13g2_decap_8 FILLER_119_473 ();
 sg13g2_decap_8 FILLER_119_480 ();
 sg13g2_decap_8 FILLER_119_487 ();
 sg13g2_decap_8 FILLER_119_494 ();
 sg13g2_decap_4 FILLER_119_501 ();
 sg13g2_decap_4 FILLER_119_517 ();
 sg13g2_decap_4 FILLER_119_539 ();
 sg13g2_decap_8 FILLER_119_547 ();
 sg13g2_decap_8 FILLER_119_554 ();
 sg13g2_decap_8 FILLER_119_561 ();
 sg13g2_decap_8 FILLER_119_568 ();
 sg13g2_decap_8 FILLER_119_575 ();
 sg13g2_decap_8 FILLER_119_582 ();
 sg13g2_decap_8 FILLER_119_589 ();
 sg13g2_decap_8 FILLER_119_596 ();
 sg13g2_decap_8 FILLER_119_603 ();
 sg13g2_decap_8 FILLER_119_610 ();
 sg13g2_fill_2 FILLER_119_617 ();
 sg13g2_fill_1 FILLER_119_619 ();
 sg13g2_decap_8 FILLER_119_625 ();
 sg13g2_decap_8 FILLER_119_632 ();
 sg13g2_decap_8 FILLER_119_639 ();
 sg13g2_decap_4 FILLER_119_646 ();
 sg13g2_decap_8 FILLER_119_656 ();
 sg13g2_decap_8 FILLER_119_663 ();
 sg13g2_decap_8 FILLER_119_670 ();
 sg13g2_decap_8 FILLER_119_677 ();
 sg13g2_fill_1 FILLER_119_684 ();
 sg13g2_decap_8 FILLER_119_703 ();
 sg13g2_decap_8 FILLER_119_710 ();
 sg13g2_decap_8 FILLER_119_717 ();
 sg13g2_decap_8 FILLER_119_724 ();
 sg13g2_decap_8 FILLER_119_731 ();
 sg13g2_decap_8 FILLER_119_738 ();
 sg13g2_decap_8 FILLER_119_745 ();
 sg13g2_decap_8 FILLER_119_752 ();
 sg13g2_fill_2 FILLER_119_759 ();
 sg13g2_fill_1 FILLER_119_761 ();
 sg13g2_decap_8 FILLER_119_787 ();
 sg13g2_decap_8 FILLER_119_794 ();
 sg13g2_decap_8 FILLER_119_801 ();
 sg13g2_decap_8 FILLER_119_808 ();
 sg13g2_decap_4 FILLER_119_823 ();
 sg13g2_decap_8 FILLER_119_835 ();
 sg13g2_decap_4 FILLER_119_842 ();
 sg13g2_fill_1 FILLER_119_846 ();
 sg13g2_decap_8 FILLER_119_851 ();
 sg13g2_decap_8 FILLER_119_858 ();
 sg13g2_decap_8 FILLER_119_865 ();
 sg13g2_fill_1 FILLER_119_872 ();
 sg13g2_fill_2 FILLER_119_894 ();
 sg13g2_fill_1 FILLER_119_896 ();
 sg13g2_decap_8 FILLER_119_910 ();
 sg13g2_fill_1 FILLER_119_917 ();
 sg13g2_decap_8 FILLER_119_931 ();
 sg13g2_decap_8 FILLER_119_938 ();
 sg13g2_decap_8 FILLER_119_945 ();
 sg13g2_decap_8 FILLER_119_952 ();
 sg13g2_fill_2 FILLER_119_959 ();
 sg13g2_decap_8 FILLER_119_981 ();
 sg13g2_decap_8 FILLER_119_988 ();
 sg13g2_decap_8 FILLER_119_995 ();
 sg13g2_decap_8 FILLER_119_1002 ();
 sg13g2_decap_4 FILLER_119_1009 ();
 sg13g2_fill_2 FILLER_119_1048 ();
 sg13g2_decap_8 FILLER_119_1063 ();
 sg13g2_decap_8 FILLER_119_1070 ();
 sg13g2_decap_8 FILLER_119_1077 ();
 sg13g2_decap_8 FILLER_119_1084 ();
 sg13g2_decap_8 FILLER_119_1091 ();
 sg13g2_decap_8 FILLER_119_1098 ();
 sg13g2_decap_8 FILLER_119_1105 ();
 sg13g2_fill_2 FILLER_119_1112 ();
 sg13g2_decap_8 FILLER_119_1119 ();
 sg13g2_decap_8 FILLER_119_1126 ();
 sg13g2_fill_2 FILLER_119_1133 ();
 sg13g2_decap_8 FILLER_119_1139 ();
 sg13g2_decap_8 FILLER_119_1146 ();
 sg13g2_decap_8 FILLER_119_1153 ();
 sg13g2_decap_8 FILLER_119_1160 ();
 sg13g2_fill_1 FILLER_119_1167 ();
 sg13g2_fill_1 FILLER_119_1175 ();
 sg13g2_decap_8 FILLER_119_1195 ();
 sg13g2_decap_8 FILLER_119_1202 ();
 sg13g2_decap_8 FILLER_119_1209 ();
 sg13g2_decap_8 FILLER_119_1216 ();
 sg13g2_decap_8 FILLER_119_1223 ();
 sg13g2_fill_2 FILLER_119_1230 ();
 sg13g2_decap_8 FILLER_119_1240 ();
 sg13g2_decap_8 FILLER_119_1247 ();
 sg13g2_decap_4 FILLER_119_1254 ();
 sg13g2_fill_2 FILLER_119_1258 ();
 sg13g2_fill_1 FILLER_119_1265 ();
 sg13g2_decap_8 FILLER_119_1274 ();
 sg13g2_decap_8 FILLER_119_1281 ();
 sg13g2_decap_8 FILLER_119_1288 ();
 sg13g2_decap_4 FILLER_119_1295 ();
 sg13g2_fill_1 FILLER_119_1299 ();
 sg13g2_decap_8 FILLER_119_1313 ();
 sg13g2_decap_8 FILLER_119_1320 ();
 sg13g2_decap_8 FILLER_119_1327 ();
 sg13g2_decap_8 FILLER_119_1334 ();
 sg13g2_decap_8 FILLER_119_1341 ();
 sg13g2_decap_4 FILLER_119_1348 ();
 sg13g2_decap_8 FILLER_119_1381 ();
 sg13g2_fill_2 FILLER_119_1388 ();
 sg13g2_decap_8 FILLER_119_1398 ();
 sg13g2_decap_8 FILLER_119_1405 ();
 sg13g2_decap_8 FILLER_119_1412 ();
 sg13g2_decap_8 FILLER_119_1419 ();
 sg13g2_decap_4 FILLER_119_1426 ();
 sg13g2_decap_8 FILLER_119_1452 ();
 sg13g2_decap_8 FILLER_119_1459 ();
 sg13g2_decap_8 FILLER_119_1466 ();
 sg13g2_decap_8 FILLER_119_1473 ();
 sg13g2_decap_8 FILLER_119_1480 ();
 sg13g2_decap_8 FILLER_119_1487 ();
 sg13g2_decap_4 FILLER_119_1494 ();
 sg13g2_fill_2 FILLER_119_1502 ();
 sg13g2_fill_1 FILLER_119_1504 ();
 sg13g2_decap_4 FILLER_119_1517 ();
 sg13g2_decap_8 FILLER_119_1526 ();
 sg13g2_decap_8 FILLER_119_1533 ();
 sg13g2_decap_8 FILLER_119_1540 ();
 sg13g2_fill_2 FILLER_119_1547 ();
 sg13g2_fill_1 FILLER_119_1549 ();
 sg13g2_decap_8 FILLER_119_1561 ();
 sg13g2_decap_8 FILLER_119_1568 ();
 sg13g2_decap_8 FILLER_119_1575 ();
 sg13g2_fill_2 FILLER_119_1592 ();
 sg13g2_decap_8 FILLER_119_1602 ();
 sg13g2_decap_8 FILLER_119_1609 ();
 sg13g2_decap_4 FILLER_119_1616 ();
 sg13g2_decap_8 FILLER_119_1629 ();
 sg13g2_decap_8 FILLER_119_1636 ();
 sg13g2_decap_8 FILLER_119_1643 ();
 sg13g2_decap_8 FILLER_119_1650 ();
 sg13g2_decap_4 FILLER_119_1657 ();
 sg13g2_fill_2 FILLER_119_1661 ();
 sg13g2_fill_1 FILLER_119_1676 ();
 sg13g2_decap_4 FILLER_119_1702 ();
 sg13g2_fill_1 FILLER_119_1726 ();
 sg13g2_fill_1 FILLER_119_1740 ();
 sg13g2_decap_8 FILLER_119_1749 ();
 sg13g2_decap_8 FILLER_119_1756 ();
 sg13g2_decap_4 FILLER_119_1763 ();
 sg13g2_fill_1 FILLER_119_1767 ();
 sg13g2_decap_8 FILLER_120_0 ();
 sg13g2_decap_8 FILLER_120_7 ();
 sg13g2_fill_1 FILLER_120_14 ();
 sg13g2_decap_4 FILLER_120_19 ();
 sg13g2_fill_2 FILLER_120_23 ();
 sg13g2_decap_8 FILLER_120_51 ();
 sg13g2_decap_8 FILLER_120_58 ();
 sg13g2_decap_8 FILLER_120_65 ();
 sg13g2_decap_8 FILLER_120_72 ();
 sg13g2_decap_8 FILLER_120_79 ();
 sg13g2_decap_8 FILLER_120_86 ();
 sg13g2_decap_8 FILLER_120_93 ();
 sg13g2_decap_8 FILLER_120_100 ();
 sg13g2_decap_8 FILLER_120_107 ();
 sg13g2_decap_8 FILLER_120_114 ();
 sg13g2_fill_1 FILLER_120_121 ();
 sg13g2_decap_8 FILLER_120_126 ();
 sg13g2_decap_4 FILLER_120_133 ();
 sg13g2_fill_1 FILLER_120_137 ();
 sg13g2_decap_8 FILLER_120_146 ();
 sg13g2_fill_2 FILLER_120_153 ();
 sg13g2_decap_8 FILLER_120_179 ();
 sg13g2_decap_8 FILLER_120_186 ();
 sg13g2_decap_8 FILLER_120_199 ();
 sg13g2_decap_8 FILLER_120_206 ();
 sg13g2_decap_8 FILLER_120_213 ();
 sg13g2_decap_8 FILLER_120_220 ();
 sg13g2_decap_8 FILLER_120_227 ();
 sg13g2_decap_8 FILLER_120_234 ();
 sg13g2_decap_8 FILLER_120_241 ();
 sg13g2_decap_8 FILLER_120_248 ();
 sg13g2_decap_8 FILLER_120_255 ();
 sg13g2_decap_8 FILLER_120_262 ();
 sg13g2_decap_8 FILLER_120_269 ();
 sg13g2_decap_8 FILLER_120_276 ();
 sg13g2_fill_1 FILLER_120_283 ();
 sg13g2_fill_2 FILLER_120_301 ();
 sg13g2_fill_1 FILLER_120_303 ();
 sg13g2_fill_1 FILLER_120_317 ();
 sg13g2_decap_8 FILLER_120_328 ();
 sg13g2_decap_8 FILLER_120_335 ();
 sg13g2_decap_4 FILLER_120_342 ();
 sg13g2_decap_8 FILLER_120_354 ();
 sg13g2_decap_8 FILLER_120_361 ();
 sg13g2_decap_8 FILLER_120_368 ();
 sg13g2_decap_8 FILLER_120_375 ();
 sg13g2_decap_8 FILLER_120_382 ();
 sg13g2_decap_8 FILLER_120_389 ();
 sg13g2_decap_4 FILLER_120_396 ();
 sg13g2_decap_8 FILLER_120_404 ();
 sg13g2_decap_8 FILLER_120_411 ();
 sg13g2_decap_4 FILLER_120_418 ();
 sg13g2_decap_8 FILLER_120_430 ();
 sg13g2_decap_4 FILLER_120_437 ();
 sg13g2_decap_8 FILLER_120_466 ();
 sg13g2_decap_8 FILLER_120_473 ();
 sg13g2_decap_8 FILLER_120_480 ();
 sg13g2_decap_8 FILLER_120_487 ();
 sg13g2_decap_8 FILLER_120_494 ();
 sg13g2_decap_8 FILLER_120_501 ();
 sg13g2_fill_2 FILLER_120_508 ();
 sg13g2_decap_8 FILLER_120_548 ();
 sg13g2_fill_2 FILLER_120_555 ();
 sg13g2_decap_8 FILLER_120_561 ();
 sg13g2_decap_8 FILLER_120_568 ();
 sg13g2_decap_8 FILLER_120_575 ();
 sg13g2_decap_8 FILLER_120_582 ();
 sg13g2_fill_1 FILLER_120_589 ();
 sg13g2_decap_8 FILLER_120_603 ();
 sg13g2_decap_8 FILLER_120_610 ();
 sg13g2_decap_8 FILLER_120_617 ();
 sg13g2_fill_1 FILLER_120_624 ();
 sg13g2_decap_4 FILLER_120_630 ();
 sg13g2_fill_2 FILLER_120_634 ();
 sg13g2_decap_8 FILLER_120_655 ();
 sg13g2_decap_8 FILLER_120_662 ();
 sg13g2_decap_8 FILLER_120_669 ();
 sg13g2_decap_8 FILLER_120_676 ();
 sg13g2_fill_2 FILLER_120_683 ();
 sg13g2_fill_1 FILLER_120_685 ();
 sg13g2_fill_1 FILLER_120_691 ();
 sg13g2_decap_8 FILLER_120_699 ();
 sg13g2_decap_8 FILLER_120_706 ();
 sg13g2_decap_8 FILLER_120_713 ();
 sg13g2_decap_8 FILLER_120_720 ();
 sg13g2_fill_2 FILLER_120_727 ();
 sg13g2_fill_1 FILLER_120_729 ();
 sg13g2_decap_4 FILLER_120_738 ();
 sg13g2_decap_8 FILLER_120_746 ();
 sg13g2_decap_8 FILLER_120_753 ();
 sg13g2_decap_8 FILLER_120_760 ();
 sg13g2_fill_2 FILLER_120_767 ();
 sg13g2_decap_8 FILLER_120_779 ();
 sg13g2_decap_8 FILLER_120_786 ();
 sg13g2_decap_8 FILLER_120_793 ();
 sg13g2_decap_8 FILLER_120_800 ();
 sg13g2_decap_8 FILLER_120_807 ();
 sg13g2_decap_8 FILLER_120_814 ();
 sg13g2_decap_8 FILLER_120_821 ();
 sg13g2_decap_8 FILLER_120_828 ();
 sg13g2_decap_8 FILLER_120_835 ();
 sg13g2_decap_8 FILLER_120_842 ();
 sg13g2_decap_4 FILLER_120_849 ();
 sg13g2_fill_1 FILLER_120_853 ();
 sg13g2_decap_8 FILLER_120_867 ();
 sg13g2_decap_8 FILLER_120_874 ();
 sg13g2_decap_4 FILLER_120_881 ();
 sg13g2_decap_8 FILLER_120_894 ();
 sg13g2_decap_8 FILLER_120_901 ();
 sg13g2_decap_8 FILLER_120_908 ();
 sg13g2_decap_8 FILLER_120_915 ();
 sg13g2_decap_8 FILLER_120_922 ();
 sg13g2_decap_8 FILLER_120_929 ();
 sg13g2_decap_8 FILLER_120_936 ();
 sg13g2_decap_8 FILLER_120_943 ();
 sg13g2_decap_4 FILLER_120_950 ();
 sg13g2_fill_2 FILLER_120_954 ();
 sg13g2_fill_2 FILLER_120_961 ();
 sg13g2_decap_8 FILLER_120_991 ();
 sg13g2_decap_4 FILLER_120_998 ();
 sg13g2_decap_4 FILLER_120_1027 ();
 sg13g2_fill_2 FILLER_120_1031 ();
 sg13g2_fill_2 FILLER_120_1037 ();
 sg13g2_fill_1 FILLER_120_1039 ();
 sg13g2_decap_8 FILLER_120_1062 ();
 sg13g2_fill_2 FILLER_120_1069 ();
 sg13g2_fill_2 FILLER_120_1092 ();
 sg13g2_decap_8 FILLER_120_1102 ();
 sg13g2_fill_2 FILLER_120_1109 ();
 sg13g2_fill_1 FILLER_120_1111 ();
 sg13g2_decap_8 FILLER_120_1120 ();
 sg13g2_decap_8 FILLER_120_1127 ();
 sg13g2_decap_8 FILLER_120_1134 ();
 sg13g2_decap_4 FILLER_120_1141 ();
 sg13g2_decap_8 FILLER_120_1158 ();
 sg13g2_decap_4 FILLER_120_1165 ();
 sg13g2_fill_1 FILLER_120_1169 ();
 sg13g2_decap_8 FILLER_120_1186 ();
 sg13g2_decap_8 FILLER_120_1193 ();
 sg13g2_fill_2 FILLER_120_1200 ();
 sg13g2_fill_1 FILLER_120_1202 ();
 sg13g2_decap_8 FILLER_120_1222 ();
 sg13g2_decap_8 FILLER_120_1229 ();
 sg13g2_decap_4 FILLER_120_1236 ();
 sg13g2_fill_2 FILLER_120_1240 ();
 sg13g2_decap_8 FILLER_120_1254 ();
 sg13g2_decap_8 FILLER_120_1261 ();
 sg13g2_decap_8 FILLER_120_1268 ();
 sg13g2_decap_8 FILLER_120_1275 ();
 sg13g2_decap_4 FILLER_120_1282 ();
 sg13g2_fill_2 FILLER_120_1286 ();
 sg13g2_decap_8 FILLER_120_1301 ();
 sg13g2_decap_8 FILLER_120_1308 ();
 sg13g2_decap_8 FILLER_120_1315 ();
 sg13g2_decap_8 FILLER_120_1322 ();
 sg13g2_decap_8 FILLER_120_1329 ();
 sg13g2_decap_4 FILLER_120_1336 ();
 sg13g2_fill_1 FILLER_120_1340 ();
 sg13g2_decap_8 FILLER_120_1346 ();
 sg13g2_decap_4 FILLER_120_1353 ();
 sg13g2_decap_4 FILLER_120_1365 ();
 sg13g2_fill_2 FILLER_120_1374 ();
 sg13g2_fill_1 FILLER_120_1376 ();
 sg13g2_decap_8 FILLER_120_1384 ();
 sg13g2_decap_8 FILLER_120_1391 ();
 sg13g2_decap_8 FILLER_120_1398 ();
 sg13g2_decap_8 FILLER_120_1405 ();
 sg13g2_decap_8 FILLER_120_1412 ();
 sg13g2_decap_8 FILLER_120_1419 ();
 sg13g2_decap_8 FILLER_120_1426 ();
 sg13g2_decap_8 FILLER_120_1433 ();
 sg13g2_fill_1 FILLER_120_1440 ();
 sg13g2_decap_8 FILLER_120_1449 ();
 sg13g2_decap_8 FILLER_120_1456 ();
 sg13g2_decap_8 FILLER_120_1463 ();
 sg13g2_decap_8 FILLER_120_1470 ();
 sg13g2_decap_8 FILLER_120_1477 ();
 sg13g2_decap_8 FILLER_120_1484 ();
 sg13g2_decap_8 FILLER_120_1491 ();
 sg13g2_decap_8 FILLER_120_1498 ();
 sg13g2_decap_8 FILLER_120_1505 ();
 sg13g2_decap_8 FILLER_120_1512 ();
 sg13g2_decap_4 FILLER_120_1519 ();
 sg13g2_decap_4 FILLER_120_1535 ();
 sg13g2_fill_1 FILLER_120_1539 ();
 sg13g2_decap_8 FILLER_120_1575 ();
 sg13g2_decap_8 FILLER_120_1582 ();
 sg13g2_decap_8 FILLER_120_1589 ();
 sg13g2_decap_8 FILLER_120_1596 ();
 sg13g2_decap_8 FILLER_120_1603 ();
 sg13g2_decap_4 FILLER_120_1610 ();
 sg13g2_fill_1 FILLER_120_1614 ();
 sg13g2_decap_8 FILLER_120_1637 ();
 sg13g2_decap_8 FILLER_120_1644 ();
 sg13g2_decap_8 FILLER_120_1651 ();
 sg13g2_decap_8 FILLER_120_1658 ();
 sg13g2_fill_2 FILLER_120_1665 ();
 sg13g2_fill_1 FILLER_120_1667 ();
 sg13g2_decap_8 FILLER_120_1673 ();
 sg13g2_decap_8 FILLER_120_1680 ();
 sg13g2_fill_2 FILLER_120_1687 ();
 sg13g2_fill_1 FILLER_120_1689 ();
 sg13g2_decap_4 FILLER_120_1695 ();
 sg13g2_fill_2 FILLER_120_1699 ();
 sg13g2_decap_8 FILLER_120_1706 ();
 sg13g2_decap_8 FILLER_120_1713 ();
 sg13g2_decap_8 FILLER_120_1720 ();
 sg13g2_decap_8 FILLER_120_1727 ();
 sg13g2_decap_8 FILLER_120_1734 ();
 sg13g2_decap_8 FILLER_120_1741 ();
 sg13g2_decap_8 FILLER_120_1748 ();
 sg13g2_decap_8 FILLER_120_1755 ();
 sg13g2_decap_4 FILLER_120_1762 ();
 sg13g2_fill_2 FILLER_120_1766 ();
 sg13g2_decap_8 FILLER_121_0 ();
 sg13g2_decap_8 FILLER_121_7 ();
 sg13g2_decap_8 FILLER_121_14 ();
 sg13g2_decap_4 FILLER_121_21 ();
 sg13g2_decap_8 FILLER_121_33 ();
 sg13g2_decap_8 FILLER_121_40 ();
 sg13g2_decap_8 FILLER_121_47 ();
 sg13g2_decap_8 FILLER_121_54 ();
 sg13g2_decap_4 FILLER_121_61 ();
 sg13g2_fill_2 FILLER_121_65 ();
 sg13g2_decap_4 FILLER_121_71 ();
 sg13g2_fill_2 FILLER_121_75 ();
 sg13g2_decap_8 FILLER_121_87 ();
 sg13g2_decap_8 FILLER_121_94 ();
 sg13g2_decap_8 FILLER_121_101 ();
 sg13g2_decap_8 FILLER_121_108 ();
 sg13g2_decap_8 FILLER_121_115 ();
 sg13g2_decap_8 FILLER_121_122 ();
 sg13g2_decap_8 FILLER_121_129 ();
 sg13g2_decap_8 FILLER_121_136 ();
 sg13g2_decap_8 FILLER_121_143 ();
 sg13g2_decap_8 FILLER_121_150 ();
 sg13g2_fill_1 FILLER_121_157 ();
 sg13g2_decap_8 FILLER_121_172 ();
 sg13g2_decap_8 FILLER_121_179 ();
 sg13g2_decap_8 FILLER_121_186 ();
 sg13g2_decap_8 FILLER_121_193 ();
 sg13g2_fill_2 FILLER_121_200 ();
 sg13g2_fill_1 FILLER_121_202 ();
 sg13g2_decap_4 FILLER_121_209 ();
 sg13g2_fill_1 FILLER_121_213 ();
 sg13g2_fill_1 FILLER_121_222 ();
 sg13g2_decap_8 FILLER_121_235 ();
 sg13g2_decap_8 FILLER_121_242 ();
 sg13g2_decap_4 FILLER_121_249 ();
 sg13g2_fill_1 FILLER_121_253 ();
 sg13g2_decap_8 FILLER_121_262 ();
 sg13g2_decap_4 FILLER_121_269 ();
 sg13g2_fill_1 FILLER_121_273 ();
 sg13g2_decap_8 FILLER_121_282 ();
 sg13g2_decap_8 FILLER_121_289 ();
 sg13g2_decap_4 FILLER_121_296 ();
 sg13g2_decap_8 FILLER_121_309 ();
 sg13g2_decap_4 FILLER_121_316 ();
 sg13g2_decap_8 FILLER_121_330 ();
 sg13g2_decap_8 FILLER_121_337 ();
 sg13g2_decap_8 FILLER_121_344 ();
 sg13g2_decap_8 FILLER_121_351 ();
 sg13g2_decap_4 FILLER_121_358 ();
 sg13g2_fill_2 FILLER_121_362 ();
 sg13g2_decap_8 FILLER_121_373 ();
 sg13g2_decap_8 FILLER_121_380 ();
 sg13g2_decap_8 FILLER_121_387 ();
 sg13g2_decap_8 FILLER_121_394 ();
 sg13g2_decap_8 FILLER_121_401 ();
 sg13g2_decap_8 FILLER_121_408 ();
 sg13g2_decap_8 FILLER_121_415 ();
 sg13g2_decap_8 FILLER_121_422 ();
 sg13g2_decap_8 FILLER_121_429 ();
 sg13g2_decap_8 FILLER_121_436 ();
 sg13g2_decap_8 FILLER_121_443 ();
 sg13g2_decap_8 FILLER_121_450 ();
 sg13g2_decap_8 FILLER_121_457 ();
 sg13g2_decap_8 FILLER_121_464 ();
 sg13g2_decap_8 FILLER_121_471 ();
 sg13g2_decap_8 FILLER_121_499 ();
 sg13g2_decap_8 FILLER_121_506 ();
 sg13g2_decap_8 FILLER_121_513 ();
 sg13g2_decap_8 FILLER_121_520 ();
 sg13g2_fill_1 FILLER_121_527 ();
 sg13g2_decap_8 FILLER_121_541 ();
 sg13g2_decap_8 FILLER_121_548 ();
 sg13g2_decap_8 FILLER_121_555 ();
 sg13g2_decap_8 FILLER_121_562 ();
 sg13g2_decap_4 FILLER_121_569 ();
 sg13g2_fill_1 FILLER_121_573 ();
 sg13g2_decap_8 FILLER_121_600 ();
 sg13g2_decap_8 FILLER_121_607 ();
 sg13g2_decap_8 FILLER_121_614 ();
 sg13g2_decap_4 FILLER_121_621 ();
 sg13g2_fill_2 FILLER_121_648 ();
 sg13g2_decap_8 FILLER_121_667 ();
 sg13g2_decap_8 FILLER_121_674 ();
 sg13g2_decap_8 FILLER_121_681 ();
 sg13g2_decap_8 FILLER_121_688 ();
 sg13g2_decap_8 FILLER_121_695 ();
 sg13g2_decap_8 FILLER_121_702 ();
 sg13g2_decap_8 FILLER_121_709 ();
 sg13g2_decap_8 FILLER_121_716 ();
 sg13g2_decap_8 FILLER_121_723 ();
 sg13g2_fill_2 FILLER_121_735 ();
 sg13g2_fill_1 FILLER_121_737 ();
 sg13g2_decap_8 FILLER_121_755 ();
 sg13g2_decap_4 FILLER_121_762 ();
 sg13g2_fill_2 FILLER_121_766 ();
 sg13g2_decap_8 FILLER_121_776 ();
 sg13g2_decap_8 FILLER_121_783 ();
 sg13g2_decap_4 FILLER_121_790 ();
 sg13g2_fill_2 FILLER_121_794 ();
 sg13g2_decap_8 FILLER_121_804 ();
 sg13g2_decap_4 FILLER_121_811 ();
 sg13g2_fill_1 FILLER_121_815 ();
 sg13g2_decap_4 FILLER_121_824 ();
 sg13g2_fill_2 FILLER_121_828 ();
 sg13g2_decap_8 FILLER_121_836 ();
 sg13g2_fill_2 FILLER_121_843 ();
 sg13g2_fill_1 FILLER_121_845 ();
 sg13g2_fill_2 FILLER_121_855 ();
 sg13g2_fill_2 FILLER_121_866 ();
 sg13g2_decap_8 FILLER_121_871 ();
 sg13g2_decap_8 FILLER_121_878 ();
 sg13g2_decap_4 FILLER_121_885 ();
 sg13g2_decap_8 FILLER_121_895 ();
 sg13g2_decap_4 FILLER_121_902 ();
 sg13g2_fill_2 FILLER_121_906 ();
 sg13g2_decap_8 FILLER_121_921 ();
 sg13g2_decap_8 FILLER_121_928 ();
 sg13g2_decap_8 FILLER_121_935 ();
 sg13g2_decap_8 FILLER_121_942 ();
 sg13g2_fill_2 FILLER_121_978 ();
 sg13g2_decap_8 FILLER_121_989 ();
 sg13g2_decap_8 FILLER_121_996 ();
 sg13g2_decap_8 FILLER_121_1003 ();
 sg13g2_decap_8 FILLER_121_1010 ();
 sg13g2_decap_8 FILLER_121_1017 ();
 sg13g2_decap_8 FILLER_121_1024 ();
 sg13g2_decap_8 FILLER_121_1031 ();
 sg13g2_decap_8 FILLER_121_1038 ();
 sg13g2_decap_8 FILLER_121_1045 ();
 sg13g2_decap_8 FILLER_121_1052 ();
 sg13g2_decap_8 FILLER_121_1059 ();
 sg13g2_decap_8 FILLER_121_1066 ();
 sg13g2_decap_4 FILLER_121_1073 ();
 sg13g2_fill_2 FILLER_121_1077 ();
 sg13g2_decap_4 FILLER_121_1092 ();
 sg13g2_fill_1 FILLER_121_1096 ();
 sg13g2_decap_8 FILLER_121_1112 ();
 sg13g2_decap_8 FILLER_121_1119 ();
 sg13g2_decap_8 FILLER_121_1126 ();
 sg13g2_decap_8 FILLER_121_1133 ();
 sg13g2_decap_8 FILLER_121_1140 ();
 sg13g2_decap_8 FILLER_121_1147 ();
 sg13g2_decap_8 FILLER_121_1154 ();
 sg13g2_decap_8 FILLER_121_1161 ();
 sg13g2_decap_8 FILLER_121_1168 ();
 sg13g2_decap_8 FILLER_121_1180 ();
 sg13g2_fill_1 FILLER_121_1187 ();
 sg13g2_decap_8 FILLER_121_1201 ();
 sg13g2_decap_4 FILLER_121_1208 ();
 sg13g2_fill_2 FILLER_121_1212 ();
 sg13g2_decap_4 FILLER_121_1235 ();
 sg13g2_decap_8 FILLER_121_1247 ();
 sg13g2_decap_8 FILLER_121_1254 ();
 sg13g2_decap_4 FILLER_121_1261 ();
 sg13g2_fill_2 FILLER_121_1265 ();
 sg13g2_decap_8 FILLER_121_1272 ();
 sg13g2_decap_8 FILLER_121_1279 ();
 sg13g2_decap_8 FILLER_121_1286 ();
 sg13g2_decap_8 FILLER_121_1293 ();
 sg13g2_decap_4 FILLER_121_1300 ();
 sg13g2_fill_1 FILLER_121_1304 ();
 sg13g2_decap_8 FILLER_121_1310 ();
 sg13g2_decap_8 FILLER_121_1317 ();
 sg13g2_decap_8 FILLER_121_1324 ();
 sg13g2_decap_4 FILLER_121_1331 ();
 sg13g2_fill_2 FILLER_121_1335 ();
 sg13g2_decap_8 FILLER_121_1352 ();
 sg13g2_decap_8 FILLER_121_1359 ();
 sg13g2_decap_8 FILLER_121_1366 ();
 sg13g2_decap_4 FILLER_121_1373 ();
 sg13g2_decap_8 FILLER_121_1388 ();
 sg13g2_decap_8 FILLER_121_1395 ();
 sg13g2_decap_8 FILLER_121_1402 ();
 sg13g2_decap_8 FILLER_121_1409 ();
 sg13g2_decap_4 FILLER_121_1416 ();
 sg13g2_fill_2 FILLER_121_1420 ();
 sg13g2_fill_2 FILLER_121_1431 ();
 sg13g2_fill_1 FILLER_121_1433 ();
 sg13g2_fill_2 FILLER_121_1442 ();
 sg13g2_fill_1 FILLER_121_1444 ();
 sg13g2_decap_8 FILLER_121_1449 ();
 sg13g2_decap_8 FILLER_121_1456 ();
 sg13g2_decap_8 FILLER_121_1463 ();
 sg13g2_decap_8 FILLER_121_1470 ();
 sg13g2_decap_4 FILLER_121_1477 ();
 sg13g2_fill_1 FILLER_121_1481 ();
 sg13g2_decap_8 FILLER_121_1487 ();
 sg13g2_decap_8 FILLER_121_1494 ();
 sg13g2_decap_8 FILLER_121_1501 ();
 sg13g2_decap_8 FILLER_121_1508 ();
 sg13g2_decap_8 FILLER_121_1515 ();
 sg13g2_decap_8 FILLER_121_1522 ();
 sg13g2_decap_4 FILLER_121_1529 ();
 sg13g2_fill_2 FILLER_121_1533 ();
 sg13g2_decap_8 FILLER_121_1543 ();
 sg13g2_fill_2 FILLER_121_1550 ();
 sg13g2_fill_1 FILLER_121_1555 ();
 sg13g2_decap_4 FILLER_121_1560 ();
 sg13g2_decap_8 FILLER_121_1576 ();
 sg13g2_decap_8 FILLER_121_1583 ();
 sg13g2_decap_8 FILLER_121_1590 ();
 sg13g2_decap_8 FILLER_121_1597 ();
 sg13g2_decap_8 FILLER_121_1613 ();
 sg13g2_decap_4 FILLER_121_1620 ();
 sg13g2_decap_8 FILLER_121_1630 ();
 sg13g2_decap_8 FILLER_121_1637 ();
 sg13g2_decap_4 FILLER_121_1644 ();
 sg13g2_decap_8 FILLER_121_1657 ();
 sg13g2_decap_8 FILLER_121_1664 ();
 sg13g2_decap_8 FILLER_121_1671 ();
 sg13g2_decap_8 FILLER_121_1678 ();
 sg13g2_decap_8 FILLER_121_1685 ();
 sg13g2_decap_8 FILLER_121_1692 ();
 sg13g2_decap_8 FILLER_121_1699 ();
 sg13g2_decap_8 FILLER_121_1706 ();
 sg13g2_decap_4 FILLER_121_1717 ();
 sg13g2_decap_8 FILLER_121_1726 ();
 sg13g2_decap_8 FILLER_121_1733 ();
 sg13g2_decap_8 FILLER_121_1740 ();
 sg13g2_decap_8 FILLER_121_1747 ();
 sg13g2_decap_8 FILLER_121_1754 ();
 sg13g2_decap_8 FILLER_121_1761 ();
 sg13g2_decap_8 FILLER_122_0 ();
 sg13g2_decap_8 FILLER_122_7 ();
 sg13g2_decap_8 FILLER_122_14 ();
 sg13g2_decap_8 FILLER_122_21 ();
 sg13g2_decap_4 FILLER_122_28 ();
 sg13g2_decap_8 FILLER_122_40 ();
 sg13g2_decap_8 FILLER_122_47 ();
 sg13g2_fill_2 FILLER_122_54 ();
 sg13g2_fill_1 FILLER_122_56 ();
 sg13g2_decap_8 FILLER_122_77 ();
 sg13g2_decap_4 FILLER_122_84 ();
 sg13g2_decap_8 FILLER_122_92 ();
 sg13g2_decap_8 FILLER_122_99 ();
 sg13g2_decap_8 FILLER_122_106 ();
 sg13g2_fill_2 FILLER_122_113 ();
 sg13g2_decap_8 FILLER_122_132 ();
 sg13g2_decap_8 FILLER_122_139 ();
 sg13g2_decap_8 FILLER_122_146 ();
 sg13g2_decap_8 FILLER_122_153 ();
 sg13g2_decap_8 FILLER_122_160 ();
 sg13g2_decap_8 FILLER_122_167 ();
 sg13g2_decap_8 FILLER_122_174 ();
 sg13g2_decap_8 FILLER_122_181 ();
 sg13g2_decap_8 FILLER_122_188 ();
 sg13g2_decap_8 FILLER_122_195 ();
 sg13g2_decap_8 FILLER_122_202 ();
 sg13g2_decap_8 FILLER_122_209 ();
 sg13g2_decap_8 FILLER_122_216 ();
 sg13g2_decap_8 FILLER_122_223 ();
 sg13g2_decap_8 FILLER_122_230 ();
 sg13g2_decap_8 FILLER_122_237 ();
 sg13g2_fill_1 FILLER_122_244 ();
 sg13g2_decap_8 FILLER_122_258 ();
 sg13g2_decap_8 FILLER_122_265 ();
 sg13g2_decap_8 FILLER_122_272 ();
 sg13g2_decap_8 FILLER_122_279 ();
 sg13g2_decap_8 FILLER_122_286 ();
 sg13g2_decap_8 FILLER_122_293 ();
 sg13g2_decap_8 FILLER_122_300 ();
 sg13g2_decap_8 FILLER_122_307 ();
 sg13g2_decap_8 FILLER_122_314 ();
 sg13g2_decap_8 FILLER_122_321 ();
 sg13g2_decap_8 FILLER_122_328 ();
 sg13g2_decap_8 FILLER_122_335 ();
 sg13g2_decap_4 FILLER_122_342 ();
 sg13g2_fill_2 FILLER_122_346 ();
 sg13g2_decap_8 FILLER_122_357 ();
 sg13g2_fill_1 FILLER_122_364 ();
 sg13g2_fill_2 FILLER_122_384 ();
 sg13g2_fill_1 FILLER_122_386 ();
 sg13g2_decap_8 FILLER_122_419 ();
 sg13g2_decap_8 FILLER_122_426 ();
 sg13g2_decap_8 FILLER_122_433 ();
 sg13g2_decap_8 FILLER_122_440 ();
 sg13g2_decap_8 FILLER_122_447 ();
 sg13g2_fill_1 FILLER_122_454 ();
 sg13g2_decap_8 FILLER_122_459 ();
 sg13g2_decap_4 FILLER_122_466 ();
 sg13g2_fill_1 FILLER_122_470 ();
 sg13g2_fill_1 FILLER_122_486 ();
 sg13g2_decap_4 FILLER_122_497 ();
 sg13g2_fill_2 FILLER_122_501 ();
 sg13g2_decap_8 FILLER_122_511 ();
 sg13g2_decap_8 FILLER_122_518 ();
 sg13g2_decap_8 FILLER_122_525 ();
 sg13g2_decap_8 FILLER_122_532 ();
 sg13g2_decap_8 FILLER_122_539 ();
 sg13g2_decap_8 FILLER_122_546 ();
 sg13g2_decap_8 FILLER_122_553 ();
 sg13g2_decap_8 FILLER_122_560 ();
 sg13g2_decap_8 FILLER_122_567 ();
 sg13g2_decap_8 FILLER_122_574 ();
 sg13g2_decap_8 FILLER_122_593 ();
 sg13g2_decap_8 FILLER_122_600 ();
 sg13g2_decap_8 FILLER_122_607 ();
 sg13g2_decap_8 FILLER_122_614 ();
 sg13g2_decap_8 FILLER_122_621 ();
 sg13g2_decap_4 FILLER_122_628 ();
 sg13g2_fill_1 FILLER_122_632 ();
 sg13g2_decap_8 FILLER_122_666 ();
 sg13g2_decap_8 FILLER_122_673 ();
 sg13g2_decap_8 FILLER_122_680 ();
 sg13g2_decap_8 FILLER_122_687 ();
 sg13g2_decap_8 FILLER_122_694 ();
 sg13g2_decap_8 FILLER_122_701 ();
 sg13g2_decap_8 FILLER_122_708 ();
 sg13g2_decap_4 FILLER_122_715 ();
 sg13g2_decap_8 FILLER_122_727 ();
 sg13g2_decap_8 FILLER_122_734 ();
 sg13g2_fill_1 FILLER_122_741 ();
 sg13g2_decap_8 FILLER_122_757 ();
 sg13g2_decap_8 FILLER_122_764 ();
 sg13g2_decap_8 FILLER_122_771 ();
 sg13g2_decap_8 FILLER_122_778 ();
 sg13g2_decap_8 FILLER_122_785 ();
 sg13g2_decap_8 FILLER_122_792 ();
 sg13g2_decap_8 FILLER_122_799 ();
 sg13g2_decap_8 FILLER_122_806 ();
 sg13g2_decap_4 FILLER_122_813 ();
 sg13g2_fill_2 FILLER_122_817 ();
 sg13g2_decap_8 FILLER_122_825 ();
 sg13g2_decap_8 FILLER_122_832 ();
 sg13g2_decap_8 FILLER_122_839 ();
 sg13g2_decap_8 FILLER_122_851 ();
 sg13g2_fill_2 FILLER_122_858 ();
 sg13g2_decap_4 FILLER_122_864 ();
 sg13g2_decap_8 FILLER_122_876 ();
 sg13g2_decap_8 FILLER_122_883 ();
 sg13g2_decap_8 FILLER_122_890 ();
 sg13g2_decap_8 FILLER_122_897 ();
 sg13g2_fill_2 FILLER_122_904 ();
 sg13g2_fill_1 FILLER_122_906 ();
 sg13g2_decap_8 FILLER_122_911 ();
 sg13g2_decap_8 FILLER_122_918 ();
 sg13g2_decap_8 FILLER_122_925 ();
 sg13g2_decap_8 FILLER_122_932 ();
 sg13g2_decap_8 FILLER_122_939 ();
 sg13g2_decap_8 FILLER_122_946 ();
 sg13g2_decap_4 FILLER_122_953 ();
 sg13g2_fill_1 FILLER_122_957 ();
 sg13g2_decap_8 FILLER_122_966 ();
 sg13g2_decap_8 FILLER_122_973 ();
 sg13g2_decap_4 FILLER_122_980 ();
 sg13g2_fill_2 FILLER_122_984 ();
 sg13g2_decap_8 FILLER_122_1012 ();
 sg13g2_decap_8 FILLER_122_1019 ();
 sg13g2_decap_8 FILLER_122_1026 ();
 sg13g2_fill_2 FILLER_122_1033 ();
 sg13g2_decap_8 FILLER_122_1043 ();
 sg13g2_decap_8 FILLER_122_1050 ();
 sg13g2_decap_8 FILLER_122_1057 ();
 sg13g2_decap_8 FILLER_122_1064 ();
 sg13g2_decap_8 FILLER_122_1071 ();
 sg13g2_decap_8 FILLER_122_1078 ();
 sg13g2_decap_8 FILLER_122_1085 ();
 sg13g2_decap_4 FILLER_122_1092 ();
 sg13g2_fill_1 FILLER_122_1096 ();
 sg13g2_decap_8 FILLER_122_1120 ();
 sg13g2_decap_8 FILLER_122_1127 ();
 sg13g2_decap_8 FILLER_122_1134 ();
 sg13g2_decap_8 FILLER_122_1141 ();
 sg13g2_decap_8 FILLER_122_1148 ();
 sg13g2_decap_8 FILLER_122_1155 ();
 sg13g2_decap_8 FILLER_122_1162 ();
 sg13g2_decap_8 FILLER_122_1169 ();
 sg13g2_decap_8 FILLER_122_1176 ();
 sg13g2_decap_8 FILLER_122_1183 ();
 sg13g2_decap_4 FILLER_122_1190 ();
 sg13g2_fill_2 FILLER_122_1194 ();
 sg13g2_decap_8 FILLER_122_1201 ();
 sg13g2_decap_8 FILLER_122_1208 ();
 sg13g2_decap_8 FILLER_122_1215 ();
 sg13g2_decap_8 FILLER_122_1222 ();
 sg13g2_decap_8 FILLER_122_1229 ();
 sg13g2_decap_8 FILLER_122_1236 ();
 sg13g2_decap_8 FILLER_122_1243 ();
 sg13g2_decap_8 FILLER_122_1254 ();
 sg13g2_decap_8 FILLER_122_1261 ();
 sg13g2_decap_8 FILLER_122_1268 ();
 sg13g2_decap_8 FILLER_122_1275 ();
 sg13g2_decap_8 FILLER_122_1282 ();
 sg13g2_decap_8 FILLER_122_1289 ();
 sg13g2_decap_8 FILLER_122_1296 ();
 sg13g2_fill_2 FILLER_122_1303 ();
 sg13g2_fill_1 FILLER_122_1305 ();
 sg13g2_fill_2 FILLER_122_1314 ();
 sg13g2_decap_8 FILLER_122_1329 ();
 sg13g2_decap_8 FILLER_122_1336 ();
 sg13g2_decap_8 FILLER_122_1343 ();
 sg13g2_decap_8 FILLER_122_1350 ();
 sg13g2_decap_8 FILLER_122_1357 ();
 sg13g2_fill_1 FILLER_122_1364 ();
 sg13g2_fill_1 FILLER_122_1369 ();
 sg13g2_decap_8 FILLER_122_1388 ();
 sg13g2_decap_8 FILLER_122_1395 ();
 sg13g2_decap_4 FILLER_122_1402 ();
 sg13g2_fill_2 FILLER_122_1406 ();
 sg13g2_decap_4 FILLER_122_1416 ();
 sg13g2_fill_1 FILLER_122_1420 ();
 sg13g2_decap_4 FILLER_122_1426 ();
 sg13g2_decap_8 FILLER_122_1459 ();
 sg13g2_decap_8 FILLER_122_1466 ();
 sg13g2_decap_8 FILLER_122_1473 ();
 sg13g2_decap_4 FILLER_122_1480 ();
 sg13g2_fill_2 FILLER_122_1484 ();
 sg13g2_fill_1 FILLER_122_1491 ();
 sg13g2_decap_8 FILLER_122_1496 ();
 sg13g2_decap_8 FILLER_122_1503 ();
 sg13g2_decap_8 FILLER_122_1510 ();
 sg13g2_decap_8 FILLER_122_1517 ();
 sg13g2_decap_4 FILLER_122_1524 ();
 sg13g2_fill_2 FILLER_122_1528 ();
 sg13g2_decap_8 FILLER_122_1534 ();
 sg13g2_decap_8 FILLER_122_1541 ();
 sg13g2_decap_8 FILLER_122_1548 ();
 sg13g2_fill_1 FILLER_122_1555 ();
 sg13g2_fill_1 FILLER_122_1559 ();
 sg13g2_decap_8 FILLER_122_1573 ();
 sg13g2_decap_8 FILLER_122_1580 ();
 sg13g2_decap_8 FILLER_122_1587 ();
 sg13g2_decap_8 FILLER_122_1594 ();
 sg13g2_decap_8 FILLER_122_1601 ();
 sg13g2_decap_8 FILLER_122_1608 ();
 sg13g2_decap_8 FILLER_122_1615 ();
 sg13g2_decap_8 FILLER_122_1622 ();
 sg13g2_decap_8 FILLER_122_1629 ();
 sg13g2_decap_8 FILLER_122_1646 ();
 sg13g2_decap_8 FILLER_122_1653 ();
 sg13g2_decap_4 FILLER_122_1660 ();
 sg13g2_decap_8 FILLER_122_1672 ();
 sg13g2_decap_8 FILLER_122_1679 ();
 sg13g2_decap_8 FILLER_122_1686 ();
 sg13g2_decap_8 FILLER_122_1693 ();
 sg13g2_decap_8 FILLER_122_1700 ();
 sg13g2_decap_8 FILLER_122_1707 ();
 sg13g2_decap_8 FILLER_122_1714 ();
 sg13g2_fill_2 FILLER_122_1721 ();
 sg13g2_fill_2 FILLER_122_1727 ();
 sg13g2_fill_1 FILLER_122_1729 ();
 sg13g2_decap_8 FILLER_122_1738 ();
 sg13g2_decap_8 FILLER_122_1745 ();
 sg13g2_decap_8 FILLER_122_1752 ();
 sg13g2_decap_8 FILLER_122_1759 ();
 sg13g2_fill_2 FILLER_122_1766 ();
 sg13g2_decap_8 FILLER_123_0 ();
 sg13g2_decap_8 FILLER_123_7 ();
 sg13g2_decap_8 FILLER_123_14 ();
 sg13g2_decap_4 FILLER_123_21 ();
 sg13g2_fill_2 FILLER_123_25 ();
 sg13g2_decap_8 FILLER_123_46 ();
 sg13g2_decap_4 FILLER_123_53 ();
 sg13g2_fill_1 FILLER_123_57 ();
 sg13g2_fill_2 FILLER_123_66 ();
 sg13g2_fill_1 FILLER_123_68 ();
 sg13g2_decap_4 FILLER_123_77 ();
 sg13g2_fill_2 FILLER_123_81 ();
 sg13g2_decap_4 FILLER_123_95 ();
 sg13g2_fill_2 FILLER_123_99 ();
 sg13g2_decap_8 FILLER_123_110 ();
 sg13g2_fill_2 FILLER_123_117 ();
 sg13g2_fill_1 FILLER_123_119 ();
 sg13g2_decap_8 FILLER_123_125 ();
 sg13g2_decap_8 FILLER_123_132 ();
 sg13g2_decap_8 FILLER_123_139 ();
 sg13g2_decap_4 FILLER_123_146 ();
 sg13g2_decap_8 FILLER_123_163 ();
 sg13g2_decap_8 FILLER_123_191 ();
 sg13g2_decap_8 FILLER_123_198 ();
 sg13g2_decap_8 FILLER_123_205 ();
 sg13g2_fill_2 FILLER_123_212 ();
 sg13g2_decap_4 FILLER_123_222 ();
 sg13g2_fill_2 FILLER_123_234 ();
 sg13g2_decap_8 FILLER_123_252 ();
 sg13g2_decap_8 FILLER_123_259 ();
 sg13g2_decap_8 FILLER_123_266 ();
 sg13g2_decap_8 FILLER_123_273 ();
 sg13g2_decap_8 FILLER_123_280 ();
 sg13g2_decap_4 FILLER_123_287 ();
 sg13g2_decap_8 FILLER_123_296 ();
 sg13g2_decap_8 FILLER_123_303 ();
 sg13g2_decap_4 FILLER_123_310 ();
 sg13g2_fill_1 FILLER_123_314 ();
 sg13g2_decap_8 FILLER_123_325 ();
 sg13g2_decap_8 FILLER_123_332 ();
 sg13g2_fill_1 FILLER_123_339 ();
 sg13g2_fill_2 FILLER_123_348 ();
 sg13g2_fill_1 FILLER_123_350 ();
 sg13g2_decap_8 FILLER_123_361 ();
 sg13g2_decap_8 FILLER_123_368 ();
 sg13g2_decap_4 FILLER_123_375 ();
 sg13g2_fill_1 FILLER_123_379 ();
 sg13g2_decap_8 FILLER_123_409 ();
 sg13g2_decap_8 FILLER_123_416 ();
 sg13g2_decap_8 FILLER_123_423 ();
 sg13g2_decap_8 FILLER_123_430 ();
 sg13g2_decap_8 FILLER_123_437 ();
 sg13g2_decap_8 FILLER_123_444 ();
 sg13g2_decap_8 FILLER_123_451 ();
 sg13g2_decap_8 FILLER_123_458 ();
 sg13g2_decap_8 FILLER_123_465 ();
 sg13g2_decap_4 FILLER_123_472 ();
 sg13g2_fill_2 FILLER_123_476 ();
 sg13g2_decap_8 FILLER_123_491 ();
 sg13g2_decap_4 FILLER_123_498 ();
 sg13g2_fill_1 FILLER_123_502 ();
 sg13g2_decap_8 FILLER_123_507 ();
 sg13g2_decap_8 FILLER_123_514 ();
 sg13g2_decap_8 FILLER_123_521 ();
 sg13g2_decap_8 FILLER_123_528 ();
 sg13g2_decap_8 FILLER_123_535 ();
 sg13g2_decap_8 FILLER_123_542 ();
 sg13g2_decap_8 FILLER_123_549 ();
 sg13g2_decap_4 FILLER_123_556 ();
 sg13g2_decap_4 FILLER_123_576 ();
 sg13g2_fill_2 FILLER_123_580 ();
 sg13g2_decap_8 FILLER_123_591 ();
 sg13g2_decap_8 FILLER_123_598 ();
 sg13g2_fill_1 FILLER_123_605 ();
 sg13g2_decap_8 FILLER_123_611 ();
 sg13g2_decap_8 FILLER_123_618 ();
 sg13g2_decap_8 FILLER_123_625 ();
 sg13g2_decap_8 FILLER_123_642 ();
 sg13g2_fill_2 FILLER_123_649 ();
 sg13g2_fill_1 FILLER_123_651 ();
 sg13g2_fill_1 FILLER_123_657 ();
 sg13g2_decap_8 FILLER_123_662 ();
 sg13g2_decap_8 FILLER_123_669 ();
 sg13g2_decap_8 FILLER_123_676 ();
 sg13g2_decap_8 FILLER_123_683 ();
 sg13g2_decap_8 FILLER_123_690 ();
 sg13g2_decap_8 FILLER_123_697 ();
 sg13g2_fill_2 FILLER_123_704 ();
 sg13g2_decap_8 FILLER_123_729 ();
 sg13g2_decap_8 FILLER_123_736 ();
 sg13g2_decap_8 FILLER_123_743 ();
 sg13g2_decap_8 FILLER_123_750 ();
 sg13g2_decap_8 FILLER_123_767 ();
 sg13g2_fill_2 FILLER_123_774 ();
 sg13g2_fill_1 FILLER_123_776 ();
 sg13g2_decap_8 FILLER_123_793 ();
 sg13g2_decap_8 FILLER_123_800 ();
 sg13g2_fill_1 FILLER_123_807 ();
 sg13g2_decap_8 FILLER_123_830 ();
 sg13g2_decap_8 FILLER_123_837 ();
 sg13g2_decap_8 FILLER_123_844 ();
 sg13g2_fill_1 FILLER_123_851 ();
 sg13g2_fill_1 FILLER_123_859 ();
 sg13g2_decap_8 FILLER_123_863 ();
 sg13g2_fill_2 FILLER_123_870 ();
 sg13g2_decap_8 FILLER_123_885 ();
 sg13g2_decap_8 FILLER_123_892 ();
 sg13g2_fill_2 FILLER_123_899 ();
 sg13g2_fill_1 FILLER_123_901 ();
 sg13g2_decap_8 FILLER_123_940 ();
 sg13g2_decap_8 FILLER_123_947 ();
 sg13g2_decap_8 FILLER_123_954 ();
 sg13g2_decap_8 FILLER_123_961 ();
 sg13g2_decap_8 FILLER_123_968 ();
 sg13g2_decap_8 FILLER_123_975 ();
 sg13g2_decap_8 FILLER_123_982 ();
 sg13g2_decap_8 FILLER_123_989 ();
 sg13g2_fill_1 FILLER_123_996 ();
 sg13g2_decap_4 FILLER_123_1001 ();
 sg13g2_fill_1 FILLER_123_1005 ();
 sg13g2_decap_8 FILLER_123_1019 ();
 sg13g2_decap_8 FILLER_123_1026 ();
 sg13g2_decap_8 FILLER_123_1033 ();
 sg13g2_decap_8 FILLER_123_1040 ();
 sg13g2_fill_2 FILLER_123_1047 ();
 sg13g2_fill_2 FILLER_123_1057 ();
 sg13g2_fill_2 FILLER_123_1064 ();
 sg13g2_fill_1 FILLER_123_1066 ();
 sg13g2_decap_8 FILLER_123_1080 ();
 sg13g2_decap_8 FILLER_123_1087 ();
 sg13g2_decap_8 FILLER_123_1094 ();
 sg13g2_decap_8 FILLER_123_1101 ();
 sg13g2_decap_8 FILLER_123_1108 ();
 sg13g2_decap_4 FILLER_123_1115 ();
 sg13g2_decap_8 FILLER_123_1125 ();
 sg13g2_decap_8 FILLER_123_1132 ();
 sg13g2_decap_8 FILLER_123_1139 ();
 sg13g2_decap_8 FILLER_123_1146 ();
 sg13g2_decap_8 FILLER_123_1153 ();
 sg13g2_decap_8 FILLER_123_1160 ();
 sg13g2_fill_1 FILLER_123_1167 ();
 sg13g2_decap_8 FILLER_123_1173 ();
 sg13g2_fill_2 FILLER_123_1180 ();
 sg13g2_fill_1 FILLER_123_1182 ();
 sg13g2_fill_2 FILLER_123_1192 ();
 sg13g2_decap_8 FILLER_123_1202 ();
 sg13g2_fill_2 FILLER_123_1209 ();
 sg13g2_decap_8 FILLER_123_1219 ();
 sg13g2_decap_8 FILLER_123_1226 ();
 sg13g2_decap_8 FILLER_123_1233 ();
 sg13g2_decap_8 FILLER_123_1240 ();
 sg13g2_decap_4 FILLER_123_1247 ();
 sg13g2_fill_2 FILLER_123_1251 ();
 sg13g2_decap_8 FILLER_123_1261 ();
 sg13g2_decap_8 FILLER_123_1268 ();
 sg13g2_decap_8 FILLER_123_1275 ();
 sg13g2_decap_8 FILLER_123_1282 ();
 sg13g2_fill_1 FILLER_123_1289 ();
 sg13g2_decap_8 FILLER_123_1296 ();
 sg13g2_decap_8 FILLER_123_1303 ();
 sg13g2_decap_8 FILLER_123_1310 ();
 sg13g2_fill_2 FILLER_123_1317 ();
 sg13g2_decap_8 FILLER_123_1325 ();
 sg13g2_decap_4 FILLER_123_1332 ();
 sg13g2_fill_1 FILLER_123_1336 ();
 sg13g2_decap_8 FILLER_123_1341 ();
 sg13g2_decap_8 FILLER_123_1348 ();
 sg13g2_decap_4 FILLER_123_1355 ();
 sg13g2_fill_1 FILLER_123_1368 ();
 sg13g2_decap_8 FILLER_123_1398 ();
 sg13g2_decap_8 FILLER_123_1405 ();
 sg13g2_decap_4 FILLER_123_1412 ();
 sg13g2_fill_1 FILLER_123_1416 ();
 sg13g2_fill_2 FILLER_123_1440 ();
 sg13g2_decap_4 FILLER_123_1447 ();
 sg13g2_fill_1 FILLER_123_1451 ();
 sg13g2_decap_8 FILLER_123_1460 ();
 sg13g2_fill_1 FILLER_123_1467 ();
 sg13g2_decap_8 FILLER_123_1476 ();
 sg13g2_fill_1 FILLER_123_1483 ();
 sg13g2_decap_8 FILLER_123_1508 ();
 sg13g2_decap_8 FILLER_123_1515 ();
 sg13g2_fill_2 FILLER_123_1522 ();
 sg13g2_fill_2 FILLER_123_1532 ();
 sg13g2_fill_1 FILLER_123_1534 ();
 sg13g2_decap_8 FILLER_123_1543 ();
 sg13g2_decap_8 FILLER_123_1550 ();
 sg13g2_decap_8 FILLER_123_1557 ();
 sg13g2_decap_8 FILLER_123_1564 ();
 sg13g2_decap_8 FILLER_123_1571 ();
 sg13g2_decap_8 FILLER_123_1578 ();
 sg13g2_decap_8 FILLER_123_1585 ();
 sg13g2_decap_8 FILLER_123_1592 ();
 sg13g2_fill_2 FILLER_123_1599 ();
 sg13g2_fill_1 FILLER_123_1601 ();
 sg13g2_fill_1 FILLER_123_1605 ();
 sg13g2_fill_1 FILLER_123_1610 ();
 sg13g2_decap_8 FILLER_123_1619 ();
 sg13g2_decap_8 FILLER_123_1626 ();
 sg13g2_decap_8 FILLER_123_1633 ();
 sg13g2_fill_1 FILLER_123_1640 ();
 sg13g2_fill_1 FILLER_123_1649 ();
 sg13g2_decap_4 FILLER_123_1663 ();
 sg13g2_fill_1 FILLER_123_1667 ();
 sg13g2_fill_1 FILLER_123_1678 ();
 sg13g2_decap_8 FILLER_123_1687 ();
 sg13g2_decap_8 FILLER_123_1694 ();
 sg13g2_decap_8 FILLER_123_1701 ();
 sg13g2_decap_8 FILLER_123_1708 ();
 sg13g2_fill_2 FILLER_123_1715 ();
 sg13g2_fill_2 FILLER_123_1741 ();
 sg13g2_fill_1 FILLER_123_1743 ();
 sg13g2_decap_8 FILLER_123_1755 ();
 sg13g2_decap_4 FILLER_123_1762 ();
 sg13g2_fill_2 FILLER_123_1766 ();
 sg13g2_decap_8 FILLER_124_0 ();
 sg13g2_decap_8 FILLER_124_7 ();
 sg13g2_decap_8 FILLER_124_14 ();
 sg13g2_decap_4 FILLER_124_21 ();
 sg13g2_fill_2 FILLER_124_25 ();
 sg13g2_decap_8 FILLER_124_53 ();
 sg13g2_decap_8 FILLER_124_60 ();
 sg13g2_decap_8 FILLER_124_67 ();
 sg13g2_decap_8 FILLER_124_74 ();
 sg13g2_decap_8 FILLER_124_81 ();
 sg13g2_decap_4 FILLER_124_88 ();
 sg13g2_fill_2 FILLER_124_96 ();
 sg13g2_decap_8 FILLER_124_122 ();
 sg13g2_decap_8 FILLER_124_129 ();
 sg13g2_decap_8 FILLER_124_136 ();
 sg13g2_decap_8 FILLER_124_143 ();
 sg13g2_fill_2 FILLER_124_166 ();
 sg13g2_fill_1 FILLER_124_168 ();
 sg13g2_decap_8 FILLER_124_173 ();
 sg13g2_decap_8 FILLER_124_180 ();
 sg13g2_decap_4 FILLER_124_187 ();
 sg13g2_fill_2 FILLER_124_191 ();
 sg13g2_decap_4 FILLER_124_199 ();
 sg13g2_fill_1 FILLER_124_203 ();
 sg13g2_decap_8 FILLER_124_209 ();
 sg13g2_decap_8 FILLER_124_216 ();
 sg13g2_decap_8 FILLER_124_223 ();
 sg13g2_decap_4 FILLER_124_230 ();
 sg13g2_fill_1 FILLER_124_234 ();
 sg13g2_decap_4 FILLER_124_241 ();
 sg13g2_fill_2 FILLER_124_245 ();
 sg13g2_decap_8 FILLER_124_252 ();
 sg13g2_decap_8 FILLER_124_259 ();
 sg13g2_decap_4 FILLER_124_266 ();
 sg13g2_fill_2 FILLER_124_270 ();
 sg13g2_decap_8 FILLER_124_292 ();
 sg13g2_decap_8 FILLER_124_299 ();
 sg13g2_decap_4 FILLER_124_306 ();
 sg13g2_decap_8 FILLER_124_318 ();
 sg13g2_decap_4 FILLER_124_325 ();
 sg13g2_decap_8 FILLER_124_342 ();
 sg13g2_fill_2 FILLER_124_349 ();
 sg13g2_fill_1 FILLER_124_351 ();
 sg13g2_decap_8 FILLER_124_361 ();
 sg13g2_decap_8 FILLER_124_368 ();
 sg13g2_decap_8 FILLER_124_375 ();
 sg13g2_decap_4 FILLER_124_382 ();
 sg13g2_fill_2 FILLER_124_386 ();
 sg13g2_decap_8 FILLER_124_395 ();
 sg13g2_decap_8 FILLER_124_402 ();
 sg13g2_decap_8 FILLER_124_409 ();
 sg13g2_decap_8 FILLER_124_416 ();
 sg13g2_decap_4 FILLER_124_423 ();
 sg13g2_fill_2 FILLER_124_427 ();
 sg13g2_fill_2 FILLER_124_436 ();
 sg13g2_decap_8 FILLER_124_454 ();
 sg13g2_decap_8 FILLER_124_461 ();
 sg13g2_fill_1 FILLER_124_468 ();
 sg13g2_decap_8 FILLER_124_474 ();
 sg13g2_decap_8 FILLER_124_481 ();
 sg13g2_fill_1 FILLER_124_488 ();
 sg13g2_fill_2 FILLER_124_499 ();
 sg13g2_decap_8 FILLER_124_514 ();
 sg13g2_decap_8 FILLER_124_521 ();
 sg13g2_decap_8 FILLER_124_528 ();
 sg13g2_decap_8 FILLER_124_535 ();
 sg13g2_decap_8 FILLER_124_547 ();
 sg13g2_decap_8 FILLER_124_554 ();
 sg13g2_decap_4 FILLER_124_561 ();
 sg13g2_fill_1 FILLER_124_565 ();
 sg13g2_decap_4 FILLER_124_575 ();
 sg13g2_decap_8 FILLER_124_596 ();
 sg13g2_decap_8 FILLER_124_603 ();
 sg13g2_decap_8 FILLER_124_610 ();
 sg13g2_decap_8 FILLER_124_617 ();
 sg13g2_decap_8 FILLER_124_624 ();
 sg13g2_decap_8 FILLER_124_639 ();
 sg13g2_decap_8 FILLER_124_646 ();
 sg13g2_decap_8 FILLER_124_653 ();
 sg13g2_decap_8 FILLER_124_660 ();
 sg13g2_decap_8 FILLER_124_667 ();
 sg13g2_decap_8 FILLER_124_674 ();
 sg13g2_fill_1 FILLER_124_681 ();
 sg13g2_fill_2 FILLER_124_687 ();
 sg13g2_fill_1 FILLER_124_689 ();
 sg13g2_fill_1 FILLER_124_699 ();
 sg13g2_decap_4 FILLER_124_709 ();
 sg13g2_fill_2 FILLER_124_713 ();
 sg13g2_decap_8 FILLER_124_720 ();
 sg13g2_decap_8 FILLER_124_727 ();
 sg13g2_decap_8 FILLER_124_734 ();
 sg13g2_decap_8 FILLER_124_741 ();
 sg13g2_decap_4 FILLER_124_748 ();
 sg13g2_fill_2 FILLER_124_764 ();
 sg13g2_decap_8 FILLER_124_778 ();
 sg13g2_decap_8 FILLER_124_785 ();
 sg13g2_decap_8 FILLER_124_792 ();
 sg13g2_decap_8 FILLER_124_799 ();
 sg13g2_fill_2 FILLER_124_806 ();
 sg13g2_decap_8 FILLER_124_835 ();
 sg13g2_decap_8 FILLER_124_842 ();
 sg13g2_decap_8 FILLER_124_849 ();
 sg13g2_fill_1 FILLER_124_856 ();
 sg13g2_decap_8 FILLER_124_881 ();
 sg13g2_decap_8 FILLER_124_888 ();
 sg13g2_decap_8 FILLER_124_895 ();
 sg13g2_decap_8 FILLER_124_902 ();
 sg13g2_decap_4 FILLER_124_909 ();
 sg13g2_decap_8 FILLER_124_917 ();
 sg13g2_fill_1 FILLER_124_924 ();
 sg13g2_decap_8 FILLER_124_942 ();
 sg13g2_decap_8 FILLER_124_949 ();
 sg13g2_decap_8 FILLER_124_956 ();
 sg13g2_decap_8 FILLER_124_963 ();
 sg13g2_decap_4 FILLER_124_970 ();
 sg13g2_decap_8 FILLER_124_982 ();
 sg13g2_fill_2 FILLER_124_989 ();
 sg13g2_decap_8 FILLER_124_995 ();
 sg13g2_decap_8 FILLER_124_1002 ();
 sg13g2_decap_8 FILLER_124_1022 ();
 sg13g2_decap_8 FILLER_124_1029 ();
 sg13g2_decap_8 FILLER_124_1036 ();
 sg13g2_decap_8 FILLER_124_1043 ();
 sg13g2_decap_4 FILLER_124_1050 ();
 sg13g2_fill_1 FILLER_124_1054 ();
 sg13g2_decap_8 FILLER_124_1076 ();
 sg13g2_decap_8 FILLER_124_1083 ();
 sg13g2_decap_8 FILLER_124_1090 ();
 sg13g2_decap_4 FILLER_124_1097 ();
 sg13g2_decap_4 FILLER_124_1118 ();
 sg13g2_fill_1 FILLER_124_1122 ();
 sg13g2_decap_8 FILLER_124_1136 ();
 sg13g2_decap_8 FILLER_124_1143 ();
 sg13g2_decap_4 FILLER_124_1150 ();
 sg13g2_fill_1 FILLER_124_1154 ();
 sg13g2_decap_8 FILLER_124_1186 ();
 sg13g2_fill_2 FILLER_124_1193 ();
 sg13g2_fill_1 FILLER_124_1195 ();
 sg13g2_decap_8 FILLER_124_1204 ();
 sg13g2_decap_8 FILLER_124_1211 ();
 sg13g2_decap_8 FILLER_124_1218 ();
 sg13g2_decap_8 FILLER_124_1225 ();
 sg13g2_decap_8 FILLER_124_1232 ();
 sg13g2_decap_4 FILLER_124_1239 ();
 sg13g2_decap_4 FILLER_124_1267 ();
 sg13g2_decap_8 FILLER_124_1298 ();
 sg13g2_fill_2 FILLER_124_1305 ();
 sg13g2_fill_1 FILLER_124_1307 ();
 sg13g2_decap_4 FILLER_124_1323 ();
 sg13g2_fill_2 FILLER_124_1327 ();
 sg13g2_fill_1 FILLER_124_1334 ();
 sg13g2_decap_8 FILLER_124_1348 ();
 sg13g2_decap_8 FILLER_124_1355 ();
 sg13g2_decap_8 FILLER_124_1362 ();
 sg13g2_fill_1 FILLER_124_1369 ();
 sg13g2_decap_8 FILLER_124_1387 ();
 sg13g2_decap_8 FILLER_124_1394 ();
 sg13g2_decap_8 FILLER_124_1401 ();
 sg13g2_decap_8 FILLER_124_1408 ();
 sg13g2_decap_4 FILLER_124_1415 ();
 sg13g2_fill_2 FILLER_124_1419 ();
 sg13g2_decap_8 FILLER_124_1437 ();
 sg13g2_decap_8 FILLER_124_1444 ();
 sg13g2_decap_8 FILLER_124_1451 ();
 sg13g2_decap_8 FILLER_124_1458 ();
 sg13g2_decap_8 FILLER_124_1465 ();
 sg13g2_decap_8 FILLER_124_1472 ();
 sg13g2_decap_8 FILLER_124_1479 ();
 sg13g2_decap_4 FILLER_124_1486 ();
 sg13g2_fill_2 FILLER_124_1490 ();
 sg13g2_decap_8 FILLER_124_1496 ();
 sg13g2_fill_1 FILLER_124_1503 ();
 sg13g2_decap_4 FILLER_124_1509 ();
 sg13g2_fill_1 FILLER_124_1513 ();
 sg13g2_decap_8 FILLER_124_1517 ();
 sg13g2_decap_8 FILLER_124_1524 ();
 sg13g2_decap_8 FILLER_124_1531 ();
 sg13g2_fill_2 FILLER_124_1538 ();
 sg13g2_fill_1 FILLER_124_1540 ();
 sg13g2_decap_8 FILLER_124_1549 ();
 sg13g2_decap_8 FILLER_124_1556 ();
 sg13g2_decap_8 FILLER_124_1563 ();
 sg13g2_decap_8 FILLER_124_1570 ();
 sg13g2_decap_8 FILLER_124_1577 ();
 sg13g2_decap_8 FILLER_124_1584 ();
 sg13g2_decap_4 FILLER_124_1591 ();
 sg13g2_fill_2 FILLER_124_1595 ();
 sg13g2_fill_1 FILLER_124_1602 ();
 sg13g2_fill_2 FILLER_124_1611 ();
 sg13g2_decap_8 FILLER_124_1625 ();
 sg13g2_decap_8 FILLER_124_1632 ();
 sg13g2_decap_8 FILLER_124_1639 ();
 sg13g2_decap_4 FILLER_124_1646 ();
 sg13g2_fill_1 FILLER_124_1650 ();
 sg13g2_decap_8 FILLER_124_1664 ();
 sg13g2_decap_8 FILLER_124_1671 ();
 sg13g2_fill_2 FILLER_124_1678 ();
 sg13g2_decap_8 FILLER_124_1692 ();
 sg13g2_decap_8 FILLER_124_1699 ();
 sg13g2_decap_8 FILLER_124_1706 ();
 sg13g2_decap_8 FILLER_124_1713 ();
 sg13g2_decap_8 FILLER_124_1720 ();
 sg13g2_decap_4 FILLER_124_1727 ();
 sg13g2_decap_8 FILLER_124_1752 ();
 sg13g2_decap_8 FILLER_124_1759 ();
 sg13g2_fill_2 FILLER_124_1766 ();
 sg13g2_decap_8 FILLER_125_0 ();
 sg13g2_decap_8 FILLER_125_7 ();
 sg13g2_decap_8 FILLER_125_14 ();
 sg13g2_decap_8 FILLER_125_21 ();
 sg13g2_fill_2 FILLER_125_28 ();
 sg13g2_fill_1 FILLER_125_30 ();
 sg13g2_decap_8 FILLER_125_55 ();
 sg13g2_decap_8 FILLER_125_62 ();
 sg13g2_decap_8 FILLER_125_69 ();
 sg13g2_decap_8 FILLER_125_76 ();
 sg13g2_fill_1 FILLER_125_91 ();
 sg13g2_decap_8 FILLER_125_102 ();
 sg13g2_decap_8 FILLER_125_109 ();
 sg13g2_decap_8 FILLER_125_116 ();
 sg13g2_decap_8 FILLER_125_123 ();
 sg13g2_decap_4 FILLER_125_130 ();
 sg13g2_fill_1 FILLER_125_134 ();
 sg13g2_decap_8 FILLER_125_140 ();
 sg13g2_decap_8 FILLER_125_147 ();
 sg13g2_fill_2 FILLER_125_154 ();
 sg13g2_fill_1 FILLER_125_156 ();
 sg13g2_decap_8 FILLER_125_209 ();
 sg13g2_decap_8 FILLER_125_216 ();
 sg13g2_fill_2 FILLER_125_223 ();
 sg13g2_fill_1 FILLER_125_225 ();
 sg13g2_decap_8 FILLER_125_242 ();
 sg13g2_decap_4 FILLER_125_249 ();
 sg13g2_fill_2 FILLER_125_253 ();
 sg13g2_fill_2 FILLER_125_267 ();
 sg13g2_fill_1 FILLER_125_269 ();
 sg13g2_decap_8 FILLER_125_274 ();
 sg13g2_decap_8 FILLER_125_281 ();
 sg13g2_decap_8 FILLER_125_300 ();
 sg13g2_decap_8 FILLER_125_307 ();
 sg13g2_decap_8 FILLER_125_314 ();
 sg13g2_decap_8 FILLER_125_321 ();
 sg13g2_decap_8 FILLER_125_328 ();
 sg13g2_fill_2 FILLER_125_335 ();
 sg13g2_fill_1 FILLER_125_337 ();
 sg13g2_decap_8 FILLER_125_346 ();
 sg13g2_decap_8 FILLER_125_353 ();
 sg13g2_decap_8 FILLER_125_360 ();
 sg13g2_decap_8 FILLER_125_367 ();
 sg13g2_decap_8 FILLER_125_374 ();
 sg13g2_decap_8 FILLER_125_381 ();
 sg13g2_decap_8 FILLER_125_388 ();
 sg13g2_decap_8 FILLER_125_395 ();
 sg13g2_decap_8 FILLER_125_402 ();
 sg13g2_decap_4 FILLER_125_409 ();
 sg13g2_decap_8 FILLER_125_421 ();
 sg13g2_decap_8 FILLER_125_461 ();
 sg13g2_decap_4 FILLER_125_468 ();
 sg13g2_decap_8 FILLER_125_475 ();
 sg13g2_decap_8 FILLER_125_482 ();
 sg13g2_fill_2 FILLER_125_489 ();
 sg13g2_fill_1 FILLER_125_491 ();
 sg13g2_decap_8 FILLER_125_521 ();
 sg13g2_decap_8 FILLER_125_528 ();
 sg13g2_decap_8 FILLER_125_535 ();
 sg13g2_decap_8 FILLER_125_542 ();
 sg13g2_decap_8 FILLER_125_549 ();
 sg13g2_decap_8 FILLER_125_556 ();
 sg13g2_decap_8 FILLER_125_563 ();
 sg13g2_decap_8 FILLER_125_570 ();
 sg13g2_decap_8 FILLER_125_577 ();
 sg13g2_fill_2 FILLER_125_602 ();
 sg13g2_fill_1 FILLER_125_604 ();
 sg13g2_fill_2 FILLER_125_608 ();
 sg13g2_decap_8 FILLER_125_615 ();
 sg13g2_decap_4 FILLER_125_622 ();
 sg13g2_decap_8 FILLER_125_638 ();
 sg13g2_decap_8 FILLER_125_645 ();
 sg13g2_decap_8 FILLER_125_652 ();
 sg13g2_decap_8 FILLER_125_659 ();
 sg13g2_decap_8 FILLER_125_666 ();
 sg13g2_decap_4 FILLER_125_673 ();
 sg13g2_fill_1 FILLER_125_677 ();
 sg13g2_decap_8 FILLER_125_714 ();
 sg13g2_decap_8 FILLER_125_721 ();
 sg13g2_decap_8 FILLER_125_728 ();
 sg13g2_decap_8 FILLER_125_735 ();
 sg13g2_fill_2 FILLER_125_742 ();
 sg13g2_fill_1 FILLER_125_744 ();
 sg13g2_decap_8 FILLER_125_753 ();
 sg13g2_fill_2 FILLER_125_760 ();
 sg13g2_decap_8 FILLER_125_770 ();
 sg13g2_decap_8 FILLER_125_777 ();
 sg13g2_decap_8 FILLER_125_784 ();
 sg13g2_decap_8 FILLER_125_791 ();
 sg13g2_decap_8 FILLER_125_798 ();
 sg13g2_decap_8 FILLER_125_805 ();
 sg13g2_fill_1 FILLER_125_829 ();
 sg13g2_decap_8 FILLER_125_835 ();
 sg13g2_decap_8 FILLER_125_842 ();
 sg13g2_decap_8 FILLER_125_849 ();
 sg13g2_decap_4 FILLER_125_856 ();
 sg13g2_decap_8 FILLER_125_863 ();
 sg13g2_decap_8 FILLER_125_870 ();
 sg13g2_decap_8 FILLER_125_877 ();
 sg13g2_decap_8 FILLER_125_884 ();
 sg13g2_decap_8 FILLER_125_891 ();
 sg13g2_decap_8 FILLER_125_898 ();
 sg13g2_decap_8 FILLER_125_905 ();
 sg13g2_decap_8 FILLER_125_912 ();
 sg13g2_decap_8 FILLER_125_919 ();
 sg13g2_fill_2 FILLER_125_926 ();
 sg13g2_fill_2 FILLER_125_937 ();
 sg13g2_fill_1 FILLER_125_939 ();
 sg13g2_decap_8 FILLER_125_944 ();
 sg13g2_decap_8 FILLER_125_951 ();
 sg13g2_decap_8 FILLER_125_958 ();
 sg13g2_decap_8 FILLER_125_965 ();
 sg13g2_decap_8 FILLER_125_972 ();
 sg13g2_decap_8 FILLER_125_979 ();
 sg13g2_fill_2 FILLER_125_986 ();
 sg13g2_fill_1 FILLER_125_988 ();
 sg13g2_decap_8 FILLER_125_997 ();
 sg13g2_decap_8 FILLER_125_1004 ();
 sg13g2_decap_8 FILLER_125_1011 ();
 sg13g2_decap_8 FILLER_125_1018 ();
 sg13g2_decap_8 FILLER_125_1025 ();
 sg13g2_decap_8 FILLER_125_1036 ();
 sg13g2_decap_8 FILLER_125_1043 ();
 sg13g2_decap_8 FILLER_125_1050 ();
 sg13g2_fill_2 FILLER_125_1057 ();
 sg13g2_decap_4 FILLER_125_1064 ();
 sg13g2_decap_8 FILLER_125_1081 ();
 sg13g2_decap_8 FILLER_125_1088 ();
 sg13g2_decap_4 FILLER_125_1095 ();
 sg13g2_fill_2 FILLER_125_1099 ();
 sg13g2_decap_8 FILLER_125_1144 ();
 sg13g2_decap_8 FILLER_125_1159 ();
 sg13g2_fill_2 FILLER_125_1166 ();
 sg13g2_fill_1 FILLER_125_1168 ();
 sg13g2_decap_8 FILLER_125_1173 ();
 sg13g2_decap_8 FILLER_125_1180 ();
 sg13g2_decap_8 FILLER_125_1187 ();
 sg13g2_decap_8 FILLER_125_1194 ();
 sg13g2_decap_8 FILLER_125_1201 ();
 sg13g2_decap_8 FILLER_125_1208 ();
 sg13g2_decap_8 FILLER_125_1215 ();
 sg13g2_decap_8 FILLER_125_1222 ();
 sg13g2_decap_8 FILLER_125_1229 ();
 sg13g2_decap_8 FILLER_125_1236 ();
 sg13g2_decap_8 FILLER_125_1243 ();
 sg13g2_decap_8 FILLER_125_1250 ();
 sg13g2_decap_8 FILLER_125_1261 ();
 sg13g2_decap_8 FILLER_125_1268 ();
 sg13g2_fill_2 FILLER_125_1275 ();
 sg13g2_fill_2 FILLER_125_1281 ();
 sg13g2_fill_1 FILLER_125_1283 ();
 sg13g2_decap_8 FILLER_125_1296 ();
 sg13g2_decap_8 FILLER_125_1303 ();
 sg13g2_decap_8 FILLER_125_1310 ();
 sg13g2_fill_2 FILLER_125_1317 ();
 sg13g2_decap_4 FILLER_125_1338 ();
 sg13g2_fill_2 FILLER_125_1354 ();
 sg13g2_fill_2 FILLER_125_1359 ();
 sg13g2_fill_1 FILLER_125_1361 ();
 sg13g2_decap_8 FILLER_125_1366 ();
 sg13g2_decap_8 FILLER_125_1373 ();
 sg13g2_decap_8 FILLER_125_1380 ();
 sg13g2_decap_8 FILLER_125_1387 ();
 sg13g2_decap_8 FILLER_125_1394 ();
 sg13g2_decap_8 FILLER_125_1401 ();
 sg13g2_decap_8 FILLER_125_1408 ();
 sg13g2_decap_8 FILLER_125_1415 ();
 sg13g2_decap_8 FILLER_125_1422 ();
 sg13g2_decap_8 FILLER_125_1429 ();
 sg13g2_decap_8 FILLER_125_1436 ();
 sg13g2_decap_8 FILLER_125_1443 ();
 sg13g2_decap_8 FILLER_125_1450 ();
 sg13g2_decap_8 FILLER_125_1457 ();
 sg13g2_decap_4 FILLER_125_1464 ();
 sg13g2_decap_8 FILLER_125_1484 ();
 sg13g2_decap_8 FILLER_125_1491 ();
 sg13g2_fill_2 FILLER_125_1498 ();
 sg13g2_fill_1 FILLER_125_1500 ();
 sg13g2_fill_1 FILLER_125_1514 ();
 sg13g2_decap_8 FILLER_125_1527 ();
 sg13g2_decap_8 FILLER_125_1534 ();
 sg13g2_decap_4 FILLER_125_1546 ();
 sg13g2_fill_2 FILLER_125_1550 ();
 sg13g2_fill_2 FILLER_125_1573 ();
 sg13g2_fill_1 FILLER_125_1575 ();
 sg13g2_decap_8 FILLER_125_1614 ();
 sg13g2_decap_8 FILLER_125_1621 ();
 sg13g2_decap_8 FILLER_125_1628 ();
 sg13g2_decap_8 FILLER_125_1635 ();
 sg13g2_decap_8 FILLER_125_1642 ();
 sg13g2_decap_4 FILLER_125_1649 ();
 sg13g2_fill_2 FILLER_125_1653 ();
 sg13g2_fill_2 FILLER_125_1660 ();
 sg13g2_fill_1 FILLER_125_1662 ();
 sg13g2_fill_2 FILLER_125_1668 ();
 sg13g2_decap_8 FILLER_125_1673 ();
 sg13g2_decap_8 FILLER_125_1680 ();
 sg13g2_decap_8 FILLER_125_1687 ();
 sg13g2_decap_8 FILLER_125_1694 ();
 sg13g2_decap_8 FILLER_125_1701 ();
 sg13g2_decap_8 FILLER_125_1708 ();
 sg13g2_decap_8 FILLER_125_1715 ();
 sg13g2_fill_2 FILLER_125_1722 ();
 sg13g2_fill_1 FILLER_125_1724 ();
 sg13g2_decap_8 FILLER_125_1734 ();
 sg13g2_decap_4 FILLER_125_1741 ();
 sg13g2_fill_1 FILLER_125_1745 ();
 sg13g2_decap_8 FILLER_125_1750 ();
 sg13g2_decap_8 FILLER_125_1757 ();
 sg13g2_decap_4 FILLER_125_1764 ();
 sg13g2_decap_8 FILLER_126_0 ();
 sg13g2_decap_8 FILLER_126_7 ();
 sg13g2_decap_8 FILLER_126_14 ();
 sg13g2_decap_8 FILLER_126_21 ();
 sg13g2_decap_8 FILLER_126_28 ();
 sg13g2_decap_8 FILLER_126_35 ();
 sg13g2_fill_2 FILLER_126_42 ();
 sg13g2_decap_4 FILLER_126_52 ();
 sg13g2_decap_8 FILLER_126_65 ();
 sg13g2_decap_8 FILLER_126_72 ();
 sg13g2_decap_8 FILLER_126_79 ();
 sg13g2_decap_8 FILLER_126_86 ();
 sg13g2_decap_8 FILLER_126_93 ();
 sg13g2_decap_8 FILLER_126_100 ();
 sg13g2_decap_8 FILLER_126_107 ();
 sg13g2_decap_8 FILLER_126_114 ();
 sg13g2_decap_4 FILLER_126_121 ();
 sg13g2_fill_2 FILLER_126_125 ();
 sg13g2_decap_8 FILLER_126_137 ();
 sg13g2_decap_8 FILLER_126_144 ();
 sg13g2_decap_8 FILLER_126_151 ();
 sg13g2_decap_8 FILLER_126_158 ();
 sg13g2_decap_8 FILLER_126_165 ();
 sg13g2_decap_8 FILLER_126_172 ();
 sg13g2_decap_8 FILLER_126_179 ();
 sg13g2_decap_8 FILLER_126_186 ();
 sg13g2_fill_2 FILLER_126_193 ();
 sg13g2_fill_1 FILLER_126_195 ();
 sg13g2_decap_8 FILLER_126_214 ();
 sg13g2_decap_8 FILLER_126_221 ();
 sg13g2_decap_8 FILLER_126_228 ();
 sg13g2_decap_8 FILLER_126_235 ();
 sg13g2_decap_8 FILLER_126_242 ();
 sg13g2_decap_8 FILLER_126_249 ();
 sg13g2_decap_8 FILLER_126_256 ();
 sg13g2_decap_8 FILLER_126_263 ();
 sg13g2_decap_8 FILLER_126_270 ();
 sg13g2_decap_4 FILLER_126_277 ();
 sg13g2_fill_1 FILLER_126_281 ();
 sg13g2_decap_8 FILLER_126_306 ();
 sg13g2_decap_8 FILLER_126_313 ();
 sg13g2_decap_8 FILLER_126_320 ();
 sg13g2_decap_8 FILLER_126_327 ();
 sg13g2_decap_4 FILLER_126_334 ();
 sg13g2_fill_2 FILLER_126_338 ();
 sg13g2_decap_8 FILLER_126_346 ();
 sg13g2_decap_8 FILLER_126_353 ();
 sg13g2_decap_4 FILLER_126_360 ();
 sg13g2_fill_2 FILLER_126_364 ();
 sg13g2_decap_8 FILLER_126_374 ();
 sg13g2_decap_8 FILLER_126_381 ();
 sg13g2_decap_8 FILLER_126_388 ();
 sg13g2_decap_8 FILLER_126_395 ();
 sg13g2_decap_8 FILLER_126_402 ();
 sg13g2_decap_8 FILLER_126_409 ();
 sg13g2_decap_8 FILLER_126_416 ();
 sg13g2_decap_8 FILLER_126_423 ();
 sg13g2_fill_2 FILLER_126_430 ();
 sg13g2_decap_4 FILLER_126_436 ();
 sg13g2_fill_1 FILLER_126_440 ();
 sg13g2_decap_4 FILLER_126_454 ();
 sg13g2_fill_1 FILLER_126_458 ();
 sg13g2_decap_8 FILLER_126_462 ();
 sg13g2_decap_8 FILLER_126_481 ();
 sg13g2_decap_8 FILLER_126_488 ();
 sg13g2_fill_2 FILLER_126_495 ();
 sg13g2_decap_8 FILLER_126_514 ();
 sg13g2_decap_8 FILLER_126_521 ();
 sg13g2_fill_2 FILLER_126_548 ();
 sg13g2_fill_1 FILLER_126_550 ();
 sg13g2_decap_8 FILLER_126_557 ();
 sg13g2_decap_8 FILLER_126_564 ();
 sg13g2_decap_8 FILLER_126_571 ();
 sg13g2_decap_8 FILLER_126_578 ();
 sg13g2_fill_2 FILLER_126_585 ();
 sg13g2_decap_8 FILLER_126_601 ();
 sg13g2_decap_4 FILLER_126_608 ();
 sg13g2_decap_8 FILLER_126_625 ();
 sg13g2_decap_8 FILLER_126_632 ();
 sg13g2_decap_8 FILLER_126_639 ();
 sg13g2_decap_8 FILLER_126_646 ();
 sg13g2_decap_8 FILLER_126_653 ();
 sg13g2_decap_8 FILLER_126_660 ();
 sg13g2_fill_2 FILLER_126_667 ();
 sg13g2_decap_8 FILLER_126_693 ();
 sg13g2_fill_2 FILLER_126_700 ();
 sg13g2_fill_1 FILLER_126_702 ();
 sg13g2_fill_2 FILLER_126_707 ();
 sg13g2_decap_8 FILLER_126_721 ();
 sg13g2_decap_8 FILLER_126_728 ();
 sg13g2_decap_8 FILLER_126_735 ();
 sg13g2_decap_8 FILLER_126_742 ();
 sg13g2_decap_8 FILLER_126_749 ();
 sg13g2_decap_8 FILLER_126_756 ();
 sg13g2_decap_8 FILLER_126_763 ();
 sg13g2_decap_8 FILLER_126_770 ();
 sg13g2_decap_8 FILLER_126_777 ();
 sg13g2_decap_8 FILLER_126_784 ();
 sg13g2_decap_8 FILLER_126_791 ();
 sg13g2_decap_8 FILLER_126_798 ();
 sg13g2_decap_8 FILLER_126_805 ();
 sg13g2_decap_8 FILLER_126_820 ();
 sg13g2_decap_8 FILLER_126_827 ();
 sg13g2_decap_8 FILLER_126_834 ();
 sg13g2_decap_8 FILLER_126_841 ();
 sg13g2_decap_8 FILLER_126_848 ();
 sg13g2_decap_4 FILLER_126_855 ();
 sg13g2_fill_2 FILLER_126_859 ();
 sg13g2_fill_2 FILLER_126_869 ();
 sg13g2_fill_1 FILLER_126_871 ();
 sg13g2_decap_8 FILLER_126_877 ();
 sg13g2_fill_2 FILLER_126_884 ();
 sg13g2_fill_1 FILLER_126_886 ();
 sg13g2_decap_8 FILLER_126_897 ();
 sg13g2_decap_8 FILLER_126_904 ();
 sg13g2_decap_8 FILLER_126_911 ();
 sg13g2_decap_8 FILLER_126_918 ();
 sg13g2_fill_2 FILLER_126_925 ();
 sg13g2_fill_2 FILLER_126_971 ();
 sg13g2_decap_8 FILLER_126_986 ();
 sg13g2_decap_8 FILLER_126_993 ();
 sg13g2_decap_8 FILLER_126_1000 ();
 sg13g2_decap_8 FILLER_126_1012 ();
 sg13g2_decap_8 FILLER_126_1019 ();
 sg13g2_fill_2 FILLER_126_1026 ();
 sg13g2_decap_8 FILLER_126_1045 ();
 sg13g2_decap_8 FILLER_126_1052 ();
 sg13g2_decap_8 FILLER_126_1059 ();
 sg13g2_decap_8 FILLER_126_1066 ();
 sg13g2_decap_8 FILLER_126_1073 ();
 sg13g2_decap_8 FILLER_126_1080 ();
 sg13g2_decap_8 FILLER_126_1087 ();
 sg13g2_decap_8 FILLER_126_1094 ();
 sg13g2_decap_8 FILLER_126_1101 ();
 sg13g2_decap_4 FILLER_126_1108 ();
 sg13g2_decap_8 FILLER_126_1116 ();
 sg13g2_decap_4 FILLER_126_1123 ();
 sg13g2_decap_8 FILLER_126_1136 ();
 sg13g2_decap_8 FILLER_126_1143 ();
 sg13g2_decap_4 FILLER_126_1150 ();
 sg13g2_fill_1 FILLER_126_1160 ();
 sg13g2_decap_8 FILLER_126_1174 ();
 sg13g2_fill_2 FILLER_126_1181 ();
 sg13g2_decap_8 FILLER_126_1199 ();
 sg13g2_fill_2 FILLER_126_1206 ();
 sg13g2_decap_8 FILLER_126_1212 ();
 sg13g2_decap_8 FILLER_126_1227 ();
 sg13g2_decap_8 FILLER_126_1239 ();
 sg13g2_decap_4 FILLER_126_1246 ();
 sg13g2_decap_8 FILLER_126_1269 ();
 sg13g2_fill_1 FILLER_126_1276 ();
 sg13g2_fill_2 FILLER_126_1285 ();
 sg13g2_decap_8 FILLER_126_1306 ();
 sg13g2_decap_4 FILLER_126_1313 ();
 sg13g2_fill_2 FILLER_126_1317 ();
 sg13g2_decap_8 FILLER_126_1336 ();
 sg13g2_decap_8 FILLER_126_1343 ();
 sg13g2_decap_8 FILLER_126_1350 ();
 sg13g2_decap_8 FILLER_126_1357 ();
 sg13g2_fill_2 FILLER_126_1364 ();
 sg13g2_fill_2 FILLER_126_1371 ();
 sg13g2_decap_8 FILLER_126_1381 ();
 sg13g2_decap_8 FILLER_126_1388 ();
 sg13g2_decap_8 FILLER_126_1395 ();
 sg13g2_decap_8 FILLER_126_1402 ();
 sg13g2_decap_8 FILLER_126_1409 ();
 sg13g2_decap_8 FILLER_126_1416 ();
 sg13g2_decap_8 FILLER_126_1423 ();
 sg13g2_decap_8 FILLER_126_1430 ();
 sg13g2_fill_1 FILLER_126_1437 ();
 sg13g2_decap_8 FILLER_126_1448 ();
 sg13g2_decap_8 FILLER_126_1455 ();
 sg13g2_decap_8 FILLER_126_1462 ();
 sg13g2_decap_8 FILLER_126_1469 ();
 sg13g2_decap_8 FILLER_126_1476 ();
 sg13g2_fill_2 FILLER_126_1483 ();
 sg13g2_fill_1 FILLER_126_1485 ();
 sg13g2_fill_2 FILLER_126_1492 ();
 sg13g2_fill_1 FILLER_126_1494 ();
 sg13g2_decap_8 FILLER_126_1500 ();
 sg13g2_fill_1 FILLER_126_1507 ();
 sg13g2_decap_8 FILLER_126_1534 ();
 sg13g2_decap_8 FILLER_126_1541 ();
 sg13g2_decap_8 FILLER_126_1548 ();
 sg13g2_decap_4 FILLER_126_1555 ();
 sg13g2_fill_2 FILLER_126_1563 ();
 sg13g2_decap_8 FILLER_126_1571 ();
 sg13g2_decap_8 FILLER_126_1578 ();
 sg13g2_decap_4 FILLER_126_1590 ();
 sg13g2_decap_8 FILLER_126_1611 ();
 sg13g2_decap_8 FILLER_126_1618 ();
 sg13g2_decap_8 FILLER_126_1625 ();
 sg13g2_decap_8 FILLER_126_1632 ();
 sg13g2_decap_8 FILLER_126_1639 ();
 sg13g2_decap_8 FILLER_126_1646 ();
 sg13g2_decap_8 FILLER_126_1653 ();
 sg13g2_decap_4 FILLER_126_1660 ();
 sg13g2_fill_2 FILLER_126_1664 ();
 sg13g2_decap_8 FILLER_126_1674 ();
 sg13g2_decap_4 FILLER_126_1681 ();
 sg13g2_fill_1 FILLER_126_1685 ();
 sg13g2_fill_1 FILLER_126_1690 ();
 sg13g2_decap_8 FILLER_126_1695 ();
 sg13g2_decap_8 FILLER_126_1702 ();
 sg13g2_decap_4 FILLER_126_1709 ();
 sg13g2_fill_1 FILLER_126_1713 ();
 sg13g2_decap_8 FILLER_126_1741 ();
 sg13g2_decap_8 FILLER_126_1748 ();
 sg13g2_decap_8 FILLER_126_1755 ();
 sg13g2_decap_4 FILLER_126_1762 ();
 sg13g2_fill_2 FILLER_126_1766 ();
 sg13g2_decap_8 FILLER_127_0 ();
 sg13g2_decap_8 FILLER_127_7 ();
 sg13g2_decap_8 FILLER_127_14 ();
 sg13g2_decap_8 FILLER_127_21 ();
 sg13g2_decap_8 FILLER_127_28 ();
 sg13g2_fill_2 FILLER_127_35 ();
 sg13g2_fill_2 FILLER_127_45 ();
 sg13g2_decap_8 FILLER_127_52 ();
 sg13g2_decap_8 FILLER_127_59 ();
 sg13g2_decap_8 FILLER_127_66 ();
 sg13g2_decap_8 FILLER_127_73 ();
 sg13g2_fill_2 FILLER_127_80 ();
 sg13g2_fill_1 FILLER_127_82 ();
 sg13g2_decap_8 FILLER_127_88 ();
 sg13g2_decap_8 FILLER_127_95 ();
 sg13g2_decap_8 FILLER_127_102 ();
 sg13g2_decap_8 FILLER_127_109 ();
 sg13g2_decap_8 FILLER_127_116 ();
 sg13g2_fill_1 FILLER_127_123 ();
 sg13g2_decap_8 FILLER_127_141 ();
 sg13g2_decap_8 FILLER_127_148 ();
 sg13g2_decap_4 FILLER_127_155 ();
 sg13g2_decap_8 FILLER_127_162 ();
 sg13g2_decap_8 FILLER_127_169 ();
 sg13g2_decap_8 FILLER_127_176 ();
 sg13g2_fill_2 FILLER_127_183 ();
 sg13g2_decap_8 FILLER_127_191 ();
 sg13g2_decap_8 FILLER_127_198 ();
 sg13g2_decap_8 FILLER_127_205 ();
 sg13g2_decap_8 FILLER_127_212 ();
 sg13g2_decap_8 FILLER_127_219 ();
 sg13g2_decap_8 FILLER_127_226 ();
 sg13g2_decap_8 FILLER_127_233 ();
 sg13g2_decap_4 FILLER_127_240 ();
 sg13g2_fill_1 FILLER_127_244 ();
 sg13g2_decap_8 FILLER_127_253 ();
 sg13g2_decap_8 FILLER_127_260 ();
 sg13g2_decap_8 FILLER_127_267 ();
 sg13g2_decap_8 FILLER_127_274 ();
 sg13g2_fill_2 FILLER_127_281 ();
 sg13g2_decap_4 FILLER_127_291 ();
 sg13g2_decap_8 FILLER_127_305 ();
 sg13g2_decap_8 FILLER_127_312 ();
 sg13g2_decap_8 FILLER_127_319 ();
 sg13g2_fill_1 FILLER_127_326 ();
 sg13g2_decap_4 FILLER_127_331 ();
 sg13g2_decap_8 FILLER_127_352 ();
 sg13g2_decap_8 FILLER_127_359 ();
 sg13g2_decap_4 FILLER_127_366 ();
 sg13g2_fill_2 FILLER_127_370 ();
 sg13g2_decap_8 FILLER_127_386 ();
 sg13g2_fill_1 FILLER_127_393 ();
 sg13g2_decap_8 FILLER_127_397 ();
 sg13g2_decap_8 FILLER_127_404 ();
 sg13g2_decap_8 FILLER_127_411 ();
 sg13g2_decap_8 FILLER_127_418 ();
 sg13g2_decap_8 FILLER_127_425 ();
 sg13g2_decap_8 FILLER_127_432 ();
 sg13g2_decap_8 FILLER_127_439 ();
 sg13g2_decap_8 FILLER_127_446 ();
 sg13g2_fill_2 FILLER_127_453 ();
 sg13g2_fill_1 FILLER_127_455 ();
 sg13g2_decap_4 FILLER_127_467 ();
 sg13g2_fill_1 FILLER_127_471 ();
 sg13g2_fill_1 FILLER_127_475 ();
 sg13g2_decap_8 FILLER_127_480 ();
 sg13g2_decap_8 FILLER_127_487 ();
 sg13g2_decap_8 FILLER_127_494 ();
 sg13g2_decap_8 FILLER_127_501 ();
 sg13g2_decap_8 FILLER_127_508 ();
 sg13g2_decap_8 FILLER_127_515 ();
 sg13g2_decap_4 FILLER_127_522 ();
 sg13g2_fill_1 FILLER_127_526 ();
 sg13g2_decap_8 FILLER_127_568 ();
 sg13g2_decap_4 FILLER_127_575 ();
 sg13g2_fill_1 FILLER_127_579 ();
 sg13g2_decap_8 FILLER_127_583 ();
 sg13g2_decap_8 FILLER_127_616 ();
 sg13g2_decap_8 FILLER_127_623 ();
 sg13g2_decap_8 FILLER_127_630 ();
 sg13g2_decap_8 FILLER_127_637 ();
 sg13g2_decap_8 FILLER_127_644 ();
 sg13g2_decap_8 FILLER_127_651 ();
 sg13g2_decap_8 FILLER_127_658 ();
 sg13g2_decap_8 FILLER_127_665 ();
 sg13g2_decap_4 FILLER_127_672 ();
 sg13g2_fill_1 FILLER_127_681 ();
 sg13g2_decap_8 FILLER_127_690 ();
 sg13g2_decap_8 FILLER_127_697 ();
 sg13g2_decap_8 FILLER_127_704 ();
 sg13g2_decap_8 FILLER_127_711 ();
 sg13g2_decap_4 FILLER_127_718 ();
 sg13g2_fill_1 FILLER_127_722 ();
 sg13g2_fill_1 FILLER_127_727 ();
 sg13g2_decap_8 FILLER_127_732 ();
 sg13g2_decap_8 FILLER_127_739 ();
 sg13g2_decap_8 FILLER_127_746 ();
 sg13g2_fill_2 FILLER_127_753 ();
 sg13g2_decap_4 FILLER_127_765 ();
 sg13g2_decap_8 FILLER_127_782 ();
 sg13g2_fill_2 FILLER_127_789 ();
 sg13g2_decap_8 FILLER_127_800 ();
 sg13g2_decap_8 FILLER_127_807 ();
 sg13g2_fill_2 FILLER_127_814 ();
 sg13g2_fill_1 FILLER_127_816 ();
 sg13g2_decap_8 FILLER_127_830 ();
 sg13g2_decap_8 FILLER_127_837 ();
 sg13g2_decap_4 FILLER_127_844 ();
 sg13g2_fill_2 FILLER_127_848 ();
 sg13g2_fill_1 FILLER_127_855 ();
 sg13g2_fill_2 FILLER_127_863 ();
 sg13g2_decap_8 FILLER_127_880 ();
 sg13g2_decap_8 FILLER_127_887 ();
 sg13g2_decap_8 FILLER_127_894 ();
 sg13g2_decap_8 FILLER_127_901 ();
 sg13g2_fill_1 FILLER_127_908 ();
 sg13g2_decap_8 FILLER_127_919 ();
 sg13g2_decap_8 FILLER_127_926 ();
 sg13g2_decap_8 FILLER_127_933 ();
 sg13g2_fill_2 FILLER_127_940 ();
 sg13g2_fill_1 FILLER_127_942 ();
 sg13g2_decap_8 FILLER_127_947 ();
 sg13g2_decap_8 FILLER_127_954 ();
 sg13g2_decap_8 FILLER_127_961 ();
 sg13g2_decap_8 FILLER_127_968 ();
 sg13g2_decap_8 FILLER_127_975 ();
 sg13g2_fill_1 FILLER_127_982 ();
 sg13g2_decap_8 FILLER_127_1003 ();
 sg13g2_decap_8 FILLER_127_1010 ();
 sg13g2_decap_8 FILLER_127_1017 ();
 sg13g2_decap_8 FILLER_127_1024 ();
 sg13g2_fill_2 FILLER_127_1031 ();
 sg13g2_fill_2 FILLER_127_1038 ();
 sg13g2_fill_1 FILLER_127_1040 ();
 sg13g2_decap_8 FILLER_127_1054 ();
 sg13g2_decap_8 FILLER_127_1061 ();
 sg13g2_decap_8 FILLER_127_1068 ();
 sg13g2_decap_8 FILLER_127_1075 ();
 sg13g2_decap_8 FILLER_127_1082 ();
 sg13g2_fill_2 FILLER_127_1089 ();
 sg13g2_decap_8 FILLER_127_1095 ();
 sg13g2_decap_8 FILLER_127_1102 ();
 sg13g2_fill_2 FILLER_127_1109 ();
 sg13g2_decap_8 FILLER_127_1117 ();
 sg13g2_decap_8 FILLER_127_1124 ();
 sg13g2_decap_8 FILLER_127_1131 ();
 sg13g2_decap_8 FILLER_127_1138 ();
 sg13g2_decap_8 FILLER_127_1145 ();
 sg13g2_decap_4 FILLER_127_1152 ();
 sg13g2_fill_2 FILLER_127_1156 ();
 sg13g2_decap_8 FILLER_127_1163 ();
 sg13g2_decap_8 FILLER_127_1170 ();
 sg13g2_decap_8 FILLER_127_1177 ();
 sg13g2_decap_8 FILLER_127_1184 ();
 sg13g2_fill_2 FILLER_127_1194 ();
 sg13g2_fill_2 FILLER_127_1211 ();
 sg13g2_decap_8 FILLER_127_1226 ();
 sg13g2_decap_8 FILLER_127_1233 ();
 sg13g2_decap_8 FILLER_127_1240 ();
 sg13g2_decap_8 FILLER_127_1247 ();
 sg13g2_decap_8 FILLER_127_1254 ();
 sg13g2_decap_8 FILLER_127_1261 ();
 sg13g2_decap_8 FILLER_127_1268 ();
 sg13g2_decap_8 FILLER_127_1275 ();
 sg13g2_fill_2 FILLER_127_1282 ();
 sg13g2_decap_8 FILLER_127_1296 ();
 sg13g2_decap_8 FILLER_127_1303 ();
 sg13g2_decap_8 FILLER_127_1310 ();
 sg13g2_decap_8 FILLER_127_1317 ();
 sg13g2_decap_8 FILLER_127_1324 ();
 sg13g2_decap_8 FILLER_127_1331 ();
 sg13g2_decap_8 FILLER_127_1338 ();
 sg13g2_decap_4 FILLER_127_1345 ();
 sg13g2_fill_2 FILLER_127_1349 ();
 sg13g2_fill_2 FILLER_127_1358 ();
 sg13g2_decap_8 FILLER_127_1372 ();
 sg13g2_decap_8 FILLER_127_1379 ();
 sg13g2_decap_8 FILLER_127_1386 ();
 sg13g2_decap_8 FILLER_127_1393 ();
 sg13g2_decap_4 FILLER_127_1400 ();
 sg13g2_fill_1 FILLER_127_1404 ();
 sg13g2_decap_8 FILLER_127_1410 ();
 sg13g2_decap_4 FILLER_127_1417 ();
 sg13g2_fill_2 FILLER_127_1421 ();
 sg13g2_fill_2 FILLER_127_1427 ();
 sg13g2_fill_2 FILLER_127_1437 ();
 sg13g2_fill_1 FILLER_127_1439 ();
 sg13g2_decap_8 FILLER_127_1453 ();
 sg13g2_decap_8 FILLER_127_1464 ();
 sg13g2_decap_8 FILLER_127_1471 ();
 sg13g2_decap_8 FILLER_127_1478 ();
 sg13g2_fill_2 FILLER_127_1485 ();
 sg13g2_fill_1 FILLER_127_1487 ();
 sg13g2_decap_8 FILLER_127_1491 ();
 sg13g2_decap_8 FILLER_127_1498 ();
 sg13g2_decap_8 FILLER_127_1505 ();
 sg13g2_decap_8 FILLER_127_1512 ();
 sg13g2_decap_4 FILLER_127_1519 ();
 sg13g2_fill_2 FILLER_127_1528 ();
 sg13g2_fill_1 FILLER_127_1530 ();
 sg13g2_fill_1 FILLER_127_1541 ();
 sg13g2_decap_8 FILLER_127_1550 ();
 sg13g2_decap_8 FILLER_127_1557 ();
 sg13g2_decap_8 FILLER_127_1564 ();
 sg13g2_decap_8 FILLER_127_1571 ();
 sg13g2_decap_8 FILLER_127_1578 ();
 sg13g2_fill_2 FILLER_127_1585 ();
 sg13g2_fill_1 FILLER_127_1587 ();
 sg13g2_decap_8 FILLER_127_1599 ();
 sg13g2_decap_8 FILLER_127_1606 ();
 sg13g2_fill_2 FILLER_127_1613 ();
 sg13g2_fill_1 FILLER_127_1615 ();
 sg13g2_fill_1 FILLER_127_1621 ();
 sg13g2_decap_8 FILLER_127_1627 ();
 sg13g2_decap_8 FILLER_127_1634 ();
 sg13g2_decap_8 FILLER_127_1641 ();
 sg13g2_decap_8 FILLER_127_1648 ();
 sg13g2_fill_2 FILLER_127_1655 ();
 sg13g2_decap_8 FILLER_127_1675 ();
 sg13g2_decap_8 FILLER_127_1682 ();
 sg13g2_decap_4 FILLER_127_1689 ();
 sg13g2_fill_2 FILLER_127_1693 ();
 sg13g2_fill_2 FILLER_127_1709 ();
 sg13g2_decap_8 FILLER_127_1740 ();
 sg13g2_decap_8 FILLER_127_1747 ();
 sg13g2_decap_8 FILLER_127_1754 ();
 sg13g2_decap_8 FILLER_127_1761 ();
 sg13g2_decap_8 FILLER_128_0 ();
 sg13g2_decap_8 FILLER_128_7 ();
 sg13g2_decap_4 FILLER_128_14 ();
 sg13g2_fill_2 FILLER_128_34 ();
 sg13g2_fill_1 FILLER_128_40 ();
 sg13g2_decap_8 FILLER_128_45 ();
 sg13g2_decap_8 FILLER_128_52 ();
 sg13g2_decap_8 FILLER_128_59 ();
 sg13g2_decap_8 FILLER_128_66 ();
 sg13g2_decap_4 FILLER_128_73 ();
 sg13g2_fill_2 FILLER_128_93 ();
 sg13g2_fill_1 FILLER_128_95 ();
 sg13g2_decap_8 FILLER_128_99 ();
 sg13g2_decap_4 FILLER_128_106 ();
 sg13g2_fill_1 FILLER_128_110 ();
 sg13g2_decap_8 FILLER_128_137 ();
 sg13g2_decap_8 FILLER_128_144 ();
 sg13g2_decap_4 FILLER_128_151 ();
 sg13g2_fill_1 FILLER_128_155 ();
 sg13g2_fill_1 FILLER_128_167 ();
 sg13g2_decap_8 FILLER_128_172 ();
 sg13g2_decap_8 FILLER_128_179 ();
 sg13g2_decap_8 FILLER_128_186 ();
 sg13g2_decap_8 FILLER_128_193 ();
 sg13g2_decap_8 FILLER_128_200 ();
 sg13g2_fill_1 FILLER_128_207 ();
 sg13g2_fill_2 FILLER_128_216 ();
 sg13g2_fill_1 FILLER_128_218 ();
 sg13g2_decap_8 FILLER_128_225 ();
 sg13g2_decap_4 FILLER_128_232 ();
 sg13g2_fill_1 FILLER_128_248 ();
 sg13g2_decap_8 FILLER_128_253 ();
 sg13g2_decap_8 FILLER_128_260 ();
 sg13g2_decap_8 FILLER_128_267 ();
 sg13g2_decap_8 FILLER_128_274 ();
 sg13g2_decap_8 FILLER_128_281 ();
 sg13g2_decap_8 FILLER_128_288 ();
 sg13g2_decap_8 FILLER_128_295 ();
 sg13g2_decap_8 FILLER_128_302 ();
 sg13g2_decap_8 FILLER_128_309 ();
 sg13g2_decap_8 FILLER_128_316 ();
 sg13g2_fill_2 FILLER_128_323 ();
 sg13g2_fill_1 FILLER_128_325 ();
 sg13g2_decap_8 FILLER_128_339 ();
 sg13g2_decap_8 FILLER_128_346 ();
 sg13g2_decap_8 FILLER_128_353 ();
 sg13g2_decap_8 FILLER_128_360 ();
 sg13g2_decap_8 FILLER_128_371 ();
 sg13g2_decap_8 FILLER_128_378 ();
 sg13g2_fill_2 FILLER_128_385 ();
 sg13g2_fill_1 FILLER_128_387 ();
 sg13g2_decap_8 FILLER_128_399 ();
 sg13g2_decap_8 FILLER_128_406 ();
 sg13g2_decap_8 FILLER_128_413 ();
 sg13g2_decap_8 FILLER_128_420 ();
 sg13g2_decap_8 FILLER_128_427 ();
 sg13g2_decap_8 FILLER_128_434 ();
 sg13g2_decap_8 FILLER_128_441 ();
 sg13g2_decap_8 FILLER_128_448 ();
 sg13g2_decap_4 FILLER_128_467 ();
 sg13g2_fill_2 FILLER_128_471 ();
 sg13g2_decap_8 FILLER_128_480 ();
 sg13g2_decap_8 FILLER_128_487 ();
 sg13g2_decap_8 FILLER_128_494 ();
 sg13g2_decap_8 FILLER_128_501 ();
 sg13g2_decap_8 FILLER_128_508 ();
 sg13g2_decap_8 FILLER_128_515 ();
 sg13g2_decap_4 FILLER_128_522 ();
 sg13g2_fill_2 FILLER_128_526 ();
 sg13g2_decap_4 FILLER_128_548 ();
 sg13g2_fill_2 FILLER_128_552 ();
 sg13g2_decap_4 FILLER_128_559 ();
 sg13g2_decap_8 FILLER_128_572 ();
 sg13g2_decap_8 FILLER_128_579 ();
 sg13g2_decap_8 FILLER_128_586 ();
 sg13g2_fill_2 FILLER_128_593 ();
 sg13g2_decap_8 FILLER_128_611 ();
 sg13g2_decap_8 FILLER_128_618 ();
 sg13g2_decap_8 FILLER_128_625 ();
 sg13g2_decap_8 FILLER_128_632 ();
 sg13g2_fill_2 FILLER_128_639 ();
 sg13g2_fill_1 FILLER_128_641 ();
 sg13g2_decap_8 FILLER_128_655 ();
 sg13g2_decap_4 FILLER_128_662 ();
 sg13g2_fill_1 FILLER_128_666 ();
 sg13g2_decap_8 FILLER_128_687 ();
 sg13g2_decap_8 FILLER_128_694 ();
 sg13g2_decap_8 FILLER_128_701 ();
 sg13g2_decap_8 FILLER_128_708 ();
 sg13g2_decap_8 FILLER_128_715 ();
 sg13g2_decap_8 FILLER_128_722 ();
 sg13g2_fill_1 FILLER_128_729 ();
 sg13g2_decap_8 FILLER_128_744 ();
 sg13g2_decap_8 FILLER_128_751 ();
 sg13g2_decap_4 FILLER_128_758 ();
 sg13g2_decap_8 FILLER_128_766 ();
 sg13g2_decap_8 FILLER_128_785 ();
 sg13g2_fill_2 FILLER_128_792 ();
 sg13g2_decap_8 FILLER_128_799 ();
 sg13g2_decap_8 FILLER_128_806 ();
 sg13g2_decap_8 FILLER_128_813 ();
 sg13g2_decap_8 FILLER_128_820 ();
 sg13g2_decap_8 FILLER_128_827 ();
 sg13g2_decap_4 FILLER_128_834 ();
 sg13g2_fill_1 FILLER_128_838 ();
 sg13g2_decap_8 FILLER_128_884 ();
 sg13g2_decap_8 FILLER_128_891 ();
 sg13g2_decap_4 FILLER_128_898 ();
 sg13g2_fill_1 FILLER_128_902 ();
 sg13g2_decap_8 FILLER_128_918 ();
 sg13g2_fill_2 FILLER_128_925 ();
 sg13g2_fill_1 FILLER_128_927 ();
 sg13g2_decap_8 FILLER_128_933 ();
 sg13g2_decap_4 FILLER_128_940 ();
 sg13g2_decap_8 FILLER_128_956 ();
 sg13g2_decap_8 FILLER_128_963 ();
 sg13g2_decap_8 FILLER_128_970 ();
 sg13g2_decap_8 FILLER_128_977 ();
 sg13g2_decap_4 FILLER_128_984 ();
 sg13g2_decap_8 FILLER_128_1016 ();
 sg13g2_decap_8 FILLER_128_1023 ();
 sg13g2_decap_8 FILLER_128_1030 ();
 sg13g2_fill_1 FILLER_128_1037 ();
 sg13g2_decap_8 FILLER_128_1057 ();
 sg13g2_decap_8 FILLER_128_1078 ();
 sg13g2_decap_4 FILLER_128_1085 ();
 sg13g2_decap_8 FILLER_128_1098 ();
 sg13g2_decap_8 FILLER_128_1105 ();
 sg13g2_decap_8 FILLER_128_1112 ();
 sg13g2_decap_4 FILLER_128_1119 ();
 sg13g2_fill_1 FILLER_128_1123 ();
 sg13g2_decap_8 FILLER_128_1132 ();
 sg13g2_decap_8 FILLER_128_1139 ();
 sg13g2_decap_8 FILLER_128_1146 ();
 sg13g2_decap_8 FILLER_128_1153 ();
 sg13g2_decap_4 FILLER_128_1160 ();
 sg13g2_fill_1 FILLER_128_1164 ();
 sg13g2_decap_8 FILLER_128_1168 ();
 sg13g2_decap_8 FILLER_128_1175 ();
 sg13g2_decap_8 FILLER_128_1182 ();
 sg13g2_fill_2 FILLER_128_1189 ();
 sg13g2_fill_2 FILLER_128_1200 ();
 sg13g2_fill_1 FILLER_128_1202 ();
 sg13g2_fill_2 FILLER_128_1213 ();
 sg13g2_decap_8 FILLER_128_1233 ();
 sg13g2_decap_8 FILLER_128_1240 ();
 sg13g2_decap_8 FILLER_128_1247 ();
 sg13g2_decap_8 FILLER_128_1270 ();
 sg13g2_decap_8 FILLER_128_1277 ();
 sg13g2_fill_2 FILLER_128_1284 ();
 sg13g2_fill_1 FILLER_128_1286 ();
 sg13g2_decap_8 FILLER_128_1296 ();
 sg13g2_fill_2 FILLER_128_1303 ();
 sg13g2_fill_1 FILLER_128_1305 ();
 sg13g2_decap_8 FILLER_128_1310 ();
 sg13g2_decap_8 FILLER_128_1317 ();
 sg13g2_decap_8 FILLER_128_1324 ();
 sg13g2_decap_8 FILLER_128_1331 ();
 sg13g2_decap_8 FILLER_128_1338 ();
 sg13g2_decap_8 FILLER_128_1345 ();
 sg13g2_fill_2 FILLER_128_1352 ();
 sg13g2_fill_1 FILLER_128_1354 ();
 sg13g2_decap_8 FILLER_128_1365 ();
 sg13g2_decap_8 FILLER_128_1372 ();
 sg13g2_decap_8 FILLER_128_1379 ();
 sg13g2_decap_8 FILLER_128_1386 ();
 sg13g2_decap_8 FILLER_128_1393 ();
 sg13g2_decap_8 FILLER_128_1400 ();
 sg13g2_decap_8 FILLER_128_1407 ();
 sg13g2_decap_4 FILLER_128_1414 ();
 sg13g2_decap_4 FILLER_128_1435 ();
 sg13g2_decap_8 FILLER_128_1464 ();
 sg13g2_decap_8 FILLER_128_1471 ();
 sg13g2_decap_8 FILLER_128_1478 ();
 sg13g2_fill_2 FILLER_128_1485 ();
 sg13g2_fill_1 FILLER_128_1487 ();
 sg13g2_decap_8 FILLER_128_1496 ();
 sg13g2_decap_8 FILLER_128_1503 ();
 sg13g2_decap_8 FILLER_128_1510 ();
 sg13g2_decap_8 FILLER_128_1517 ();
 sg13g2_decap_8 FILLER_128_1524 ();
 sg13g2_decap_8 FILLER_128_1531 ();
 sg13g2_decap_8 FILLER_128_1538 ();
 sg13g2_decap_8 FILLER_128_1545 ();
 sg13g2_decap_8 FILLER_128_1552 ();
 sg13g2_decap_8 FILLER_128_1559 ();
 sg13g2_decap_8 FILLER_128_1566 ();
 sg13g2_decap_8 FILLER_128_1573 ();
 sg13g2_decap_8 FILLER_128_1580 ();
 sg13g2_decap_8 FILLER_128_1587 ();
 sg13g2_decap_8 FILLER_128_1594 ();
 sg13g2_decap_8 FILLER_128_1601 ();
 sg13g2_fill_1 FILLER_128_1608 ();
 sg13g2_decap_8 FILLER_128_1632 ();
 sg13g2_decap_8 FILLER_128_1639 ();
 sg13g2_decap_8 FILLER_128_1646 ();
 sg13g2_decap_4 FILLER_128_1653 ();
 sg13g2_fill_2 FILLER_128_1660 ();
 sg13g2_fill_1 FILLER_128_1662 ();
 sg13g2_decap_8 FILLER_128_1667 ();
 sg13g2_fill_1 FILLER_128_1674 ();
 sg13g2_decap_8 FILLER_128_1678 ();
 sg13g2_decap_8 FILLER_128_1685 ();
 sg13g2_decap_8 FILLER_128_1692 ();
 sg13g2_decap_8 FILLER_128_1699 ();
 sg13g2_decap_8 FILLER_128_1706 ();
 sg13g2_decap_4 FILLER_128_1713 ();
 sg13g2_fill_1 FILLER_128_1717 ();
 sg13g2_fill_1 FILLER_128_1723 ();
 sg13g2_decap_8 FILLER_128_1736 ();
 sg13g2_decap_8 FILLER_128_1743 ();
 sg13g2_decap_8 FILLER_128_1750 ();
 sg13g2_decap_8 FILLER_128_1757 ();
 sg13g2_decap_4 FILLER_128_1764 ();
 sg13g2_decap_8 FILLER_129_0 ();
 sg13g2_decap_4 FILLER_129_7 ();
 sg13g2_fill_1 FILLER_129_11 ();
 sg13g2_decap_8 FILLER_129_42 ();
 sg13g2_decap_8 FILLER_129_49 ();
 sg13g2_fill_2 FILLER_129_56 ();
 sg13g2_fill_1 FILLER_129_58 ();
 sg13g2_decap_8 FILLER_129_64 ();
 sg13g2_fill_2 FILLER_129_71 ();
 sg13g2_fill_2 FILLER_129_78 ();
 sg13g2_fill_1 FILLER_129_80 ();
 sg13g2_decap_8 FILLER_129_85 ();
 sg13g2_decap_8 FILLER_129_92 ();
 sg13g2_decap_8 FILLER_129_99 ();
 sg13g2_fill_2 FILLER_129_106 ();
 sg13g2_decap_8 FILLER_129_112 ();
 sg13g2_fill_2 FILLER_129_119 ();
 sg13g2_fill_1 FILLER_129_121 ();
 sg13g2_decap_8 FILLER_129_133 ();
 sg13g2_decap_8 FILLER_129_140 ();
 sg13g2_decap_8 FILLER_129_147 ();
 sg13g2_fill_2 FILLER_129_162 ();
 sg13g2_fill_1 FILLER_129_164 ();
 sg13g2_decap_8 FILLER_129_186 ();
 sg13g2_decap_8 FILLER_129_193 ();
 sg13g2_decap_4 FILLER_129_200 ();
 sg13g2_fill_2 FILLER_129_204 ();
 sg13g2_decap_8 FILLER_129_210 ();
 sg13g2_decap_8 FILLER_129_217 ();
 sg13g2_fill_2 FILLER_129_224 ();
 sg13g2_decap_8 FILLER_129_242 ();
 sg13g2_decap_8 FILLER_129_249 ();
 sg13g2_fill_2 FILLER_129_256 ();
 sg13g2_decap_8 FILLER_129_271 ();
 sg13g2_decap_8 FILLER_129_278 ();
 sg13g2_fill_2 FILLER_129_285 ();
 sg13g2_fill_1 FILLER_129_287 ();
 sg13g2_decap_8 FILLER_129_292 ();
 sg13g2_decap_8 FILLER_129_299 ();
 sg13g2_decap_8 FILLER_129_306 ();
 sg13g2_decap_4 FILLER_129_313 ();
 sg13g2_fill_1 FILLER_129_317 ();
 sg13g2_decap_4 FILLER_129_330 ();
 sg13g2_fill_1 FILLER_129_334 ();
 sg13g2_decap_8 FILLER_129_351 ();
 sg13g2_fill_2 FILLER_129_358 ();
 sg13g2_decap_8 FILLER_129_368 ();
 sg13g2_decap_8 FILLER_129_375 ();
 sg13g2_decap_8 FILLER_129_382 ();
 sg13g2_decap_8 FILLER_129_389 ();
 sg13g2_decap_4 FILLER_129_396 ();
 sg13g2_fill_2 FILLER_129_400 ();
 sg13g2_decap_8 FILLER_129_436 ();
 sg13g2_decap_8 FILLER_129_443 ();
 sg13g2_fill_2 FILLER_129_450 ();
 sg13g2_fill_1 FILLER_129_457 ();
 sg13g2_decap_8 FILLER_129_472 ();
 sg13g2_decap_8 FILLER_129_479 ();
 sg13g2_decap_8 FILLER_129_486 ();
 sg13g2_decap_8 FILLER_129_493 ();
 sg13g2_decap_4 FILLER_129_500 ();
 sg13g2_decap_8 FILLER_129_508 ();
 sg13g2_decap_8 FILLER_129_515 ();
 sg13g2_decap_8 FILLER_129_522 ();
 sg13g2_decap_8 FILLER_129_529 ();
 sg13g2_decap_8 FILLER_129_536 ();
 sg13g2_decap_8 FILLER_129_543 ();
 sg13g2_decap_8 FILLER_129_550 ();
 sg13g2_decap_8 FILLER_129_557 ();
 sg13g2_decap_8 FILLER_129_564 ();
 sg13g2_decap_8 FILLER_129_571 ();
 sg13g2_decap_8 FILLER_129_578 ();
 sg13g2_decap_8 FILLER_129_585 ();
 sg13g2_decap_8 FILLER_129_592 ();
 sg13g2_decap_8 FILLER_129_599 ();
 sg13g2_decap_8 FILLER_129_606 ();
 sg13g2_decap_4 FILLER_129_613 ();
 sg13g2_fill_2 FILLER_129_617 ();
 sg13g2_decap_8 FILLER_129_623 ();
 sg13g2_decap_8 FILLER_129_630 ();
 sg13g2_fill_2 FILLER_129_637 ();
 sg13g2_decap_8 FILLER_129_654 ();
 sg13g2_decap_8 FILLER_129_661 ();
 sg13g2_decap_8 FILLER_129_668 ();
 sg13g2_decap_8 FILLER_129_692 ();
 sg13g2_decap_8 FILLER_129_699 ();
 sg13g2_decap_8 FILLER_129_706 ();
 sg13g2_decap_4 FILLER_129_713 ();
 sg13g2_decap_8 FILLER_129_736 ();
 sg13g2_decap_8 FILLER_129_743 ();
 sg13g2_decap_8 FILLER_129_775 ();
 sg13g2_decap_8 FILLER_129_782 ();
 sg13g2_decap_8 FILLER_129_789 ();
 sg13g2_decap_8 FILLER_129_796 ();
 sg13g2_decap_8 FILLER_129_803 ();
 sg13g2_decap_8 FILLER_129_810 ();
 sg13g2_decap_8 FILLER_129_817 ();
 sg13g2_decap_8 FILLER_129_824 ();
 sg13g2_fill_1 FILLER_129_831 ();
 sg13g2_decap_4 FILLER_129_840 ();
 sg13g2_fill_1 FILLER_129_844 ();
 sg13g2_decap_8 FILLER_129_870 ();
 sg13g2_decap_8 FILLER_129_877 ();
 sg13g2_decap_8 FILLER_129_884 ();
 sg13g2_decap_8 FILLER_129_891 ();
 sg13g2_decap_8 FILLER_129_898 ();
 sg13g2_decap_8 FILLER_129_905 ();
 sg13g2_decap_8 FILLER_129_912 ();
 sg13g2_decap_8 FILLER_129_919 ();
 sg13g2_decap_8 FILLER_129_926 ();
 sg13g2_decap_8 FILLER_129_959 ();
 sg13g2_decap_8 FILLER_129_966 ();
 sg13g2_decap_8 FILLER_129_973 ();
 sg13g2_decap_8 FILLER_129_980 ();
 sg13g2_decap_8 FILLER_129_987 ();
 sg13g2_decap_8 FILLER_129_994 ();
 sg13g2_decap_4 FILLER_129_1001 ();
 sg13g2_fill_1 FILLER_129_1005 ();
 sg13g2_decap_8 FILLER_129_1020 ();
 sg13g2_decap_8 FILLER_129_1027 ();
 sg13g2_decap_4 FILLER_129_1034 ();
 sg13g2_fill_2 FILLER_129_1038 ();
 sg13g2_decap_8 FILLER_129_1058 ();
 sg13g2_decap_8 FILLER_129_1065 ();
 sg13g2_decap_8 FILLER_129_1072 ();
 sg13g2_fill_2 FILLER_129_1079 ();
 sg13g2_fill_2 FILLER_129_1089 ();
 sg13g2_fill_1 FILLER_129_1091 ();
 sg13g2_decap_8 FILLER_129_1104 ();
 sg13g2_decap_8 FILLER_129_1111 ();
 sg13g2_decap_8 FILLER_129_1118 ();
 sg13g2_fill_2 FILLER_129_1125 ();
 sg13g2_decap_8 FILLER_129_1141 ();
 sg13g2_decap_8 FILLER_129_1148 ();
 sg13g2_decap_8 FILLER_129_1155 ();
 sg13g2_fill_2 FILLER_129_1162 ();
 sg13g2_fill_1 FILLER_129_1164 ();
 sg13g2_decap_8 FILLER_129_1172 ();
 sg13g2_decap_8 FILLER_129_1179 ();
 sg13g2_decap_8 FILLER_129_1186 ();
 sg13g2_decap_8 FILLER_129_1193 ();
 sg13g2_decap_4 FILLER_129_1200 ();
 sg13g2_fill_1 FILLER_129_1204 ();
 sg13g2_decap_8 FILLER_129_1218 ();
 sg13g2_decap_8 FILLER_129_1225 ();
 sg13g2_fill_1 FILLER_129_1232 ();
 sg13g2_fill_1 FILLER_129_1255 ();
 sg13g2_decap_8 FILLER_129_1269 ();
 sg13g2_decap_8 FILLER_129_1276 ();
 sg13g2_decap_8 FILLER_129_1283 ();
 sg13g2_decap_8 FILLER_129_1290 ();
 sg13g2_decap_4 FILLER_129_1297 ();
 sg13g2_fill_1 FILLER_129_1305 ();
 sg13g2_decap_8 FILLER_129_1326 ();
 sg13g2_decap_8 FILLER_129_1333 ();
 sg13g2_decap_8 FILLER_129_1340 ();
 sg13g2_decap_8 FILLER_129_1347 ();
 sg13g2_fill_2 FILLER_129_1354 ();
 sg13g2_decap_8 FILLER_129_1389 ();
 sg13g2_decap_8 FILLER_129_1396 ();
 sg13g2_decap_8 FILLER_129_1403 ();
 sg13g2_decap_4 FILLER_129_1410 ();
 sg13g2_fill_1 FILLER_129_1414 ();
 sg13g2_decap_8 FILLER_129_1423 ();
 sg13g2_decap_8 FILLER_129_1430 ();
 sg13g2_fill_2 FILLER_129_1437 ();
 sg13g2_decap_8 FILLER_129_1454 ();
 sg13g2_decap_8 FILLER_129_1461 ();
 sg13g2_decap_8 FILLER_129_1468 ();
 sg13g2_decap_4 FILLER_129_1475 ();
 sg13g2_decap_8 FILLER_129_1484 ();
 sg13g2_decap_4 FILLER_129_1491 ();
 sg13g2_fill_2 FILLER_129_1495 ();
 sg13g2_decap_8 FILLER_129_1506 ();
 sg13g2_decap_8 FILLER_129_1513 ();
 sg13g2_decap_8 FILLER_129_1520 ();
 sg13g2_decap_8 FILLER_129_1527 ();
 sg13g2_decap_8 FILLER_129_1534 ();
 sg13g2_fill_2 FILLER_129_1541 ();
 sg13g2_fill_1 FILLER_129_1543 ();
 sg13g2_decap_8 FILLER_129_1557 ();
 sg13g2_decap_8 FILLER_129_1564 ();
 sg13g2_decap_8 FILLER_129_1571 ();
 sg13g2_decap_8 FILLER_129_1578 ();
 sg13g2_decap_8 FILLER_129_1585 ();
 sg13g2_decap_8 FILLER_129_1592 ();
 sg13g2_decap_8 FILLER_129_1599 ();
 sg13g2_decap_8 FILLER_129_1606 ();
 sg13g2_decap_4 FILLER_129_1613 ();
 sg13g2_fill_1 FILLER_129_1617 ();
 sg13g2_fill_2 FILLER_129_1622 ();
 sg13g2_decap_8 FILLER_129_1636 ();
 sg13g2_decap_8 FILLER_129_1643 ();
 sg13g2_fill_2 FILLER_129_1650 ();
 sg13g2_fill_1 FILLER_129_1652 ();
 sg13g2_fill_2 FILLER_129_1661 ();
 sg13g2_decap_8 FILLER_129_1688 ();
 sg13g2_decap_8 FILLER_129_1695 ();
 sg13g2_decap_8 FILLER_129_1702 ();
 sg13g2_decap_8 FILLER_129_1709 ();
 sg13g2_decap_4 FILLER_129_1716 ();
 sg13g2_fill_2 FILLER_129_1720 ();
 sg13g2_decap_8 FILLER_129_1726 ();
 sg13g2_decap_8 FILLER_129_1733 ();
 sg13g2_fill_1 FILLER_129_1740 ();
 sg13g2_decap_8 FILLER_129_1746 ();
 sg13g2_decap_8 FILLER_129_1753 ();
 sg13g2_decap_8 FILLER_129_1760 ();
 sg13g2_fill_1 FILLER_129_1767 ();
 sg13g2_decap_8 FILLER_130_0 ();
 sg13g2_decap_8 FILLER_130_7 ();
 sg13g2_decap_4 FILLER_130_14 ();
 sg13g2_fill_2 FILLER_130_22 ();
 sg13g2_fill_1 FILLER_130_24 ();
 sg13g2_decap_8 FILLER_130_33 ();
 sg13g2_decap_8 FILLER_130_40 ();
 sg13g2_fill_1 FILLER_130_47 ();
 sg13g2_decap_8 FILLER_130_75 ();
 sg13g2_decap_8 FILLER_130_82 ();
 sg13g2_decap_8 FILLER_130_89 ();
 sg13g2_decap_8 FILLER_130_96 ();
 sg13g2_fill_1 FILLER_130_103 ();
 sg13g2_decap_8 FILLER_130_127 ();
 sg13g2_decap_8 FILLER_130_134 ();
 sg13g2_fill_1 FILLER_130_141 ();
 sg13g2_decap_8 FILLER_130_151 ();
 sg13g2_fill_1 FILLER_130_158 ();
 sg13g2_decap_8 FILLER_130_166 ();
 sg13g2_decap_4 FILLER_130_173 ();
 sg13g2_fill_1 FILLER_130_177 ();
 sg13g2_decap_8 FILLER_130_183 ();
 sg13g2_decap_8 FILLER_130_190 ();
 sg13g2_decap_8 FILLER_130_197 ();
 sg13g2_decap_8 FILLER_130_204 ();
 sg13g2_decap_8 FILLER_130_211 ();
 sg13g2_decap_8 FILLER_130_218 ();
 sg13g2_decap_4 FILLER_130_225 ();
 sg13g2_fill_1 FILLER_130_229 ();
 sg13g2_fill_2 FILLER_130_238 ();
 sg13g2_decap_8 FILLER_130_245 ();
 sg13g2_decap_8 FILLER_130_252 ();
 sg13g2_decap_8 FILLER_130_259 ();
 sg13g2_decap_8 FILLER_130_266 ();
 sg13g2_fill_2 FILLER_130_273 ();
 sg13g2_fill_1 FILLER_130_275 ();
 sg13g2_decap_8 FILLER_130_281 ();
 sg13g2_decap_8 FILLER_130_288 ();
 sg13g2_decap_4 FILLER_130_295 ();
 sg13g2_decap_8 FILLER_130_308 ();
 sg13g2_decap_8 FILLER_130_315 ();
 sg13g2_decap_8 FILLER_130_322 ();
 sg13g2_fill_2 FILLER_130_329 ();
 sg13g2_fill_1 FILLER_130_331 ();
 sg13g2_decap_8 FILLER_130_337 ();
 sg13g2_decap_8 FILLER_130_344 ();
 sg13g2_decap_8 FILLER_130_351 ();
 sg13g2_fill_1 FILLER_130_358 ();
 sg13g2_fill_2 FILLER_130_368 ();
 sg13g2_fill_1 FILLER_130_370 ();
 sg13g2_fill_2 FILLER_130_387 ();
 sg13g2_decap_8 FILLER_130_397 ();
 sg13g2_decap_8 FILLER_130_404 ();
 sg13g2_fill_1 FILLER_130_411 ();
 sg13g2_fill_2 FILLER_130_425 ();
 sg13g2_decap_8 FILLER_130_439 ();
 sg13g2_decap_8 FILLER_130_446 ();
 sg13g2_decap_8 FILLER_130_453 ();
 sg13g2_fill_2 FILLER_130_460 ();
 sg13g2_decap_8 FILLER_130_470 ();
 sg13g2_decap_8 FILLER_130_477 ();
 sg13g2_decap_8 FILLER_130_484 ();
 sg13g2_fill_2 FILLER_130_491 ();
 sg13g2_fill_1 FILLER_130_493 ();
 sg13g2_decap_8 FILLER_130_499 ();
 sg13g2_decap_8 FILLER_130_506 ();
 sg13g2_decap_8 FILLER_130_513 ();
 sg13g2_decap_8 FILLER_130_520 ();
 sg13g2_decap_8 FILLER_130_527 ();
 sg13g2_decap_8 FILLER_130_534 ();
 sg13g2_decap_4 FILLER_130_541 ();
 sg13g2_fill_1 FILLER_130_545 ();
 sg13g2_fill_2 FILLER_130_556 ();
 sg13g2_fill_2 FILLER_130_563 ();
 sg13g2_fill_1 FILLER_130_565 ();
 sg13g2_decap_8 FILLER_130_572 ();
 sg13g2_fill_2 FILLER_130_579 ();
 sg13g2_decap_4 FILLER_130_589 ();
 sg13g2_fill_1 FILLER_130_593 ();
 sg13g2_fill_1 FILLER_130_606 ();
 sg13g2_fill_2 FILLER_130_613 ();
 sg13g2_decap_8 FILLER_130_625 ();
 sg13g2_decap_8 FILLER_130_632 ();
 sg13g2_fill_2 FILLER_130_639 ();
 sg13g2_fill_1 FILLER_130_641 ();
 sg13g2_decap_8 FILLER_130_645 ();
 sg13g2_decap_8 FILLER_130_652 ();
 sg13g2_decap_8 FILLER_130_659 ();
 sg13g2_decap_8 FILLER_130_666 ();
 sg13g2_decap_8 FILLER_130_673 ();
 sg13g2_decap_8 FILLER_130_684 ();
 sg13g2_decap_8 FILLER_130_691 ();
 sg13g2_decap_8 FILLER_130_698 ();
 sg13g2_decap_8 FILLER_130_705 ();
 sg13g2_decap_8 FILLER_130_712 ();
 sg13g2_decap_4 FILLER_130_719 ();
 sg13g2_decap_4 FILLER_130_731 ();
 sg13g2_fill_1 FILLER_130_735 ();
 sg13g2_decap_8 FILLER_130_740 ();
 sg13g2_fill_2 FILLER_130_747 ();
 sg13g2_fill_1 FILLER_130_749 ();
 sg13g2_decap_8 FILLER_130_766 ();
 sg13g2_decap_8 FILLER_130_773 ();
 sg13g2_decap_8 FILLER_130_780 ();
 sg13g2_decap_8 FILLER_130_787 ();
 sg13g2_decap_8 FILLER_130_794 ();
 sg13g2_fill_2 FILLER_130_801 ();
 sg13g2_decap_8 FILLER_130_815 ();
 sg13g2_decap_8 FILLER_130_822 ();
 sg13g2_decap_8 FILLER_130_829 ();
 sg13g2_decap_8 FILLER_130_836 ();
 sg13g2_decap_8 FILLER_130_843 ();
 sg13g2_fill_1 FILLER_130_850 ();
 sg13g2_decap_8 FILLER_130_859 ();
 sg13g2_decap_8 FILLER_130_866 ();
 sg13g2_decap_8 FILLER_130_873 ();
 sg13g2_decap_8 FILLER_130_880 ();
 sg13g2_decap_8 FILLER_130_887 ();
 sg13g2_decap_8 FILLER_130_894 ();
 sg13g2_decap_8 FILLER_130_901 ();
 sg13g2_decap_8 FILLER_130_908 ();
 sg13g2_decap_8 FILLER_130_915 ();
 sg13g2_decap_8 FILLER_130_922 ();
 sg13g2_decap_4 FILLER_130_929 ();
 sg13g2_fill_1 FILLER_130_933 ();
 sg13g2_fill_1 FILLER_130_945 ();
 sg13g2_decap_8 FILLER_130_950 ();
 sg13g2_decap_8 FILLER_130_957 ();
 sg13g2_decap_8 FILLER_130_964 ();
 sg13g2_fill_2 FILLER_130_971 ();
 sg13g2_fill_1 FILLER_130_973 ();
 sg13g2_decap_8 FILLER_130_980 ();
 sg13g2_decap_8 FILLER_130_987 ();
 sg13g2_decap_8 FILLER_130_994 ();
 sg13g2_decap_8 FILLER_130_1001 ();
 sg13g2_fill_2 FILLER_130_1008 ();
 sg13g2_decap_8 FILLER_130_1014 ();
 sg13g2_decap_8 FILLER_130_1021 ();
 sg13g2_decap_8 FILLER_130_1028 ();
 sg13g2_decap_8 FILLER_130_1035 ();
 sg13g2_fill_1 FILLER_130_1042 ();
 sg13g2_fill_1 FILLER_130_1056 ();
 sg13g2_decap_8 FILLER_130_1070 ();
 sg13g2_decap_8 FILLER_130_1077 ();
 sg13g2_decap_8 FILLER_130_1090 ();
 sg13g2_decap_8 FILLER_130_1097 ();
 sg13g2_decap_8 FILLER_130_1104 ();
 sg13g2_fill_2 FILLER_130_1111 ();
 sg13g2_decap_8 FILLER_130_1125 ();
 sg13g2_decap_8 FILLER_130_1132 ();
 sg13g2_decap_8 FILLER_130_1139 ();
 sg13g2_fill_2 FILLER_130_1146 ();
 sg13g2_decap_4 FILLER_130_1166 ();
 sg13g2_fill_2 FILLER_130_1186 ();
 sg13g2_fill_1 FILLER_130_1188 ();
 sg13g2_decap_8 FILLER_130_1202 ();
 sg13g2_decap_4 FILLER_130_1209 ();
 sg13g2_fill_2 FILLER_130_1213 ();
 sg13g2_decap_8 FILLER_130_1223 ();
 sg13g2_decap_8 FILLER_130_1230 ();
 sg13g2_decap_8 FILLER_130_1237 ();
 sg13g2_decap_8 FILLER_130_1244 ();
 sg13g2_decap_8 FILLER_130_1251 ();
 sg13g2_fill_2 FILLER_130_1258 ();
 sg13g2_fill_1 FILLER_130_1260 ();
 sg13g2_decap_8 FILLER_130_1269 ();
 sg13g2_decap_8 FILLER_130_1276 ();
 sg13g2_fill_2 FILLER_130_1283 ();
 sg13g2_fill_1 FILLER_130_1285 ();
 sg13g2_fill_1 FILLER_130_1311 ();
 sg13g2_decap_8 FILLER_130_1317 ();
 sg13g2_decap_8 FILLER_130_1324 ();
 sg13g2_decap_8 FILLER_130_1331 ();
 sg13g2_decap_8 FILLER_130_1338 ();
 sg13g2_decap_8 FILLER_130_1345 ();
 sg13g2_decap_4 FILLER_130_1352 ();
 sg13g2_decap_8 FILLER_130_1369 ();
 sg13g2_decap_4 FILLER_130_1376 ();
 sg13g2_fill_2 FILLER_130_1380 ();
 sg13g2_fill_1 FILLER_130_1399 ();
 sg13g2_decap_8 FILLER_130_1406 ();
 sg13g2_decap_8 FILLER_130_1413 ();
 sg13g2_decap_8 FILLER_130_1420 ();
 sg13g2_decap_8 FILLER_130_1427 ();
 sg13g2_decap_8 FILLER_130_1434 ();
 sg13g2_fill_2 FILLER_130_1441 ();
 sg13g2_decap_4 FILLER_130_1448 ();
 sg13g2_fill_2 FILLER_130_1452 ();
 sg13g2_decap_8 FILLER_130_1459 ();
 sg13g2_decap_8 FILLER_130_1466 ();
 sg13g2_decap_8 FILLER_130_1473 ();
 sg13g2_decap_8 FILLER_130_1480 ();
 sg13g2_decap_8 FILLER_130_1491 ();
 sg13g2_decap_8 FILLER_130_1502 ();
 sg13g2_decap_8 FILLER_130_1509 ();
 sg13g2_decap_8 FILLER_130_1516 ();
 sg13g2_decap_8 FILLER_130_1523 ();
 sg13g2_fill_1 FILLER_130_1547 ();
 sg13g2_decap_8 FILLER_130_1574 ();
 sg13g2_decap_8 FILLER_130_1581 ();
 sg13g2_decap_8 FILLER_130_1588 ();
 sg13g2_decap_8 FILLER_130_1595 ();
 sg13g2_decap_8 FILLER_130_1602 ();
 sg13g2_decap_8 FILLER_130_1609 ();
 sg13g2_decap_8 FILLER_130_1616 ();
 sg13g2_decap_8 FILLER_130_1623 ();
 sg13g2_decap_8 FILLER_130_1630 ();
 sg13g2_decap_8 FILLER_130_1637 ();
 sg13g2_decap_8 FILLER_130_1644 ();
 sg13g2_fill_2 FILLER_130_1651 ();
 sg13g2_fill_1 FILLER_130_1653 ();
 sg13g2_decap_4 FILLER_130_1662 ();
 sg13g2_fill_2 FILLER_130_1666 ();
 sg13g2_decap_8 FILLER_130_1686 ();
 sg13g2_decap_8 FILLER_130_1693 ();
 sg13g2_decap_8 FILLER_130_1700 ();
 sg13g2_decap_8 FILLER_130_1707 ();
 sg13g2_decap_8 FILLER_130_1714 ();
 sg13g2_decap_8 FILLER_130_1721 ();
 sg13g2_decap_4 FILLER_130_1728 ();
 sg13g2_fill_1 FILLER_130_1732 ();
 sg13g2_decap_8 FILLER_130_1759 ();
 sg13g2_fill_2 FILLER_130_1766 ();
 sg13g2_decap_8 FILLER_131_0 ();
 sg13g2_decap_8 FILLER_131_7 ();
 sg13g2_decap_8 FILLER_131_14 ();
 sg13g2_decap_8 FILLER_131_21 ();
 sg13g2_decap_8 FILLER_131_28 ();
 sg13g2_decap_8 FILLER_131_35 ();
 sg13g2_decap_8 FILLER_131_42 ();
 sg13g2_decap_8 FILLER_131_49 ();
 sg13g2_decap_4 FILLER_131_56 ();
 sg13g2_decap_8 FILLER_131_79 ();
 sg13g2_decap_8 FILLER_131_86 ();
 sg13g2_decap_8 FILLER_131_93 ();
 sg13g2_decap_8 FILLER_131_100 ();
 sg13g2_decap_8 FILLER_131_107 ();
 sg13g2_decap_8 FILLER_131_114 ();
 sg13g2_decap_8 FILLER_131_121 ();
 sg13g2_decap_8 FILLER_131_128 ();
 sg13g2_fill_2 FILLER_131_135 ();
 sg13g2_fill_2 FILLER_131_145 ();
 sg13g2_decap_8 FILLER_131_151 ();
 sg13g2_decap_8 FILLER_131_158 ();
 sg13g2_decap_8 FILLER_131_165 ();
 sg13g2_fill_2 FILLER_131_172 ();
 sg13g2_decap_8 FILLER_131_184 ();
 sg13g2_decap_8 FILLER_131_191 ();
 sg13g2_decap_8 FILLER_131_198 ();
 sg13g2_decap_8 FILLER_131_205 ();
 sg13g2_fill_2 FILLER_131_212 ();
 sg13g2_fill_1 FILLER_131_214 ();
 sg13g2_decap_4 FILLER_131_223 ();
 sg13g2_fill_1 FILLER_131_227 ();
 sg13g2_decap_4 FILLER_131_232 ();
 sg13g2_fill_2 FILLER_131_236 ();
 sg13g2_decap_8 FILLER_131_247 ();
 sg13g2_fill_2 FILLER_131_254 ();
 sg13g2_decap_8 FILLER_131_259 ();
 sg13g2_decap_4 FILLER_131_266 ();
 sg13g2_fill_2 FILLER_131_270 ();
 sg13g2_fill_2 FILLER_131_287 ();
 sg13g2_fill_2 FILLER_131_297 ();
 sg13g2_fill_1 FILLER_131_299 ();
 sg13g2_decap_8 FILLER_131_311 ();
 sg13g2_decap_8 FILLER_131_318 ();
 sg13g2_decap_8 FILLER_131_325 ();
 sg13g2_decap_8 FILLER_131_332 ();
 sg13g2_decap_8 FILLER_131_339 ();
 sg13g2_decap_8 FILLER_131_346 ();
 sg13g2_decap_4 FILLER_131_379 ();
 sg13g2_fill_2 FILLER_131_383 ();
 sg13g2_decap_8 FILLER_131_402 ();
 sg13g2_decap_8 FILLER_131_409 ();
 sg13g2_decap_8 FILLER_131_416 ();
 sg13g2_decap_8 FILLER_131_423 ();
 sg13g2_fill_1 FILLER_131_430 ();
 sg13g2_decap_8 FILLER_131_436 ();
 sg13g2_decap_8 FILLER_131_443 ();
 sg13g2_fill_2 FILLER_131_450 ();
 sg13g2_fill_1 FILLER_131_452 ();
 sg13g2_decap_8 FILLER_131_457 ();
 sg13g2_decap_8 FILLER_131_464 ();
 sg13g2_decap_8 FILLER_131_471 ();
 sg13g2_fill_2 FILLER_131_478 ();
 sg13g2_fill_1 FILLER_131_480 ();
 sg13g2_fill_2 FILLER_131_502 ();
 sg13g2_fill_1 FILLER_131_504 ();
 sg13g2_decap_4 FILLER_131_514 ();
 sg13g2_fill_2 FILLER_131_518 ();
 sg13g2_decap_4 FILLER_131_528 ();
 sg13g2_fill_1 FILLER_131_532 ();
 sg13g2_decap_8 FILLER_131_547 ();
 sg13g2_decap_8 FILLER_131_554 ();
 sg13g2_decap_8 FILLER_131_561 ();
 sg13g2_fill_2 FILLER_131_568 ();
 sg13g2_fill_2 FILLER_131_584 ();
 sg13g2_decap_4 FILLER_131_605 ();
 sg13g2_fill_1 FILLER_131_609 ();
 sg13g2_decap_8 FILLER_131_623 ();
 sg13g2_fill_2 FILLER_131_630 ();
 sg13g2_fill_2 FILLER_131_640 ();
 sg13g2_fill_1 FILLER_131_642 ();
 sg13g2_decap_8 FILLER_131_655 ();
 sg13g2_decap_8 FILLER_131_662 ();
 sg13g2_fill_2 FILLER_131_669 ();
 sg13g2_decap_4 FILLER_131_692 ();
 sg13g2_fill_1 FILLER_131_696 ();
 sg13g2_decap_8 FILLER_131_710 ();
 sg13g2_decap_4 FILLER_131_717 ();
 sg13g2_fill_2 FILLER_131_721 ();
 sg13g2_fill_1 FILLER_131_728 ();
 sg13g2_decap_8 FILLER_131_734 ();
 sg13g2_fill_1 FILLER_131_741 ();
 sg13g2_decap_8 FILLER_131_751 ();
 sg13g2_decap_8 FILLER_131_758 ();
 sg13g2_decap_8 FILLER_131_774 ();
 sg13g2_decap_8 FILLER_131_781 ();
 sg13g2_decap_8 FILLER_131_788 ();
 sg13g2_fill_1 FILLER_131_795 ();
 sg13g2_decap_8 FILLER_131_821 ();
 sg13g2_decap_8 FILLER_131_828 ();
 sg13g2_decap_8 FILLER_131_835 ();
 sg13g2_decap_8 FILLER_131_842 ();
 sg13g2_decap_4 FILLER_131_849 ();
 sg13g2_decap_8 FILLER_131_861 ();
 sg13g2_fill_2 FILLER_131_868 ();
 sg13g2_decap_8 FILLER_131_878 ();
 sg13g2_decap_8 FILLER_131_885 ();
 sg13g2_decap_8 FILLER_131_892 ();
 sg13g2_decap_4 FILLER_131_899 ();
 sg13g2_fill_2 FILLER_131_903 ();
 sg13g2_decap_8 FILLER_131_909 ();
 sg13g2_decap_4 FILLER_131_916 ();
 sg13g2_fill_1 FILLER_131_920 ();
 sg13g2_decap_4 FILLER_131_928 ();
 sg13g2_fill_2 FILLER_131_932 ();
 sg13g2_decap_8 FILLER_131_953 ();
 sg13g2_decap_8 FILLER_131_960 ();
 sg13g2_decap_8 FILLER_131_967 ();
 sg13g2_decap_8 FILLER_131_974 ();
 sg13g2_decap_8 FILLER_131_981 ();
 sg13g2_decap_8 FILLER_131_988 ();
 sg13g2_decap_8 FILLER_131_995 ();
 sg13g2_decap_8 FILLER_131_1002 ();
 sg13g2_decap_8 FILLER_131_1009 ();
 sg13g2_decap_8 FILLER_131_1016 ();
 sg13g2_decap_8 FILLER_131_1023 ();
 sg13g2_decap_8 FILLER_131_1030 ();
 sg13g2_decap_8 FILLER_131_1037 ();
 sg13g2_decap_8 FILLER_131_1044 ();
 sg13g2_decap_8 FILLER_131_1051 ();
 sg13g2_decap_8 FILLER_131_1058 ();
 sg13g2_decap_8 FILLER_131_1065 ();
 sg13g2_decap_4 FILLER_131_1072 ();
 sg13g2_decap_8 FILLER_131_1093 ();
 sg13g2_decap_4 FILLER_131_1100 ();
 sg13g2_fill_2 FILLER_131_1104 ();
 sg13g2_decap_8 FILLER_131_1137 ();
 sg13g2_decap_8 FILLER_131_1144 ();
 sg13g2_fill_2 FILLER_131_1151 ();
 sg13g2_decap_8 FILLER_131_1160 ();
 sg13g2_fill_2 FILLER_131_1167 ();
 sg13g2_fill_1 FILLER_131_1169 ();
 sg13g2_decap_4 FILLER_131_1176 ();
 sg13g2_decap_8 FILLER_131_1206 ();
 sg13g2_decap_8 FILLER_131_1213 ();
 sg13g2_decap_8 FILLER_131_1220 ();
 sg13g2_decap_8 FILLER_131_1227 ();
 sg13g2_decap_8 FILLER_131_1234 ();
 sg13g2_fill_1 FILLER_131_1241 ();
 sg13g2_decap_8 FILLER_131_1247 ();
 sg13g2_decap_8 FILLER_131_1254 ();
 sg13g2_decap_8 FILLER_131_1261 ();
 sg13g2_decap_8 FILLER_131_1268 ();
 sg13g2_fill_1 FILLER_131_1275 ();
 sg13g2_decap_4 FILLER_131_1292 ();
 sg13g2_decap_8 FILLER_131_1316 ();
 sg13g2_decap_4 FILLER_131_1323 ();
 sg13g2_decap_8 FILLER_131_1331 ();
 sg13g2_decap_8 FILLER_131_1338 ();
 sg13g2_decap_8 FILLER_131_1345 ();
 sg13g2_decap_8 FILLER_131_1352 ();
 sg13g2_decap_8 FILLER_131_1359 ();
 sg13g2_decap_8 FILLER_131_1366 ();
 sg13g2_decap_8 FILLER_131_1373 ();
 sg13g2_decap_8 FILLER_131_1380 ();
 sg13g2_fill_1 FILLER_131_1387 ();
 sg13g2_fill_2 FILLER_131_1402 ();
 sg13g2_fill_1 FILLER_131_1404 ();
 sg13g2_decap_8 FILLER_131_1417 ();
 sg13g2_decap_8 FILLER_131_1424 ();
 sg13g2_decap_8 FILLER_131_1431 ();
 sg13g2_decap_8 FILLER_131_1438 ();
 sg13g2_fill_2 FILLER_131_1445 ();
 sg13g2_decap_8 FILLER_131_1455 ();
 sg13g2_fill_1 FILLER_131_1462 ();
 sg13g2_decap_8 FILLER_131_1471 ();
 sg13g2_decap_8 FILLER_131_1478 ();
 sg13g2_decap_8 FILLER_131_1514 ();
 sg13g2_decap_8 FILLER_131_1521 ();
 sg13g2_decap_8 FILLER_131_1528 ();
 sg13g2_decap_4 FILLER_131_1535 ();
 sg13g2_fill_2 FILLER_131_1539 ();
 sg13g2_decap_4 FILLER_131_1545 ();
 sg13g2_fill_2 FILLER_131_1549 ();
 sg13g2_fill_2 FILLER_131_1555 ();
 sg13g2_fill_1 FILLER_131_1557 ();
 sg13g2_decap_8 FILLER_131_1572 ();
 sg13g2_decap_8 FILLER_131_1579 ();
 sg13g2_fill_2 FILLER_131_1586 ();
 sg13g2_decap_8 FILLER_131_1592 ();
 sg13g2_decap_8 FILLER_131_1599 ();
 sg13g2_decap_8 FILLER_131_1606 ();
 sg13g2_decap_8 FILLER_131_1613 ();
 sg13g2_decap_8 FILLER_131_1620 ();
 sg13g2_decap_8 FILLER_131_1627 ();
 sg13g2_decap_8 FILLER_131_1634 ();
 sg13g2_decap_8 FILLER_131_1641 ();
 sg13g2_decap_8 FILLER_131_1648 ();
 sg13g2_decap_8 FILLER_131_1655 ();
 sg13g2_fill_2 FILLER_131_1662 ();
 sg13g2_fill_1 FILLER_131_1664 ();
 sg13g2_fill_1 FILLER_131_1673 ();
 sg13g2_decap_8 FILLER_131_1679 ();
 sg13g2_decap_8 FILLER_131_1686 ();
 sg13g2_decap_8 FILLER_131_1693 ();
 sg13g2_decap_8 FILLER_131_1700 ();
 sg13g2_decap_8 FILLER_131_1707 ();
 sg13g2_decap_8 FILLER_131_1714 ();
 sg13g2_decap_8 FILLER_131_1721 ();
 sg13g2_decap_8 FILLER_131_1728 ();
 sg13g2_fill_2 FILLER_131_1735 ();
 sg13g2_decap_8 FILLER_131_1749 ();
 sg13g2_decap_8 FILLER_131_1756 ();
 sg13g2_decap_4 FILLER_131_1763 ();
 sg13g2_fill_1 FILLER_131_1767 ();
 sg13g2_decap_8 FILLER_132_0 ();
 sg13g2_decap_8 FILLER_132_7 ();
 sg13g2_decap_8 FILLER_132_14 ();
 sg13g2_decap_8 FILLER_132_21 ();
 sg13g2_decap_8 FILLER_132_28 ();
 sg13g2_decap_8 FILLER_132_35 ();
 sg13g2_decap_8 FILLER_132_42 ();
 sg13g2_decap_4 FILLER_132_49 ();
 sg13g2_fill_1 FILLER_132_53 ();
 sg13g2_fill_2 FILLER_132_62 ();
 sg13g2_fill_1 FILLER_132_64 ();
 sg13g2_decap_8 FILLER_132_75 ();
 sg13g2_decap_8 FILLER_132_82 ();
 sg13g2_decap_8 FILLER_132_89 ();
 sg13g2_decap_8 FILLER_132_96 ();
 sg13g2_fill_1 FILLER_132_103 ();
 sg13g2_fill_1 FILLER_132_107 ();
 sg13g2_decap_8 FILLER_132_129 ();
 sg13g2_decap_8 FILLER_132_136 ();
 sg13g2_decap_8 FILLER_132_143 ();
 sg13g2_decap_8 FILLER_132_150 ();
 sg13g2_decap_8 FILLER_132_157 ();
 sg13g2_decap_4 FILLER_132_164 ();
 sg13g2_fill_2 FILLER_132_168 ();
 sg13g2_fill_2 FILLER_132_184 ();
 sg13g2_fill_1 FILLER_132_186 ();
 sg13g2_decap_8 FILLER_132_191 ();
 sg13g2_decap_8 FILLER_132_198 ();
 sg13g2_decap_8 FILLER_132_205 ();
 sg13g2_decap_8 FILLER_132_212 ();
 sg13g2_fill_1 FILLER_132_219 ();
 sg13g2_decap_8 FILLER_132_244 ();
 sg13g2_decap_4 FILLER_132_251 ();
 sg13g2_fill_1 FILLER_132_255 ();
 sg13g2_decap_8 FILLER_132_268 ();
 sg13g2_decap_8 FILLER_132_275 ();
 sg13g2_decap_4 FILLER_132_291 ();
 sg13g2_fill_1 FILLER_132_295 ();
 sg13g2_decap_4 FILLER_132_308 ();
 sg13g2_fill_2 FILLER_132_312 ();
 sg13g2_fill_1 FILLER_132_327 ();
 sg13g2_decap_8 FILLER_132_337 ();
 sg13g2_decap_8 FILLER_132_344 ();
 sg13g2_decap_8 FILLER_132_351 ();
 sg13g2_decap_8 FILLER_132_362 ();
 sg13g2_decap_4 FILLER_132_369 ();
 sg13g2_fill_1 FILLER_132_373 ();
 sg13g2_decap_4 FILLER_132_380 ();
 sg13g2_fill_1 FILLER_132_384 ();
 sg13g2_decap_8 FILLER_132_406 ();
 sg13g2_decap_8 FILLER_132_413 ();
 sg13g2_fill_2 FILLER_132_420 ();
 sg13g2_fill_1 FILLER_132_443 ();
 sg13g2_decap_8 FILLER_132_465 ();
 sg13g2_decap_8 FILLER_132_472 ();
 sg13g2_decap_8 FILLER_132_479 ();
 sg13g2_decap_8 FILLER_132_486 ();
 sg13g2_fill_2 FILLER_132_493 ();
 sg13g2_fill_1 FILLER_132_495 ();
 sg13g2_decap_8 FILLER_132_501 ();
 sg13g2_fill_1 FILLER_132_508 ();
 sg13g2_decap_8 FILLER_132_523 ();
 sg13g2_fill_2 FILLER_132_530 ();
 sg13g2_decap_8 FILLER_132_548 ();
 sg13g2_decap_8 FILLER_132_555 ();
 sg13g2_decap_8 FILLER_132_562 ();
 sg13g2_decap_8 FILLER_132_573 ();
 sg13g2_decap_8 FILLER_132_580 ();
 sg13g2_decap_8 FILLER_132_587 ();
 sg13g2_decap_8 FILLER_132_626 ();
 sg13g2_decap_8 FILLER_132_633 ();
 sg13g2_decap_8 FILLER_132_640 ();
 sg13g2_decap_8 FILLER_132_647 ();
 sg13g2_decap_8 FILLER_132_654 ();
 sg13g2_decap_8 FILLER_132_661 ();
 sg13g2_decap_8 FILLER_132_668 ();
 sg13g2_decap_8 FILLER_132_675 ();
 sg13g2_decap_8 FILLER_132_682 ();
 sg13g2_decap_8 FILLER_132_689 ();
 sg13g2_fill_2 FILLER_132_696 ();
 sg13g2_fill_1 FILLER_132_698 ();
 sg13g2_fill_1 FILLER_132_704 ();
 sg13g2_decap_8 FILLER_132_714 ();
 sg13g2_decap_8 FILLER_132_721 ();
 sg13g2_decap_8 FILLER_132_728 ();
 sg13g2_decap_8 FILLER_132_735 ();
 sg13g2_decap_4 FILLER_132_742 ();
 sg13g2_fill_1 FILLER_132_746 ();
 sg13g2_decap_4 FILLER_132_750 ();
 sg13g2_fill_2 FILLER_132_758 ();
 sg13g2_decap_8 FILLER_132_780 ();
 sg13g2_decap_8 FILLER_132_787 ();
 sg13g2_fill_2 FILLER_132_794 ();
 sg13g2_decap_8 FILLER_132_816 ();
 sg13g2_decap_8 FILLER_132_823 ();
 sg13g2_decap_8 FILLER_132_830 ();
 sg13g2_decap_8 FILLER_132_837 ();
 sg13g2_decap_8 FILLER_132_844 ();
 sg13g2_decap_8 FILLER_132_851 ();
 sg13g2_decap_8 FILLER_132_858 ();
 sg13g2_fill_2 FILLER_132_865 ();
 sg13g2_fill_2 FILLER_132_880 ();
 sg13g2_decap_4 FILLER_132_890 ();
 sg13g2_fill_1 FILLER_132_933 ();
 sg13g2_fill_1 FILLER_132_945 ();
 sg13g2_fill_2 FILLER_132_951 ();
 sg13g2_decap_8 FILLER_132_961 ();
 sg13g2_fill_1 FILLER_132_968 ();
 sg13g2_decap_8 FILLER_132_974 ();
 sg13g2_fill_1 FILLER_132_981 ();
 sg13g2_fill_2 FILLER_132_987 ();
 sg13g2_fill_1 FILLER_132_989 ();
 sg13g2_decap_4 FILLER_132_1003 ();
 sg13g2_fill_2 FILLER_132_1007 ();
 sg13g2_fill_1 FILLER_132_1013 ();
 sg13g2_decap_8 FILLER_132_1018 ();
 sg13g2_decap_8 FILLER_132_1025 ();
 sg13g2_decap_8 FILLER_132_1032 ();
 sg13g2_decap_8 FILLER_132_1039 ();
 sg13g2_decap_8 FILLER_132_1046 ();
 sg13g2_decap_8 FILLER_132_1053 ();
 sg13g2_decap_8 FILLER_132_1060 ();
 sg13g2_fill_2 FILLER_132_1067 ();
 sg13g2_fill_2 FILLER_132_1076 ();
 sg13g2_decap_8 FILLER_132_1098 ();
 sg13g2_fill_1 FILLER_132_1105 ();
 sg13g2_decap_4 FILLER_132_1116 ();
 sg13g2_fill_1 FILLER_132_1120 ();
 sg13g2_decap_8 FILLER_132_1133 ();
 sg13g2_decap_8 FILLER_132_1140 ();
 sg13g2_decap_8 FILLER_132_1147 ();
 sg13g2_decap_4 FILLER_132_1154 ();
 sg13g2_decap_4 FILLER_132_1183 ();
 sg13g2_fill_2 FILLER_132_1201 ();
 sg13g2_decap_8 FILLER_132_1215 ();
 sg13g2_decap_4 FILLER_132_1222 ();
 sg13g2_fill_1 FILLER_132_1226 ();
 sg13g2_decap_8 FILLER_132_1235 ();
 sg13g2_decap_8 FILLER_132_1242 ();
 sg13g2_decap_8 FILLER_132_1249 ();
 sg13g2_decap_8 FILLER_132_1256 ();
 sg13g2_decap_8 FILLER_132_1263 ();
 sg13g2_decap_4 FILLER_132_1270 ();
 sg13g2_fill_2 FILLER_132_1274 ();
 sg13g2_decap_4 FILLER_132_1288 ();
 sg13g2_decap_8 FILLER_132_1300 ();
 sg13g2_decap_8 FILLER_132_1307 ();
 sg13g2_decap_8 FILLER_132_1314 ();
 sg13g2_decap_4 FILLER_132_1321 ();
 sg13g2_fill_1 FILLER_132_1325 ();
 sg13g2_decap_8 FILLER_132_1336 ();
 sg13g2_decap_8 FILLER_132_1343 ();
 sg13g2_fill_2 FILLER_132_1350 ();
 sg13g2_fill_1 FILLER_132_1356 ();
 sg13g2_decap_8 FILLER_132_1361 ();
 sg13g2_decap_8 FILLER_132_1368 ();
 sg13g2_decap_8 FILLER_132_1375 ();
 sg13g2_decap_8 FILLER_132_1382 ();
 sg13g2_decap_8 FILLER_132_1389 ();
 sg13g2_fill_1 FILLER_132_1396 ();
 sg13g2_decap_8 FILLER_132_1406 ();
 sg13g2_decap_4 FILLER_132_1413 ();
 sg13g2_fill_1 FILLER_132_1417 ();
 sg13g2_decap_4 FILLER_132_1426 ();
 sg13g2_decap_8 FILLER_132_1434 ();
 sg13g2_decap_8 FILLER_132_1441 ();
 sg13g2_fill_1 FILLER_132_1448 ();
 sg13g2_decap_8 FILLER_132_1454 ();
 sg13g2_decap_8 FILLER_132_1461 ();
 sg13g2_decap_8 FILLER_132_1468 ();
 sg13g2_decap_8 FILLER_132_1475 ();
 sg13g2_decap_4 FILLER_132_1482 ();
 sg13g2_decap_8 FILLER_132_1516 ();
 sg13g2_decap_8 FILLER_132_1523 ();
 sg13g2_decap_8 FILLER_132_1530 ();
 sg13g2_decap_4 FILLER_132_1537 ();
 sg13g2_decap_8 FILLER_132_1561 ();
 sg13g2_decap_8 FILLER_132_1568 ();
 sg13g2_fill_2 FILLER_132_1575 ();
 sg13g2_fill_1 FILLER_132_1577 ();
 sg13g2_fill_2 FILLER_132_1604 ();
 sg13g2_fill_1 FILLER_132_1606 ();
 sg13g2_fill_1 FILLER_132_1611 ();
 sg13g2_decap_8 FILLER_132_1625 ();
 sg13g2_decap_8 FILLER_132_1632 ();
 sg13g2_decap_8 FILLER_132_1639 ();
 sg13g2_decap_8 FILLER_132_1646 ();
 sg13g2_fill_2 FILLER_132_1653 ();
 sg13g2_fill_1 FILLER_132_1655 ();
 sg13g2_decap_8 FILLER_132_1666 ();
 sg13g2_fill_1 FILLER_132_1673 ();
 sg13g2_decap_8 FILLER_132_1679 ();
 sg13g2_decap_8 FILLER_132_1686 ();
 sg13g2_decap_8 FILLER_132_1693 ();
 sg13g2_decap_8 FILLER_132_1700 ();
 sg13g2_decap_8 FILLER_132_1707 ();
 sg13g2_decap_8 FILLER_132_1714 ();
 sg13g2_decap_8 FILLER_132_1721 ();
 sg13g2_fill_2 FILLER_132_1728 ();
 sg13g2_decap_8 FILLER_132_1755 ();
 sg13g2_decap_4 FILLER_132_1762 ();
 sg13g2_fill_2 FILLER_132_1766 ();
 sg13g2_decap_8 FILLER_133_0 ();
 sg13g2_decap_8 FILLER_133_7 ();
 sg13g2_fill_2 FILLER_133_14 ();
 sg13g2_decap_8 FILLER_133_33 ();
 sg13g2_decap_8 FILLER_133_40 ();
 sg13g2_decap_8 FILLER_133_47 ();
 sg13g2_decap_8 FILLER_133_54 ();
 sg13g2_decap_8 FILLER_133_61 ();
 sg13g2_decap_8 FILLER_133_68 ();
 sg13g2_decap_8 FILLER_133_75 ();
 sg13g2_decap_8 FILLER_133_82 ();
 sg13g2_decap_8 FILLER_133_89 ();
 sg13g2_decap_4 FILLER_133_96 ();
 sg13g2_fill_1 FILLER_133_100 ();
 sg13g2_decap_8 FILLER_133_118 ();
 sg13g2_decap_8 FILLER_133_125 ();
 sg13g2_decap_8 FILLER_133_132 ();
 sg13g2_decap_8 FILLER_133_139 ();
 sg13g2_decap_8 FILLER_133_146 ();
 sg13g2_decap_8 FILLER_133_153 ();
 sg13g2_decap_8 FILLER_133_160 ();
 sg13g2_decap_4 FILLER_133_177 ();
 sg13g2_fill_1 FILLER_133_181 ();
 sg13g2_decap_8 FILLER_133_203 ();
 sg13g2_decap_8 FILLER_133_210 ();
 sg13g2_fill_1 FILLER_133_217 ();
 sg13g2_fill_2 FILLER_133_230 ();
 sg13g2_fill_1 FILLER_133_232 ();
 sg13g2_decap_8 FILLER_133_255 ();
 sg13g2_decap_8 FILLER_133_262 ();
 sg13g2_decap_4 FILLER_133_269 ();
 sg13g2_fill_2 FILLER_133_273 ();
 sg13g2_decap_8 FILLER_133_298 ();
 sg13g2_decap_8 FILLER_133_305 ();
 sg13g2_decap_8 FILLER_133_312 ();
 sg13g2_decap_8 FILLER_133_319 ();
 sg13g2_decap_8 FILLER_133_326 ();
 sg13g2_decap_8 FILLER_133_333 ();
 sg13g2_decap_8 FILLER_133_340 ();
 sg13g2_decap_8 FILLER_133_347 ();
 sg13g2_decap_8 FILLER_133_354 ();
 sg13g2_decap_8 FILLER_133_361 ();
 sg13g2_fill_2 FILLER_133_368 ();
 sg13g2_fill_1 FILLER_133_370 ();
 sg13g2_decap_8 FILLER_133_381 ();
 sg13g2_decap_8 FILLER_133_388 ();
 sg13g2_decap_8 FILLER_133_395 ();
 sg13g2_decap_4 FILLER_133_402 ();
 sg13g2_fill_2 FILLER_133_406 ();
 sg13g2_decap_4 FILLER_133_417 ();
 sg13g2_fill_1 FILLER_133_421 ();
 sg13g2_decap_8 FILLER_133_438 ();
 sg13g2_decap_8 FILLER_133_445 ();
 sg13g2_decap_8 FILLER_133_452 ();
 sg13g2_fill_2 FILLER_133_459 ();
 sg13g2_decap_8 FILLER_133_470 ();
 sg13g2_fill_1 FILLER_133_477 ();
 sg13g2_decap_8 FILLER_133_482 ();
 sg13g2_decap_8 FILLER_133_489 ();
 sg13g2_decap_8 FILLER_133_496 ();
 sg13g2_fill_2 FILLER_133_503 ();
 sg13g2_fill_1 FILLER_133_505 ();
 sg13g2_decap_8 FILLER_133_515 ();
 sg13g2_decap_8 FILLER_133_522 ();
 sg13g2_decap_8 FILLER_133_529 ();
 sg13g2_decap_4 FILLER_133_536 ();
 sg13g2_fill_2 FILLER_133_540 ();
 sg13g2_decap_8 FILLER_133_550 ();
 sg13g2_decap_8 FILLER_133_557 ();
 sg13g2_fill_1 FILLER_133_564 ();
 sg13g2_decap_8 FILLER_133_573 ();
 sg13g2_decap_8 FILLER_133_580 ();
 sg13g2_fill_1 FILLER_133_587 ();
 sg13g2_fill_2 FILLER_133_596 ();
 sg13g2_decap_4 FILLER_133_606 ();
 sg13g2_fill_2 FILLER_133_610 ();
 sg13g2_decap_8 FILLER_133_625 ();
 sg13g2_fill_2 FILLER_133_632 ();
 sg13g2_decap_8 FILLER_133_646 ();
 sg13g2_decap_8 FILLER_133_653 ();
 sg13g2_decap_8 FILLER_133_660 ();
 sg13g2_decap_8 FILLER_133_667 ();
 sg13g2_decap_8 FILLER_133_674 ();
 sg13g2_decap_8 FILLER_133_681 ();
 sg13g2_decap_8 FILLER_133_688 ();
 sg13g2_fill_2 FILLER_133_695 ();
 sg13g2_decap_8 FILLER_133_710 ();
 sg13g2_decap_8 FILLER_133_717 ();
 sg13g2_decap_8 FILLER_133_724 ();
 sg13g2_decap_8 FILLER_133_731 ();
 sg13g2_decap_8 FILLER_133_738 ();
 sg13g2_decap_8 FILLER_133_745 ();
 sg13g2_decap_8 FILLER_133_752 ();
 sg13g2_decap_8 FILLER_133_772 ();
 sg13g2_decap_8 FILLER_133_779 ();
 sg13g2_decap_8 FILLER_133_786 ();
 sg13g2_decap_8 FILLER_133_793 ();
 sg13g2_decap_4 FILLER_133_800 ();
 sg13g2_fill_1 FILLER_133_804 ();
 sg13g2_decap_8 FILLER_133_809 ();
 sg13g2_decap_8 FILLER_133_816 ();
 sg13g2_decap_8 FILLER_133_823 ();
 sg13g2_fill_1 FILLER_133_830 ();
 sg13g2_decap_4 FILLER_133_837 ();
 sg13g2_fill_1 FILLER_133_841 ();
 sg13g2_decap_8 FILLER_133_850 ();
 sg13g2_decap_8 FILLER_133_857 ();
 sg13g2_decap_8 FILLER_133_864 ();
 sg13g2_decap_8 FILLER_133_871 ();
 sg13g2_decap_8 FILLER_133_878 ();
 sg13g2_decap_8 FILLER_133_885 ();
 sg13g2_decap_8 FILLER_133_892 ();
 sg13g2_fill_1 FILLER_133_899 ();
 sg13g2_decap_8 FILLER_133_905 ();
 sg13g2_decap_8 FILLER_133_912 ();
 sg13g2_decap_8 FILLER_133_919 ();
 sg13g2_decap_8 FILLER_133_926 ();
 sg13g2_decap_4 FILLER_133_933 ();
 sg13g2_decap_8 FILLER_133_963 ();
 sg13g2_decap_8 FILLER_133_970 ();
 sg13g2_decap_8 FILLER_133_977 ();
 sg13g2_decap_8 FILLER_133_984 ();
 sg13g2_decap_8 FILLER_133_991 ();
 sg13g2_fill_2 FILLER_133_1037 ();
 sg13g2_decap_8 FILLER_133_1044 ();
 sg13g2_decap_8 FILLER_133_1051 ();
 sg13g2_decap_8 FILLER_133_1058 ();
 sg13g2_fill_1 FILLER_133_1065 ();
 sg13g2_decap_4 FILLER_133_1070 ();
 sg13g2_fill_1 FILLER_133_1074 ();
 sg13g2_fill_1 FILLER_133_1083 ();
 sg13g2_decap_8 FILLER_133_1101 ();
 sg13g2_fill_2 FILLER_133_1108 ();
 sg13g2_fill_1 FILLER_133_1110 ();
 sg13g2_decap_8 FILLER_133_1115 ();
 sg13g2_decap_8 FILLER_133_1122 ();
 sg13g2_decap_8 FILLER_133_1129 ();
 sg13g2_decap_8 FILLER_133_1136 ();
 sg13g2_decap_8 FILLER_133_1143 ();
 sg13g2_decap_8 FILLER_133_1150 ();
 sg13g2_decap_8 FILLER_133_1157 ();
 sg13g2_decap_4 FILLER_133_1164 ();
 sg13g2_fill_2 FILLER_133_1168 ();
 sg13g2_decap_8 FILLER_133_1173 ();
 sg13g2_decap_8 FILLER_133_1180 ();
 sg13g2_fill_2 FILLER_133_1187 ();
 sg13g2_fill_1 FILLER_133_1189 ();
 sg13g2_fill_1 FILLER_133_1199 ();
 sg13g2_fill_1 FILLER_133_1214 ();
 sg13g2_decap_8 FILLER_133_1228 ();
 sg13g2_fill_2 FILLER_133_1235 ();
 sg13g2_decap_8 FILLER_133_1257 ();
 sg13g2_decap_8 FILLER_133_1264 ();
 sg13g2_decap_8 FILLER_133_1271 ();
 sg13g2_decap_8 FILLER_133_1278 ();
 sg13g2_decap_8 FILLER_133_1285 ();
 sg13g2_decap_8 FILLER_133_1292 ();
 sg13g2_decap_8 FILLER_133_1299 ();
 sg13g2_decap_8 FILLER_133_1311 ();
 sg13g2_decap_8 FILLER_133_1318 ();
 sg13g2_decap_8 FILLER_133_1325 ();
 sg13g2_fill_1 FILLER_133_1344 ();
 sg13g2_decap_8 FILLER_133_1383 ();
 sg13g2_fill_1 FILLER_133_1390 ();
 sg13g2_decap_8 FILLER_133_1417 ();
 sg13g2_fill_1 FILLER_133_1424 ();
 sg13g2_decap_8 FILLER_133_1433 ();
 sg13g2_decap_4 FILLER_133_1440 ();
 sg13g2_fill_1 FILLER_133_1457 ();
 sg13g2_decap_8 FILLER_133_1466 ();
 sg13g2_decap_8 FILLER_133_1473 ();
 sg13g2_decap_8 FILLER_133_1480 ();
 sg13g2_decap_8 FILLER_133_1487 ();
 sg13g2_decap_8 FILLER_133_1494 ();
 sg13g2_decap_8 FILLER_133_1516 ();
 sg13g2_decap_8 FILLER_133_1523 ();
 sg13g2_decap_8 FILLER_133_1530 ();
 sg13g2_decap_8 FILLER_133_1537 ();
 sg13g2_decap_8 FILLER_133_1544 ();
 sg13g2_decap_4 FILLER_133_1551 ();
 sg13g2_fill_1 FILLER_133_1555 ();
 sg13g2_decap_8 FILLER_133_1564 ();
 sg13g2_decap_8 FILLER_133_1571 ();
 sg13g2_decap_8 FILLER_133_1578 ();
 sg13g2_decap_8 FILLER_133_1585 ();
 sg13g2_decap_4 FILLER_133_1592 ();
 sg13g2_fill_2 FILLER_133_1596 ();
 sg13g2_decap_8 FILLER_133_1629 ();
 sg13g2_decap_8 FILLER_133_1636 ();
 sg13g2_decap_8 FILLER_133_1643 ();
 sg13g2_decap_8 FILLER_133_1650 ();
 sg13g2_decap_8 FILLER_133_1665 ();
 sg13g2_decap_8 FILLER_133_1685 ();
 sg13g2_decap_8 FILLER_133_1692 ();
 sg13g2_decap_8 FILLER_133_1699 ();
 sg13g2_decap_4 FILLER_133_1706 ();
 sg13g2_fill_1 FILLER_133_1710 ();
 sg13g2_decap_8 FILLER_133_1727 ();
 sg13g2_decap_8 FILLER_133_1749 ();
 sg13g2_decap_8 FILLER_133_1756 ();
 sg13g2_decap_4 FILLER_133_1763 ();
 sg13g2_fill_1 FILLER_133_1767 ();
 sg13g2_decap_8 FILLER_134_0 ();
 sg13g2_decap_8 FILLER_134_7 ();
 sg13g2_decap_4 FILLER_134_14 ();
 sg13g2_fill_1 FILLER_134_18 ();
 sg13g2_decap_8 FILLER_134_33 ();
 sg13g2_decap_8 FILLER_134_40 ();
 sg13g2_fill_2 FILLER_134_47 ();
 sg13g2_decap_8 FILLER_134_77 ();
 sg13g2_decap_8 FILLER_134_84 ();
 sg13g2_decap_8 FILLER_134_91 ();
 sg13g2_fill_1 FILLER_134_106 ();
 sg13g2_decap_8 FILLER_134_124 ();
 sg13g2_decap_8 FILLER_134_131 ();
 sg13g2_decap_8 FILLER_134_138 ();
 sg13g2_decap_8 FILLER_134_145 ();
 sg13g2_decap_8 FILLER_134_152 ();
 sg13g2_decap_4 FILLER_134_159 ();
 sg13g2_fill_2 FILLER_134_163 ();
 sg13g2_decap_4 FILLER_134_173 ();
 sg13g2_fill_1 FILLER_134_177 ();
 sg13g2_decap_8 FILLER_134_196 ();
 sg13g2_decap_8 FILLER_134_207 ();
 sg13g2_decap_8 FILLER_134_214 ();
 sg13g2_decap_8 FILLER_134_221 ();
 sg13g2_decap_8 FILLER_134_228 ();
 sg13g2_fill_1 FILLER_134_235 ();
 sg13g2_decap_8 FILLER_134_252 ();
 sg13g2_decap_8 FILLER_134_259 ();
 sg13g2_decap_8 FILLER_134_266 ();
 sg13g2_decap_8 FILLER_134_273 ();
 sg13g2_decap_8 FILLER_134_280 ();
 sg13g2_decap_8 FILLER_134_295 ();
 sg13g2_decap_8 FILLER_134_302 ();
 sg13g2_decap_8 FILLER_134_309 ();
 sg13g2_fill_2 FILLER_134_316 ();
 sg13g2_fill_1 FILLER_134_318 ();
 sg13g2_decap_8 FILLER_134_345 ();
 sg13g2_fill_2 FILLER_134_352 ();
 sg13g2_decap_4 FILLER_134_362 ();
 sg13g2_fill_2 FILLER_134_371 ();
 sg13g2_decap_8 FILLER_134_381 ();
 sg13g2_decap_4 FILLER_134_388 ();
 sg13g2_fill_2 FILLER_134_406 ();
 sg13g2_decap_8 FILLER_134_422 ();
 sg13g2_decap_8 FILLER_134_429 ();
 sg13g2_decap_8 FILLER_134_436 ();
 sg13g2_decap_8 FILLER_134_443 ();
 sg13g2_decap_8 FILLER_134_450 ();
 sg13g2_decap_8 FILLER_134_457 ();
 sg13g2_decap_4 FILLER_134_464 ();
 sg13g2_decap_8 FILLER_134_472 ();
 sg13g2_decap_8 FILLER_134_479 ();
 sg13g2_fill_2 FILLER_134_486 ();
 sg13g2_decap_8 FILLER_134_496 ();
 sg13g2_decap_4 FILLER_134_503 ();
 sg13g2_fill_2 FILLER_134_507 ();
 sg13g2_decap_8 FILLER_134_512 ();
 sg13g2_decap_8 FILLER_134_519 ();
 sg13g2_fill_1 FILLER_134_526 ();
 sg13g2_decap_4 FILLER_134_538 ();
 sg13g2_fill_1 FILLER_134_542 ();
 sg13g2_decap_8 FILLER_134_562 ();
 sg13g2_decap_8 FILLER_134_569 ();
 sg13g2_decap_8 FILLER_134_576 ();
 sg13g2_decap_8 FILLER_134_583 ();
 sg13g2_decap_4 FILLER_134_590 ();
 sg13g2_fill_2 FILLER_134_594 ();
 sg13g2_decap_8 FILLER_134_600 ();
 sg13g2_decap_8 FILLER_134_607 ();
 sg13g2_decap_8 FILLER_134_614 ();
 sg13g2_decap_8 FILLER_134_621 ();
 sg13g2_fill_1 FILLER_134_654 ();
 sg13g2_fill_1 FILLER_134_663 ();
 sg13g2_decap_8 FILLER_134_671 ();
 sg13g2_decap_8 FILLER_134_678 ();
 sg13g2_decap_8 FILLER_134_685 ();
 sg13g2_decap_8 FILLER_134_692 ();
 sg13g2_fill_1 FILLER_134_699 ();
 sg13g2_decap_8 FILLER_134_713 ();
 sg13g2_decap_8 FILLER_134_720 ();
 sg13g2_fill_2 FILLER_134_727 ();
 sg13g2_decap_8 FILLER_134_732 ();
 sg13g2_decap_8 FILLER_134_743 ();
 sg13g2_decap_8 FILLER_134_750 ();
 sg13g2_decap_8 FILLER_134_757 ();
 sg13g2_decap_8 FILLER_134_764 ();
 sg13g2_decap_8 FILLER_134_771 ();
 sg13g2_decap_8 FILLER_134_778 ();
 sg13g2_decap_8 FILLER_134_785 ();
 sg13g2_decap_8 FILLER_134_792 ();
 sg13g2_decap_8 FILLER_134_799 ();
 sg13g2_decap_8 FILLER_134_806 ();
 sg13g2_decap_8 FILLER_134_813 ();
 sg13g2_decap_8 FILLER_134_820 ();
 sg13g2_fill_2 FILLER_134_827 ();
 sg13g2_decap_8 FILLER_134_837 ();
 sg13g2_decap_8 FILLER_134_848 ();
 sg13g2_decap_4 FILLER_134_855 ();
 sg13g2_decap_8 FILLER_134_864 ();
 sg13g2_decap_8 FILLER_134_871 ();
 sg13g2_decap_8 FILLER_134_878 ();
 sg13g2_decap_8 FILLER_134_885 ();
 sg13g2_decap_4 FILLER_134_892 ();
 sg13g2_fill_2 FILLER_134_896 ();
 sg13g2_decap_8 FILLER_134_902 ();
 sg13g2_decap_8 FILLER_134_909 ();
 sg13g2_decap_8 FILLER_134_916 ();
 sg13g2_decap_8 FILLER_134_923 ();
 sg13g2_decap_8 FILLER_134_930 ();
 sg13g2_decap_8 FILLER_134_937 ();
 sg13g2_decap_4 FILLER_134_944 ();
 sg13g2_decap_8 FILLER_134_958 ();
 sg13g2_decap_8 FILLER_134_965 ();
 sg13g2_fill_2 FILLER_134_972 ();
 sg13g2_fill_1 FILLER_134_974 ();
 sg13g2_fill_2 FILLER_134_993 ();
 sg13g2_decap_8 FILLER_134_1016 ();
 sg13g2_decap_8 FILLER_134_1023 ();
 sg13g2_decap_4 FILLER_134_1030 ();
 sg13g2_fill_1 FILLER_134_1034 ();
 sg13g2_decap_8 FILLER_134_1048 ();
 sg13g2_decap_4 FILLER_134_1055 ();
 sg13g2_decap_8 FILLER_134_1067 ();
 sg13g2_decap_4 FILLER_134_1074 ();
 sg13g2_decap_8 FILLER_134_1107 ();
 sg13g2_decap_8 FILLER_134_1114 ();
 sg13g2_decap_8 FILLER_134_1121 ();
 sg13g2_decap_8 FILLER_134_1128 ();
 sg13g2_decap_8 FILLER_134_1135 ();
 sg13g2_fill_2 FILLER_134_1142 ();
 sg13g2_decap_8 FILLER_134_1153 ();
 sg13g2_decap_8 FILLER_134_1160 ();
 sg13g2_fill_2 FILLER_134_1167 ();
 sg13g2_fill_1 FILLER_134_1169 ();
 sg13g2_decap_8 FILLER_134_1173 ();
 sg13g2_decap_8 FILLER_134_1180 ();
 sg13g2_decap_8 FILLER_134_1187 ();
 sg13g2_decap_4 FILLER_134_1194 ();
 sg13g2_fill_1 FILLER_134_1198 ();
 sg13g2_decap_8 FILLER_134_1215 ();
 sg13g2_decap_8 FILLER_134_1222 ();
 sg13g2_fill_1 FILLER_134_1240 ();
 sg13g2_decap_8 FILLER_134_1265 ();
 sg13g2_fill_2 FILLER_134_1272 ();
 sg13g2_fill_1 FILLER_134_1274 ();
 sg13g2_decap_8 FILLER_134_1281 ();
 sg13g2_fill_1 FILLER_134_1288 ();
 sg13g2_decap_8 FILLER_134_1297 ();
 sg13g2_decap_8 FILLER_134_1304 ();
 sg13g2_decap_8 FILLER_134_1311 ();
 sg13g2_decap_8 FILLER_134_1318 ();
 sg13g2_decap_8 FILLER_134_1325 ();
 sg13g2_decap_8 FILLER_134_1332 ();
 sg13g2_decap_4 FILLER_134_1339 ();
 sg13g2_fill_1 FILLER_134_1343 ();
 sg13g2_decap_8 FILLER_134_1368 ();
 sg13g2_decap_8 FILLER_134_1375 ();
 sg13g2_decap_8 FILLER_134_1382 ();
 sg13g2_decap_8 FILLER_134_1389 ();
 sg13g2_decap_8 FILLER_134_1396 ();
 sg13g2_decap_8 FILLER_134_1403 ();
 sg13g2_decap_8 FILLER_134_1410 ();
 sg13g2_decap_8 FILLER_134_1417 ();
 sg13g2_decap_8 FILLER_134_1424 ();
 sg13g2_decap_8 FILLER_134_1431 ();
 sg13g2_decap_8 FILLER_134_1438 ();
 sg13g2_decap_8 FILLER_134_1445 ();
 sg13g2_fill_1 FILLER_134_1452 ();
 sg13g2_decap_8 FILLER_134_1458 ();
 sg13g2_decap_8 FILLER_134_1465 ();
 sg13g2_decap_8 FILLER_134_1472 ();
 sg13g2_decap_8 FILLER_134_1479 ();
 sg13g2_decap_8 FILLER_134_1486 ();
 sg13g2_decap_8 FILLER_134_1493 ();
 sg13g2_decap_4 FILLER_134_1507 ();
 sg13g2_decap_8 FILLER_134_1527 ();
 sg13g2_decap_8 FILLER_134_1534 ();
 sg13g2_decap_8 FILLER_134_1541 ();
 sg13g2_decap_4 FILLER_134_1548 ();
 sg13g2_fill_2 FILLER_134_1552 ();
 sg13g2_decap_8 FILLER_134_1557 ();
 sg13g2_decap_8 FILLER_134_1564 ();
 sg13g2_decap_8 FILLER_134_1571 ();
 sg13g2_decap_8 FILLER_134_1578 ();
 sg13g2_decap_8 FILLER_134_1585 ();
 sg13g2_fill_2 FILLER_134_1602 ();
 sg13g2_fill_1 FILLER_134_1604 ();
 sg13g2_fill_1 FILLER_134_1618 ();
 sg13g2_decap_8 FILLER_134_1628 ();
 sg13g2_decap_8 FILLER_134_1635 ();
 sg13g2_decap_8 FILLER_134_1642 ();
 sg13g2_decap_8 FILLER_134_1649 ();
 sg13g2_decap_8 FILLER_134_1656 ();
 sg13g2_decap_8 FILLER_134_1663 ();
 sg13g2_fill_2 FILLER_134_1670 ();
 sg13g2_decap_4 FILLER_134_1678 ();
 sg13g2_decap_8 FILLER_134_1690 ();
 sg13g2_decap_4 FILLER_134_1697 ();
 sg13g2_fill_1 FILLER_134_1701 ();
 sg13g2_decap_8 FILLER_134_1724 ();
 sg13g2_decap_8 FILLER_134_1731 ();
 sg13g2_decap_8 FILLER_134_1738 ();
 sg13g2_decap_8 FILLER_134_1745 ();
 sg13g2_decap_8 FILLER_134_1752 ();
 sg13g2_decap_8 FILLER_134_1759 ();
 sg13g2_fill_2 FILLER_134_1766 ();
 sg13g2_decap_8 FILLER_135_0 ();
 sg13g2_decap_8 FILLER_135_7 ();
 sg13g2_decap_8 FILLER_135_14 ();
 sg13g2_decap_8 FILLER_135_21 ();
 sg13g2_decap_8 FILLER_135_28 ();
 sg13g2_fill_2 FILLER_135_35 ();
 sg13g2_fill_1 FILLER_135_37 ();
 sg13g2_fill_1 FILLER_135_63 ();
 sg13g2_decap_8 FILLER_135_69 ();
 sg13g2_decap_8 FILLER_135_76 ();
 sg13g2_decap_8 FILLER_135_83 ();
 sg13g2_decap_8 FILLER_135_90 ();
 sg13g2_decap_4 FILLER_135_97 ();
 sg13g2_decap_8 FILLER_135_127 ();
 sg13g2_decap_8 FILLER_135_134 ();
 sg13g2_decap_8 FILLER_135_141 ();
 sg13g2_decap_8 FILLER_135_148 ();
 sg13g2_decap_8 FILLER_135_155 ();
 sg13g2_decap_8 FILLER_135_162 ();
 sg13g2_decap_8 FILLER_135_169 ();
 sg13g2_decap_8 FILLER_135_176 ();
 sg13g2_decap_4 FILLER_135_183 ();
 sg13g2_decap_8 FILLER_135_195 ();
 sg13g2_decap_8 FILLER_135_202 ();
 sg13g2_decap_8 FILLER_135_209 ();
 sg13g2_decap_8 FILLER_135_216 ();
 sg13g2_decap_8 FILLER_135_223 ();
 sg13g2_decap_8 FILLER_135_230 ();
 sg13g2_decap_8 FILLER_135_237 ();
 sg13g2_decap_8 FILLER_135_244 ();
 sg13g2_decap_8 FILLER_135_251 ();
 sg13g2_decap_8 FILLER_135_258 ();
 sg13g2_decap_4 FILLER_135_265 ();
 sg13g2_fill_1 FILLER_135_269 ();
 sg13g2_decap_8 FILLER_135_273 ();
 sg13g2_decap_8 FILLER_135_280 ();
 sg13g2_decap_8 FILLER_135_287 ();
 sg13g2_decap_8 FILLER_135_294 ();
 sg13g2_decap_8 FILLER_135_301 ();
 sg13g2_decap_8 FILLER_135_308 ();
 sg13g2_decap_8 FILLER_135_315 ();
 sg13g2_decap_4 FILLER_135_322 ();
 sg13g2_fill_2 FILLER_135_326 ();
 sg13g2_decap_8 FILLER_135_368 ();
 sg13g2_decap_8 FILLER_135_375 ();
 sg13g2_decap_8 FILLER_135_382 ();
 sg13g2_decap_8 FILLER_135_389 ();
 sg13g2_decap_8 FILLER_135_396 ();
 sg13g2_decap_4 FILLER_135_411 ();
 sg13g2_fill_2 FILLER_135_415 ();
 sg13g2_decap_8 FILLER_135_427 ();
 sg13g2_decap_8 FILLER_135_434 ();
 sg13g2_decap_8 FILLER_135_441 ();
 sg13g2_decap_8 FILLER_135_448 ();
 sg13g2_fill_2 FILLER_135_455 ();
 sg13g2_decap_8 FILLER_135_465 ();
 sg13g2_decap_4 FILLER_135_472 ();
 sg13g2_decap_8 FILLER_135_480 ();
 sg13g2_decap_8 FILLER_135_487 ();
 sg13g2_decap_8 FILLER_135_494 ();
 sg13g2_fill_2 FILLER_135_501 ();
 sg13g2_decap_8 FILLER_135_513 ();
 sg13g2_decap_8 FILLER_135_520 ();
 sg13g2_decap_8 FILLER_135_527 ();
 sg13g2_fill_2 FILLER_135_534 ();
 sg13g2_decap_8 FILLER_135_540 ();
 sg13g2_decap_8 FILLER_135_547 ();
 sg13g2_fill_2 FILLER_135_554 ();
 sg13g2_fill_1 FILLER_135_556 ();
 sg13g2_decap_8 FILLER_135_562 ();
 sg13g2_decap_8 FILLER_135_569 ();
 sg13g2_fill_2 FILLER_135_576 ();
 sg13g2_fill_1 FILLER_135_578 ();
 sg13g2_decap_8 FILLER_135_587 ();
 sg13g2_fill_1 FILLER_135_601 ();
 sg13g2_decap_8 FILLER_135_605 ();
 sg13g2_decap_8 FILLER_135_612 ();
 sg13g2_decap_8 FILLER_135_619 ();
 sg13g2_decap_8 FILLER_135_626 ();
 sg13g2_decap_8 FILLER_135_669 ();
 sg13g2_decap_8 FILLER_135_676 ();
 sg13g2_decap_8 FILLER_135_683 ();
 sg13g2_decap_8 FILLER_135_690 ();
 sg13g2_decap_8 FILLER_135_697 ();
 sg13g2_decap_8 FILLER_135_704 ();
 sg13g2_decap_8 FILLER_135_711 ();
 sg13g2_decap_4 FILLER_135_718 ();
 sg13g2_fill_1 FILLER_135_722 ();
 sg13g2_fill_2 FILLER_135_739 ();
 sg13g2_decap_8 FILLER_135_746 ();
 sg13g2_decap_8 FILLER_135_753 ();
 sg13g2_decap_8 FILLER_135_760 ();
 sg13g2_decap_8 FILLER_135_767 ();
 sg13g2_decap_8 FILLER_135_774 ();
 sg13g2_fill_2 FILLER_135_781 ();
 sg13g2_fill_1 FILLER_135_783 ();
 sg13g2_decap_8 FILLER_135_802 ();
 sg13g2_decap_8 FILLER_135_809 ();
 sg13g2_decap_8 FILLER_135_816 ();
 sg13g2_decap_8 FILLER_135_823 ();
 sg13g2_decap_8 FILLER_135_830 ();
 sg13g2_decap_8 FILLER_135_837 ();
 sg13g2_decap_4 FILLER_135_844 ();
 sg13g2_fill_1 FILLER_135_848 ();
 sg13g2_fill_2 FILLER_135_862 ();
 sg13g2_fill_2 FILLER_135_873 ();
 sg13g2_fill_1 FILLER_135_875 ();
 sg13g2_decap_8 FILLER_135_879 ();
 sg13g2_decap_4 FILLER_135_886 ();
 sg13g2_fill_2 FILLER_135_890 ();
 sg13g2_decap_8 FILLER_135_917 ();
 sg13g2_decap_8 FILLER_135_924 ();
 sg13g2_decap_4 FILLER_135_931 ();
 sg13g2_fill_1 FILLER_135_935 ();
 sg13g2_fill_1 FILLER_135_948 ();
 sg13g2_decap_8 FILLER_135_961 ();
 sg13g2_decap_8 FILLER_135_968 ();
 sg13g2_fill_2 FILLER_135_975 ();
 sg13g2_fill_1 FILLER_135_977 ();
 sg13g2_fill_2 FILLER_135_983 ();
 sg13g2_decap_8 FILLER_135_989 ();
 sg13g2_decap_4 FILLER_135_996 ();
 sg13g2_decap_8 FILLER_135_1008 ();
 sg13g2_decap_8 FILLER_135_1015 ();
 sg13g2_decap_8 FILLER_135_1022 ();
 sg13g2_fill_1 FILLER_135_1029 ();
 sg13g2_decap_8 FILLER_135_1042 ();
 sg13g2_decap_8 FILLER_135_1049 ();
 sg13g2_decap_8 FILLER_135_1056 ();
 sg13g2_decap_8 FILLER_135_1063 ();
 sg13g2_decap_4 FILLER_135_1070 ();
 sg13g2_decap_4 FILLER_135_1082 ();
 sg13g2_fill_1 FILLER_135_1086 ();
 sg13g2_decap_8 FILLER_135_1099 ();
 sg13g2_decap_8 FILLER_135_1106 ();
 sg13g2_decap_8 FILLER_135_1113 ();
 sg13g2_decap_8 FILLER_135_1120 ();
 sg13g2_fill_1 FILLER_135_1127 ();
 sg13g2_decap_8 FILLER_135_1136 ();
 sg13g2_decap_8 FILLER_135_1143 ();
 sg13g2_decap_8 FILLER_135_1150 ();
 sg13g2_decap_8 FILLER_135_1157 ();
 sg13g2_decap_4 FILLER_135_1164 ();
 sg13g2_fill_1 FILLER_135_1168 ();
 sg13g2_decap_8 FILLER_135_1174 ();
 sg13g2_decap_8 FILLER_135_1181 ();
 sg13g2_decap_8 FILLER_135_1188 ();
 sg13g2_fill_2 FILLER_135_1195 ();
 sg13g2_fill_1 FILLER_135_1197 ();
 sg13g2_decap_8 FILLER_135_1205 ();
 sg13g2_decap_8 FILLER_135_1212 ();
 sg13g2_decap_8 FILLER_135_1219 ();
 sg13g2_decap_4 FILLER_135_1226 ();
 sg13g2_fill_2 FILLER_135_1230 ();
 sg13g2_decap_8 FILLER_135_1254 ();
 sg13g2_decap_8 FILLER_135_1261 ();
 sg13g2_decap_4 FILLER_135_1268 ();
 sg13g2_fill_2 FILLER_135_1272 ();
 sg13g2_decap_8 FILLER_135_1295 ();
 sg13g2_decap_8 FILLER_135_1302 ();
 sg13g2_decap_8 FILLER_135_1309 ();
 sg13g2_decap_8 FILLER_135_1316 ();
 sg13g2_decap_8 FILLER_135_1323 ();
 sg13g2_decap_8 FILLER_135_1330 ();
 sg13g2_decap_8 FILLER_135_1337 ();
 sg13g2_decap_8 FILLER_135_1344 ();
 sg13g2_decap_8 FILLER_135_1351 ();
 sg13g2_decap_8 FILLER_135_1358 ();
 sg13g2_decap_8 FILLER_135_1365 ();
 sg13g2_decap_8 FILLER_135_1372 ();
 sg13g2_decap_8 FILLER_135_1379 ();
 sg13g2_decap_8 FILLER_135_1386 ();
 sg13g2_decap_8 FILLER_135_1393 ();
 sg13g2_decap_8 FILLER_135_1400 ();
 sg13g2_decap_8 FILLER_135_1407 ();
 sg13g2_decap_8 FILLER_135_1414 ();
 sg13g2_decap_8 FILLER_135_1421 ();
 sg13g2_decap_8 FILLER_135_1428 ();
 sg13g2_decap_8 FILLER_135_1435 ();
 sg13g2_fill_2 FILLER_135_1442 ();
 sg13g2_fill_2 FILLER_135_1448 ();
 sg13g2_decap_4 FILLER_135_1454 ();
 sg13g2_fill_2 FILLER_135_1458 ();
 sg13g2_decap_8 FILLER_135_1464 ();
 sg13g2_decap_8 FILLER_135_1471 ();
 sg13g2_decap_8 FILLER_135_1478 ();
 sg13g2_decap_8 FILLER_135_1485 ();
 sg13g2_decap_8 FILLER_135_1492 ();
 sg13g2_decap_8 FILLER_135_1499 ();
 sg13g2_decap_8 FILLER_135_1506 ();
 sg13g2_decap_8 FILLER_135_1513 ();
 sg13g2_decap_8 FILLER_135_1520 ();
 sg13g2_decap_8 FILLER_135_1527 ();
 sg13g2_decap_8 FILLER_135_1534 ();
 sg13g2_fill_2 FILLER_135_1541 ();
 sg13g2_decap_8 FILLER_135_1568 ();
 sg13g2_decap_8 FILLER_135_1575 ();
 sg13g2_decap_8 FILLER_135_1582 ();
 sg13g2_decap_8 FILLER_135_1589 ();
 sg13g2_decap_8 FILLER_135_1596 ();
 sg13g2_decap_8 FILLER_135_1603 ();
 sg13g2_decap_8 FILLER_135_1610 ();
 sg13g2_decap_8 FILLER_135_1617 ();
 sg13g2_decap_8 FILLER_135_1624 ();
 sg13g2_decap_8 FILLER_135_1631 ();
 sg13g2_decap_8 FILLER_135_1638 ();
 sg13g2_decap_8 FILLER_135_1645 ();
 sg13g2_decap_8 FILLER_135_1652 ();
 sg13g2_decap_8 FILLER_135_1659 ();
 sg13g2_decap_8 FILLER_135_1666 ();
 sg13g2_fill_2 FILLER_135_1673 ();
 sg13g2_fill_2 FILLER_135_1688 ();
 sg13g2_decap_8 FILLER_135_1707 ();
 sg13g2_decap_8 FILLER_135_1714 ();
 sg13g2_decap_8 FILLER_135_1721 ();
 sg13g2_fill_2 FILLER_135_1728 ();
 sg13g2_decap_8 FILLER_135_1738 ();
 sg13g2_decap_8 FILLER_135_1745 ();
 sg13g2_decap_8 FILLER_135_1752 ();
 sg13g2_decap_8 FILLER_135_1759 ();
 sg13g2_fill_2 FILLER_135_1766 ();
 sg13g2_decap_8 FILLER_136_0 ();
 sg13g2_decap_8 FILLER_136_7 ();
 sg13g2_decap_8 FILLER_136_14 ();
 sg13g2_decap_4 FILLER_136_21 ();
 sg13g2_fill_1 FILLER_136_25 ();
 sg13g2_decap_4 FILLER_136_45 ();
 sg13g2_fill_1 FILLER_136_49 ();
 sg13g2_decap_8 FILLER_136_63 ();
 sg13g2_decap_8 FILLER_136_70 ();
 sg13g2_decap_8 FILLER_136_77 ();
 sg13g2_decap_8 FILLER_136_84 ();
 sg13g2_decap_8 FILLER_136_91 ();
 sg13g2_decap_8 FILLER_136_98 ();
 sg13g2_fill_2 FILLER_136_105 ();
 sg13g2_fill_1 FILLER_136_107 ();
 sg13g2_decap_8 FILLER_136_121 ();
 sg13g2_decap_8 FILLER_136_128 ();
 sg13g2_decap_8 FILLER_136_135 ();
 sg13g2_decap_4 FILLER_136_146 ();
 sg13g2_fill_2 FILLER_136_150 ();
 sg13g2_decap_8 FILLER_136_174 ();
 sg13g2_decap_4 FILLER_136_181 ();
 sg13g2_fill_1 FILLER_136_185 ();
 sg13g2_decap_8 FILLER_136_198 ();
 sg13g2_decap_8 FILLER_136_205 ();
 sg13g2_decap_8 FILLER_136_216 ();
 sg13g2_decap_8 FILLER_136_223 ();
 sg13g2_decap_8 FILLER_136_230 ();
 sg13g2_decap_8 FILLER_136_237 ();
 sg13g2_decap_8 FILLER_136_244 ();
 sg13g2_decap_8 FILLER_136_251 ();
 sg13g2_decap_4 FILLER_136_258 ();
 sg13g2_fill_1 FILLER_136_262 ();
 sg13g2_fill_2 FILLER_136_268 ();
 sg13g2_decap_8 FILLER_136_275 ();
 sg13g2_decap_8 FILLER_136_282 ();
 sg13g2_decap_8 FILLER_136_289 ();
 sg13g2_decap_4 FILLER_136_296 ();
 sg13g2_decap_8 FILLER_136_314 ();
 sg13g2_decap_8 FILLER_136_321 ();
 sg13g2_decap_8 FILLER_136_328 ();
 sg13g2_decap_4 FILLER_136_335 ();
 sg13g2_fill_2 FILLER_136_339 ();
 sg13g2_decap_8 FILLER_136_345 ();
 sg13g2_decap_8 FILLER_136_352 ();
 sg13g2_fill_1 FILLER_136_359 ();
 sg13g2_decap_8 FILLER_136_373 ();
 sg13g2_decap_8 FILLER_136_380 ();
 sg13g2_decap_8 FILLER_136_387 ();
 sg13g2_decap_8 FILLER_136_394 ();
 sg13g2_decap_8 FILLER_136_401 ();
 sg13g2_decap_8 FILLER_136_408 ();
 sg13g2_decap_8 FILLER_136_423 ();
 sg13g2_decap_4 FILLER_136_430 ();
 sg13g2_fill_2 FILLER_136_434 ();
 sg13g2_decap_8 FILLER_136_440 ();
 sg13g2_decap_8 FILLER_136_447 ();
 sg13g2_decap_4 FILLER_136_454 ();
 sg13g2_fill_2 FILLER_136_458 ();
 sg13g2_fill_2 FILLER_136_465 ();
 sg13g2_fill_1 FILLER_136_467 ();
 sg13g2_decap_8 FILLER_136_472 ();
 sg13g2_decap_8 FILLER_136_479 ();
 sg13g2_decap_4 FILLER_136_486 ();
 sg13g2_decap_8 FILLER_136_496 ();
 sg13g2_decap_8 FILLER_136_503 ();
 sg13g2_decap_8 FILLER_136_525 ();
 sg13g2_decap_8 FILLER_136_532 ();
 sg13g2_decap_8 FILLER_136_539 ();
 sg13g2_decap_8 FILLER_136_546 ();
 sg13g2_decap_8 FILLER_136_553 ();
 sg13g2_decap_8 FILLER_136_560 ();
 sg13g2_decap_4 FILLER_136_567 ();
 sg13g2_decap_8 FILLER_136_576 ();
 sg13g2_decap_8 FILLER_136_583 ();
 sg13g2_fill_1 FILLER_136_590 ();
 sg13g2_decap_8 FILLER_136_613 ();
 sg13g2_decap_8 FILLER_136_620 ();
 sg13g2_decap_8 FILLER_136_627 ();
 sg13g2_fill_2 FILLER_136_634 ();
 sg13g2_fill_1 FILLER_136_636 ();
 sg13g2_decap_8 FILLER_136_645 ();
 sg13g2_decap_8 FILLER_136_652 ();
 sg13g2_decap_8 FILLER_136_659 ();
 sg13g2_decap_8 FILLER_136_666 ();
 sg13g2_decap_8 FILLER_136_673 ();
 sg13g2_decap_8 FILLER_136_705 ();
 sg13g2_decap_4 FILLER_136_712 ();
 sg13g2_fill_1 FILLER_136_716 ();
 sg13g2_decap_8 FILLER_136_733 ();
 sg13g2_fill_1 FILLER_136_740 ();
 sg13g2_decap_4 FILLER_136_749 ();
 sg13g2_decap_8 FILLER_136_761 ();
 sg13g2_decap_8 FILLER_136_768 ();
 sg13g2_decap_8 FILLER_136_775 ();
 sg13g2_decap_8 FILLER_136_782 ();
 sg13g2_decap_4 FILLER_136_789 ();
 sg13g2_fill_1 FILLER_136_793 ();
 sg13g2_fill_2 FILLER_136_802 ();
 sg13g2_decap_8 FILLER_136_817 ();
 sg13g2_decap_8 FILLER_136_824 ();
 sg13g2_fill_2 FILLER_136_831 ();
 sg13g2_decap_4 FILLER_136_841 ();
 sg13g2_decap_8 FILLER_136_861 ();
 sg13g2_decap_8 FILLER_136_868 ();
 sg13g2_fill_1 FILLER_136_875 ();
 sg13g2_decap_8 FILLER_136_894 ();
 sg13g2_decap_8 FILLER_136_901 ();
 sg13g2_decap_8 FILLER_136_908 ();
 sg13g2_decap_8 FILLER_136_915 ();
 sg13g2_decap_8 FILLER_136_922 ();
 sg13g2_decap_8 FILLER_136_929 ();
 sg13g2_decap_8 FILLER_136_936 ();
 sg13g2_decap_8 FILLER_136_943 ();
 sg13g2_decap_8 FILLER_136_950 ();
 sg13g2_decap_8 FILLER_136_957 ();
 sg13g2_decap_8 FILLER_136_964 ();
 sg13g2_decap_8 FILLER_136_971 ();
 sg13g2_fill_2 FILLER_136_978 ();
 sg13g2_fill_1 FILLER_136_980 ();
 sg13g2_fill_1 FILLER_136_990 ();
 sg13g2_decap_8 FILLER_136_996 ();
 sg13g2_decap_8 FILLER_136_1003 ();
 sg13g2_decap_8 FILLER_136_1010 ();
 sg13g2_decap_8 FILLER_136_1017 ();
 sg13g2_decap_8 FILLER_136_1024 ();
 sg13g2_decap_8 FILLER_136_1031 ();
 sg13g2_decap_8 FILLER_136_1038 ();
 sg13g2_decap_8 FILLER_136_1045 ();
 sg13g2_decap_4 FILLER_136_1072 ();
 sg13g2_fill_1 FILLER_136_1076 ();
 sg13g2_decap_8 FILLER_136_1080 ();
 sg13g2_decap_8 FILLER_136_1087 ();
 sg13g2_decap_8 FILLER_136_1094 ();
 sg13g2_fill_1 FILLER_136_1101 ();
 sg13g2_decap_8 FILLER_136_1106 ();
 sg13g2_decap_8 FILLER_136_1113 ();
 sg13g2_decap_4 FILLER_136_1120 ();
 sg13g2_decap_8 FILLER_136_1128 ();
 sg13g2_decap_8 FILLER_136_1135 ();
 sg13g2_decap_8 FILLER_136_1142 ();
 sg13g2_decap_8 FILLER_136_1149 ();
 sg13g2_decap_8 FILLER_136_1180 ();
 sg13g2_decap_8 FILLER_136_1216 ();
 sg13g2_decap_8 FILLER_136_1223 ();
 sg13g2_decap_8 FILLER_136_1230 ();
 sg13g2_decap_4 FILLER_136_1237 ();
 sg13g2_decap_8 FILLER_136_1250 ();
 sg13g2_decap_8 FILLER_136_1257 ();
 sg13g2_decap_8 FILLER_136_1264 ();
 sg13g2_fill_2 FILLER_136_1285 ();
 sg13g2_decap_4 FILLER_136_1299 ();
 sg13g2_fill_2 FILLER_136_1303 ();
 sg13g2_decap_8 FILLER_136_1313 ();
 sg13g2_decap_8 FILLER_136_1320 ();
 sg13g2_decap_8 FILLER_136_1327 ();
 sg13g2_decap_8 FILLER_136_1337 ();
 sg13g2_decap_8 FILLER_136_1344 ();
 sg13g2_fill_1 FILLER_136_1351 ();
 sg13g2_decap_8 FILLER_136_1362 ();
 sg13g2_decap_8 FILLER_136_1369 ();
 sg13g2_decap_8 FILLER_136_1376 ();
 sg13g2_decap_8 FILLER_136_1383 ();
 sg13g2_decap_8 FILLER_136_1390 ();
 sg13g2_decap_8 FILLER_136_1405 ();
 sg13g2_decap_8 FILLER_136_1412 ();
 sg13g2_fill_2 FILLER_136_1419 ();
 sg13g2_decap_8 FILLER_136_1429 ();
 sg13g2_fill_2 FILLER_136_1436 ();
 sg13g2_decap_8 FILLER_136_1472 ();
 sg13g2_decap_8 FILLER_136_1479 ();
 sg13g2_decap_8 FILLER_136_1486 ();
 sg13g2_decap_8 FILLER_136_1493 ();
 sg13g2_decap_8 FILLER_136_1500 ();
 sg13g2_fill_2 FILLER_136_1507 ();
 sg13g2_fill_1 FILLER_136_1509 ();
 sg13g2_decap_4 FILLER_136_1518 ();
 sg13g2_fill_2 FILLER_136_1522 ();
 sg13g2_decap_8 FILLER_136_1532 ();
 sg13g2_decap_8 FILLER_136_1539 ();
 sg13g2_decap_8 FILLER_136_1546 ();
 sg13g2_fill_2 FILLER_136_1553 ();
 sg13g2_fill_1 FILLER_136_1555 ();
 sg13g2_decap_8 FILLER_136_1570 ();
 sg13g2_decap_8 FILLER_136_1577 ();
 sg13g2_decap_8 FILLER_136_1584 ();
 sg13g2_decap_8 FILLER_136_1591 ();
 sg13g2_decap_4 FILLER_136_1598 ();
 sg13g2_decap_4 FILLER_136_1607 ();
 sg13g2_fill_1 FILLER_136_1611 ();
 sg13g2_decap_8 FILLER_136_1616 ();
 sg13g2_decap_8 FILLER_136_1636 ();
 sg13g2_decap_8 FILLER_136_1643 ();
 sg13g2_decap_8 FILLER_136_1650 ();
 sg13g2_decap_8 FILLER_136_1657 ();
 sg13g2_fill_2 FILLER_136_1664 ();
 sg13g2_decap_4 FILLER_136_1674 ();
 sg13g2_fill_2 FILLER_136_1678 ();
 sg13g2_decap_4 FILLER_136_1701 ();
 sg13g2_fill_1 FILLER_136_1705 ();
 sg13g2_decap_8 FILLER_136_1709 ();
 sg13g2_decap_8 FILLER_136_1721 ();
 sg13g2_decap_8 FILLER_136_1728 ();
 sg13g2_decap_8 FILLER_136_1735 ();
 sg13g2_decap_8 FILLER_136_1742 ();
 sg13g2_decap_8 FILLER_136_1749 ();
 sg13g2_decap_8 FILLER_136_1756 ();
 sg13g2_decap_4 FILLER_136_1763 ();
 sg13g2_fill_1 FILLER_136_1767 ();
 sg13g2_decap_8 FILLER_137_0 ();
 sg13g2_decap_8 FILLER_137_7 ();
 sg13g2_decap_8 FILLER_137_14 ();
 sg13g2_decap_8 FILLER_137_21 ();
 sg13g2_decap_8 FILLER_137_28 ();
 sg13g2_decap_8 FILLER_137_44 ();
 sg13g2_decap_8 FILLER_137_65 ();
 sg13g2_decap_8 FILLER_137_72 ();
 sg13g2_decap_8 FILLER_137_79 ();
 sg13g2_decap_8 FILLER_137_86 ();
 sg13g2_decap_8 FILLER_137_93 ();
 sg13g2_decap_8 FILLER_137_100 ();
 sg13g2_decap_8 FILLER_137_107 ();
 sg13g2_decap_8 FILLER_137_114 ();
 sg13g2_decap_8 FILLER_137_121 ();
 sg13g2_decap_8 FILLER_137_128 ();
 sg13g2_fill_1 FILLER_137_135 ();
 sg13g2_fill_1 FILLER_137_153 ();
 sg13g2_decap_8 FILLER_137_162 ();
 sg13g2_decap_8 FILLER_137_169 ();
 sg13g2_decap_8 FILLER_137_176 ();
 sg13g2_decap_8 FILLER_137_183 ();
 sg13g2_decap_8 FILLER_137_190 ();
 sg13g2_decap_8 FILLER_137_197 ();
 sg13g2_decap_8 FILLER_137_204 ();
 sg13g2_fill_2 FILLER_137_211 ();
 sg13g2_fill_1 FILLER_137_213 ();
 sg13g2_decap_8 FILLER_137_222 ();
 sg13g2_decap_8 FILLER_137_229 ();
 sg13g2_decap_8 FILLER_137_236 ();
 sg13g2_fill_2 FILLER_137_243 ();
 sg13g2_fill_1 FILLER_137_245 ();
 sg13g2_decap_8 FILLER_137_250 ();
 sg13g2_fill_2 FILLER_137_273 ();
 sg13g2_fill_1 FILLER_137_275 ();
 sg13g2_decap_8 FILLER_137_288 ();
 sg13g2_decap_8 FILLER_137_295 ();
 sg13g2_decap_8 FILLER_137_302 ();
 sg13g2_decap_8 FILLER_137_309 ();
 sg13g2_decap_8 FILLER_137_316 ();
 sg13g2_decap_8 FILLER_137_323 ();
 sg13g2_decap_8 FILLER_137_356 ();
 sg13g2_decap_8 FILLER_137_363 ();
 sg13g2_decap_8 FILLER_137_370 ();
 sg13g2_decap_8 FILLER_137_377 ();
 sg13g2_decap_8 FILLER_137_384 ();
 sg13g2_fill_2 FILLER_137_391 ();
 sg13g2_fill_1 FILLER_137_393 ();
 sg13g2_decap_8 FILLER_137_398 ();
 sg13g2_fill_2 FILLER_137_405 ();
 sg13g2_fill_1 FILLER_137_407 ();
 sg13g2_decap_8 FILLER_137_420 ();
 sg13g2_decap_4 FILLER_137_427 ();
 sg13g2_fill_2 FILLER_137_448 ();
 sg13g2_fill_1 FILLER_137_450 ();
 sg13g2_decap_8 FILLER_137_479 ();
 sg13g2_decap_8 FILLER_137_486 ();
 sg13g2_decap_8 FILLER_137_493 ();
 sg13g2_decap_8 FILLER_137_500 ();
 sg13g2_fill_2 FILLER_137_525 ();
 sg13g2_decap_8 FILLER_137_534 ();
 sg13g2_decap_8 FILLER_137_541 ();
 sg13g2_decap_8 FILLER_137_548 ();
 sg13g2_decap_8 FILLER_137_555 ();
 sg13g2_decap_8 FILLER_137_562 ();
 sg13g2_decap_4 FILLER_137_569 ();
 sg13g2_fill_1 FILLER_137_573 ();
 sg13g2_decap_8 FILLER_137_613 ();
 sg13g2_decap_8 FILLER_137_620 ();
 sg13g2_decap_8 FILLER_137_627 ();
 sg13g2_decap_8 FILLER_137_634 ();
 sg13g2_decap_8 FILLER_137_641 ();
 sg13g2_decap_8 FILLER_137_648 ();
 sg13g2_decap_8 FILLER_137_655 ();
 sg13g2_decap_8 FILLER_137_662 ();
 sg13g2_decap_8 FILLER_137_669 ();
 sg13g2_decap_8 FILLER_137_676 ();
 sg13g2_decap_8 FILLER_137_683 ();
 sg13g2_decap_8 FILLER_137_690 ();
 sg13g2_fill_1 FILLER_137_697 ();
 sg13g2_decap_8 FILLER_137_710 ();
 sg13g2_decap_8 FILLER_137_717 ();
 sg13g2_fill_1 FILLER_137_724 ();
 sg13g2_decap_8 FILLER_137_731 ();
 sg13g2_decap_8 FILLER_137_738 ();
 sg13g2_decap_4 FILLER_137_745 ();
 sg13g2_fill_2 FILLER_137_749 ();
 sg13g2_decap_8 FILLER_137_771 ();
 sg13g2_decap_8 FILLER_137_778 ();
 sg13g2_fill_2 FILLER_137_785 ();
 sg13g2_fill_1 FILLER_137_800 ();
 sg13g2_decap_8 FILLER_137_813 ();
 sg13g2_decap_8 FILLER_137_820 ();
 sg13g2_decap_8 FILLER_137_827 ();
 sg13g2_decap_8 FILLER_137_834 ();
 sg13g2_decap_8 FILLER_137_841 ();
 sg13g2_decap_8 FILLER_137_848 ();
 sg13g2_decap_8 FILLER_137_855 ();
 sg13g2_decap_8 FILLER_137_862 ();
 sg13g2_decap_8 FILLER_137_869 ();
 sg13g2_fill_2 FILLER_137_876 ();
 sg13g2_fill_1 FILLER_137_878 ();
 sg13g2_decap_8 FILLER_137_882 ();
 sg13g2_decap_8 FILLER_137_889 ();
 sg13g2_decap_8 FILLER_137_896 ();
 sg13g2_decap_8 FILLER_137_903 ();
 sg13g2_decap_8 FILLER_137_910 ();
 sg13g2_decap_8 FILLER_137_917 ();
 sg13g2_decap_8 FILLER_137_924 ();
 sg13g2_decap_4 FILLER_137_931 ();
 sg13g2_fill_1 FILLER_137_935 ();
 sg13g2_decap_8 FILLER_137_939 ();
 sg13g2_decap_8 FILLER_137_946 ();
 sg13g2_decap_8 FILLER_137_953 ();
 sg13g2_decap_8 FILLER_137_960 ();
 sg13g2_fill_1 FILLER_137_967 ();
 sg13g2_decap_4 FILLER_137_974 ();
 sg13g2_decap_8 FILLER_137_990 ();
 sg13g2_decap_8 FILLER_137_997 ();
 sg13g2_decap_8 FILLER_137_1004 ();
 sg13g2_decap_8 FILLER_137_1011 ();
 sg13g2_decap_8 FILLER_137_1018 ();
 sg13g2_decap_8 FILLER_137_1025 ();
 sg13g2_decap_8 FILLER_137_1032 ();
 sg13g2_decap_4 FILLER_137_1039 ();
 sg13g2_fill_2 FILLER_137_1043 ();
 sg13g2_decap_4 FILLER_137_1050 ();
 sg13g2_fill_1 FILLER_137_1054 ();
 sg13g2_decap_8 FILLER_137_1063 ();
 sg13g2_decap_8 FILLER_137_1070 ();
 sg13g2_decap_8 FILLER_137_1082 ();
 sg13g2_fill_2 FILLER_137_1089 ();
 sg13g2_fill_1 FILLER_137_1091 ();
 sg13g2_decap_8 FILLER_137_1096 ();
 sg13g2_decap_4 FILLER_137_1103 ();
 sg13g2_fill_2 FILLER_137_1107 ();
 sg13g2_decap_8 FILLER_137_1152 ();
 sg13g2_fill_1 FILLER_137_1159 ();
 sg13g2_fill_1 FILLER_137_1167 ();
 sg13g2_fill_2 FILLER_137_1178 ();
 sg13g2_fill_1 FILLER_137_1180 ();
 sg13g2_decap_8 FILLER_137_1186 ();
 sg13g2_decap_4 FILLER_137_1193 ();
 sg13g2_fill_1 FILLER_137_1197 ();
 sg13g2_fill_2 FILLER_137_1211 ();
 sg13g2_fill_2 FILLER_137_1217 ();
 sg13g2_fill_2 FILLER_137_1232 ();
 sg13g2_fill_1 FILLER_137_1234 ();
 sg13g2_fill_2 FILLER_137_1243 ();
 sg13g2_fill_1 FILLER_137_1245 ();
 sg13g2_decap_8 FILLER_137_1254 ();
 sg13g2_decap_8 FILLER_137_1261 ();
 sg13g2_decap_8 FILLER_137_1268 ();
 sg13g2_decap_4 FILLER_137_1275 ();
 sg13g2_fill_1 FILLER_137_1279 ();
 sg13g2_fill_2 FILLER_137_1297 ();
 sg13g2_decap_8 FILLER_137_1316 ();
 sg13g2_decap_4 FILLER_137_1323 ();
 sg13g2_fill_2 FILLER_137_1327 ();
 sg13g2_decap_8 FILLER_137_1338 ();
 sg13g2_fill_2 FILLER_137_1345 ();
 sg13g2_decap_8 FILLER_137_1351 ();
 sg13g2_decap_8 FILLER_137_1358 ();
 sg13g2_decap_8 FILLER_137_1365 ();
 sg13g2_decap_8 FILLER_137_1372 ();
 sg13g2_decap_8 FILLER_137_1379 ();
 sg13g2_decap_8 FILLER_137_1410 ();
 sg13g2_decap_8 FILLER_137_1417 ();
 sg13g2_decap_8 FILLER_137_1424 ();
 sg13g2_decap_4 FILLER_137_1439 ();
 sg13g2_fill_2 FILLER_137_1443 ();
 sg13g2_decap_8 FILLER_137_1479 ();
 sg13g2_decap_8 FILLER_137_1486 ();
 sg13g2_decap_8 FILLER_137_1493 ();
 sg13g2_fill_2 FILLER_137_1500 ();
 sg13g2_fill_1 FILLER_137_1502 ();
 sg13g2_decap_8 FILLER_137_1508 ();
 sg13g2_decap_4 FILLER_137_1515 ();
 sg13g2_decap_8 FILLER_137_1527 ();
 sg13g2_decap_8 FILLER_137_1534 ();
 sg13g2_decap_8 FILLER_137_1541 ();
 sg13g2_decap_8 FILLER_137_1548 ();
 sg13g2_decap_8 FILLER_137_1555 ();
 sg13g2_decap_8 FILLER_137_1562 ();
 sg13g2_decap_8 FILLER_137_1569 ();
 sg13g2_decap_8 FILLER_137_1576 ();
 sg13g2_decap_8 FILLER_137_1583 ();
 sg13g2_decap_8 FILLER_137_1590 ();
 sg13g2_decap_4 FILLER_137_1597 ();
 sg13g2_decap_8 FILLER_137_1640 ();
 sg13g2_decap_8 FILLER_137_1647 ();
 sg13g2_decap_8 FILLER_137_1654 ();
 sg13g2_decap_8 FILLER_137_1661 ();
 sg13g2_fill_2 FILLER_137_1668 ();
 sg13g2_fill_1 FILLER_137_1670 ();
 sg13g2_decap_8 FILLER_137_1683 ();
 sg13g2_decap_8 FILLER_137_1690 ();
 sg13g2_decap_4 FILLER_137_1697 ();
 sg13g2_fill_2 FILLER_137_1701 ();
 sg13g2_decap_4 FILLER_137_1711 ();
 sg13g2_decap_8 FILLER_137_1720 ();
 sg13g2_decap_8 FILLER_137_1727 ();
 sg13g2_decap_8 FILLER_137_1734 ();
 sg13g2_decap_8 FILLER_137_1741 ();
 sg13g2_decap_8 FILLER_137_1748 ();
 sg13g2_decap_8 FILLER_137_1755 ();
 sg13g2_decap_4 FILLER_137_1762 ();
 sg13g2_fill_2 FILLER_137_1766 ();
 sg13g2_decap_8 FILLER_138_0 ();
 sg13g2_decap_8 FILLER_138_7 ();
 sg13g2_decap_8 FILLER_138_14 ();
 sg13g2_decap_4 FILLER_138_21 ();
 sg13g2_fill_2 FILLER_138_25 ();
 sg13g2_decap_8 FILLER_138_36 ();
 sg13g2_decap_8 FILLER_138_43 ();
 sg13g2_decap_8 FILLER_138_50 ();
 sg13g2_decap_8 FILLER_138_57 ();
 sg13g2_decap_8 FILLER_138_64 ();
 sg13g2_decap_8 FILLER_138_71 ();
 sg13g2_decap_8 FILLER_138_78 ();
 sg13g2_decap_8 FILLER_138_85 ();
 sg13g2_decap_4 FILLER_138_92 ();
 sg13g2_decap_8 FILLER_138_104 ();
 sg13g2_decap_8 FILLER_138_111 ();
 sg13g2_decap_8 FILLER_138_118 ();
 sg13g2_fill_2 FILLER_138_125 ();
 sg13g2_decap_8 FILLER_138_135 ();
 sg13g2_decap_8 FILLER_138_155 ();
 sg13g2_decap_4 FILLER_138_162 ();
 sg13g2_decap_8 FILLER_138_182 ();
 sg13g2_decap_8 FILLER_138_189 ();
 sg13g2_decap_4 FILLER_138_196 ();
 sg13g2_fill_2 FILLER_138_200 ();
 sg13g2_decap_8 FILLER_138_210 ();
 sg13g2_decap_4 FILLER_138_217 ();
 sg13g2_fill_2 FILLER_138_221 ();
 sg13g2_decap_8 FILLER_138_226 ();
 sg13g2_fill_2 FILLER_138_233 ();
 sg13g2_fill_1 FILLER_138_235 ();
 sg13g2_decap_4 FILLER_138_255 ();
 sg13g2_fill_1 FILLER_138_259 ();
 sg13g2_fill_2 FILLER_138_268 ();
 sg13g2_fill_1 FILLER_138_270 ();
 sg13g2_decap_8 FILLER_138_276 ();
 sg13g2_decap_8 FILLER_138_283 ();
 sg13g2_fill_1 FILLER_138_290 ();
 sg13g2_decap_8 FILLER_138_295 ();
 sg13g2_decap_8 FILLER_138_302 ();
 sg13g2_decap_8 FILLER_138_309 ();
 sg13g2_decap_8 FILLER_138_316 ();
 sg13g2_fill_2 FILLER_138_323 ();
 sg13g2_fill_1 FILLER_138_325 ();
 sg13g2_decap_8 FILLER_138_335 ();
 sg13g2_decap_8 FILLER_138_342 ();
 sg13g2_decap_8 FILLER_138_349 ();
 sg13g2_decap_8 FILLER_138_356 ();
 sg13g2_fill_2 FILLER_138_363 ();
 sg13g2_fill_1 FILLER_138_365 ();
 sg13g2_decap_8 FILLER_138_379 ();
 sg13g2_decap_8 FILLER_138_386 ();
 sg13g2_decap_4 FILLER_138_398 ();
 sg13g2_fill_2 FILLER_138_406 ();
 sg13g2_decap_8 FILLER_138_429 ();
 sg13g2_decap_4 FILLER_138_436 ();
 sg13g2_fill_1 FILLER_138_440 ();
 sg13g2_decap_4 FILLER_138_449 ();
 sg13g2_fill_1 FILLER_138_453 ();
 sg13g2_decap_8 FILLER_138_482 ();
 sg13g2_decap_8 FILLER_138_489 ();
 sg13g2_decap_8 FILLER_138_496 ();
 sg13g2_decap_8 FILLER_138_503 ();
 sg13g2_fill_1 FILLER_138_515 ();
 sg13g2_fill_2 FILLER_138_525 ();
 sg13g2_fill_1 FILLER_138_527 ();
 sg13g2_decap_4 FILLER_138_541 ();
 sg13g2_fill_1 FILLER_138_545 ();
 sg13g2_fill_1 FILLER_138_550 ();
 sg13g2_decap_8 FILLER_138_555 ();
 sg13g2_decap_8 FILLER_138_562 ();
 sg13g2_decap_8 FILLER_138_569 ();
 sg13g2_decap_8 FILLER_138_576 ();
 sg13g2_decap_4 FILLER_138_583 ();
 sg13g2_fill_1 FILLER_138_587 ();
 sg13g2_decap_8 FILLER_138_610 ();
 sg13g2_decap_8 FILLER_138_617 ();
 sg13g2_fill_1 FILLER_138_624 ();
 sg13g2_decap_8 FILLER_138_630 ();
 sg13g2_decap_8 FILLER_138_641 ();
 sg13g2_decap_8 FILLER_138_648 ();
 sg13g2_decap_8 FILLER_138_655 ();
 sg13g2_decap_8 FILLER_138_662 ();
 sg13g2_fill_2 FILLER_138_669 ();
 sg13g2_decap_8 FILLER_138_683 ();
 sg13g2_decap_4 FILLER_138_690 ();
 sg13g2_fill_2 FILLER_138_694 ();
 sg13g2_decap_8 FILLER_138_701 ();
 sg13g2_decap_8 FILLER_138_708 ();
 sg13g2_decap_8 FILLER_138_715 ();
 sg13g2_decap_8 FILLER_138_722 ();
 sg13g2_decap_8 FILLER_138_729 ();
 sg13g2_decap_8 FILLER_138_736 ();
 sg13g2_decap_8 FILLER_138_743 ();
 sg13g2_decap_4 FILLER_138_750 ();
 sg13g2_decap_8 FILLER_138_765 ();
 sg13g2_decap_8 FILLER_138_772 ();
 sg13g2_decap_8 FILLER_138_779 ();
 sg13g2_decap_8 FILLER_138_786 ();
 sg13g2_decap_4 FILLER_138_793 ();
 sg13g2_fill_1 FILLER_138_797 ();
 sg13g2_fill_1 FILLER_138_821 ();
 sg13g2_decap_8 FILLER_138_826 ();
 sg13g2_fill_1 FILLER_138_833 ();
 sg13g2_decap_8 FILLER_138_851 ();
 sg13g2_decap_8 FILLER_138_858 ();
 sg13g2_fill_2 FILLER_138_877 ();
 sg13g2_decap_8 FILLER_138_889 ();
 sg13g2_decap_8 FILLER_138_896 ();
 sg13g2_decap_8 FILLER_138_903 ();
 sg13g2_decap_8 FILLER_138_910 ();
 sg13g2_decap_8 FILLER_138_917 ();
 sg13g2_fill_2 FILLER_138_924 ();
 sg13g2_fill_1 FILLER_138_943 ();
 sg13g2_decap_8 FILLER_138_949 ();
 sg13g2_decap_8 FILLER_138_956 ();
 sg13g2_decap_8 FILLER_138_963 ();
 sg13g2_decap_8 FILLER_138_970 ();
 sg13g2_decap_8 FILLER_138_977 ();
 sg13g2_decap_8 FILLER_138_984 ();
 sg13g2_decap_8 FILLER_138_991 ();
 sg13g2_decap_4 FILLER_138_998 ();
 sg13g2_fill_2 FILLER_138_1002 ();
 sg13g2_decap_8 FILLER_138_1012 ();
 sg13g2_decap_8 FILLER_138_1019 ();
 sg13g2_decap_8 FILLER_138_1026 ();
 sg13g2_decap_8 FILLER_138_1033 ();
 sg13g2_fill_2 FILLER_138_1040 ();
 sg13g2_decap_8 FILLER_138_1047 ();
 sg13g2_decap_8 FILLER_138_1054 ();
 sg13g2_fill_2 FILLER_138_1061 ();
 sg13g2_fill_1 FILLER_138_1063 ();
 sg13g2_decap_4 FILLER_138_1080 ();
 sg13g2_fill_2 FILLER_138_1084 ();
 sg13g2_fill_2 FILLER_138_1090 ();
 sg13g2_fill_2 FILLER_138_1104 ();
 sg13g2_decap_8 FILLER_138_1117 ();
 sg13g2_decap_8 FILLER_138_1124 ();
 sg13g2_decap_4 FILLER_138_1148 ();
 sg13g2_fill_1 FILLER_138_1169 ();
 sg13g2_decap_8 FILLER_138_1178 ();
 sg13g2_decap_8 FILLER_138_1185 ();
 sg13g2_decap_8 FILLER_138_1192 ();
 sg13g2_fill_2 FILLER_138_1199 ();
 sg13g2_decap_8 FILLER_138_1209 ();
 sg13g2_fill_2 FILLER_138_1216 ();
 sg13g2_fill_1 FILLER_138_1218 ();
 sg13g2_decap_8 FILLER_138_1235 ();
 sg13g2_decap_8 FILLER_138_1242 ();
 sg13g2_decap_4 FILLER_138_1249 ();
 sg13g2_fill_1 FILLER_138_1253 ();
 sg13g2_decap_8 FILLER_138_1262 ();
 sg13g2_decap_8 FILLER_138_1269 ();
 sg13g2_decap_8 FILLER_138_1276 ();
 sg13g2_decap_8 FILLER_138_1283 ();
 sg13g2_decap_8 FILLER_138_1290 ();
 sg13g2_decap_4 FILLER_138_1297 ();
 sg13g2_fill_1 FILLER_138_1301 ();
 sg13g2_decap_8 FILLER_138_1307 ();
 sg13g2_decap_8 FILLER_138_1314 ();
 sg13g2_fill_2 FILLER_138_1321 ();
 sg13g2_fill_1 FILLER_138_1323 ();
 sg13g2_fill_1 FILLER_138_1332 ();
 sg13g2_fill_2 FILLER_138_1341 ();
 sg13g2_fill_2 FILLER_138_1356 ();
 sg13g2_decap_8 FILLER_138_1366 ();
 sg13g2_decap_8 FILLER_138_1373 ();
 sg13g2_fill_1 FILLER_138_1380 ();
 sg13g2_fill_2 FILLER_138_1390 ();
 sg13g2_decap_8 FILLER_138_1404 ();
 sg13g2_fill_2 FILLER_138_1411 ();
 sg13g2_fill_1 FILLER_138_1413 ();
 sg13g2_decap_8 FILLER_138_1419 ();
 sg13g2_decap_8 FILLER_138_1426 ();
 sg13g2_decap_8 FILLER_138_1433 ();
 sg13g2_decap_8 FILLER_138_1440 ();
 sg13g2_decap_8 FILLER_138_1447 ();
 sg13g2_decap_4 FILLER_138_1454 ();
 sg13g2_fill_1 FILLER_138_1458 ();
 sg13g2_fill_1 FILLER_138_1464 ();
 sg13g2_decap_8 FILLER_138_1483 ();
 sg13g2_decap_4 FILLER_138_1490 ();
 sg13g2_fill_2 FILLER_138_1494 ();
 sg13g2_fill_1 FILLER_138_1509 ();
 sg13g2_fill_2 FILLER_138_1518 ();
 sg13g2_decap_8 FILLER_138_1533 ();
 sg13g2_decap_8 FILLER_138_1540 ();
 sg13g2_decap_4 FILLER_138_1547 ();
 sg13g2_fill_1 FILLER_138_1551 ();
 sg13g2_decap_8 FILLER_138_1568 ();
 sg13g2_decap_8 FILLER_138_1575 ();
 sg13g2_decap_8 FILLER_138_1582 ();
 sg13g2_decap_8 FILLER_138_1589 ();
 sg13g2_decap_8 FILLER_138_1596 ();
 sg13g2_fill_2 FILLER_138_1603 ();
 sg13g2_decap_8 FILLER_138_1618 ();
 sg13g2_decap_8 FILLER_138_1625 ();
 sg13g2_decap_8 FILLER_138_1632 ();
 sg13g2_decap_8 FILLER_138_1639 ();
 sg13g2_decap_8 FILLER_138_1646 ();
 sg13g2_decap_8 FILLER_138_1653 ();
 sg13g2_decap_4 FILLER_138_1660 ();
 sg13g2_fill_2 FILLER_138_1672 ();
 sg13g2_fill_1 FILLER_138_1674 ();
 sg13g2_decap_8 FILLER_138_1695 ();
 sg13g2_decap_8 FILLER_138_1702 ();
 sg13g2_decap_8 FILLER_138_1709 ();
 sg13g2_decap_8 FILLER_138_1716 ();
 sg13g2_decap_8 FILLER_138_1723 ();
 sg13g2_decap_8 FILLER_138_1730 ();
 sg13g2_decap_8 FILLER_138_1737 ();
 sg13g2_decap_8 FILLER_138_1744 ();
 sg13g2_decap_8 FILLER_138_1751 ();
 sg13g2_decap_8 FILLER_138_1758 ();
 sg13g2_fill_2 FILLER_138_1765 ();
 sg13g2_fill_1 FILLER_138_1767 ();
 sg13g2_decap_8 FILLER_139_0 ();
 sg13g2_decap_8 FILLER_139_7 ();
 sg13g2_decap_8 FILLER_139_14 ();
 sg13g2_decap_4 FILLER_139_21 ();
 sg13g2_fill_1 FILLER_139_25 ();
 sg13g2_decap_8 FILLER_139_43 ();
 sg13g2_decap_8 FILLER_139_50 ();
 sg13g2_decap_8 FILLER_139_57 ();
 sg13g2_decap_8 FILLER_139_64 ();
 sg13g2_decap_8 FILLER_139_71 ();
 sg13g2_decap_4 FILLER_139_78 ();
 sg13g2_fill_2 FILLER_139_82 ();
 sg13g2_decap_8 FILLER_139_105 ();
 sg13g2_decap_8 FILLER_139_112 ();
 sg13g2_decap_8 FILLER_139_119 ();
 sg13g2_decap_8 FILLER_139_126 ();
 sg13g2_decap_8 FILLER_139_133 ();
 sg13g2_decap_4 FILLER_139_140 ();
 sg13g2_fill_1 FILLER_139_144 ();
 sg13g2_decap_8 FILLER_139_152 ();
 sg13g2_decap_4 FILLER_139_159 ();
 sg13g2_decap_8 FILLER_139_176 ();
 sg13g2_decap_8 FILLER_139_183 ();
 sg13g2_decap_4 FILLER_139_190 ();
 sg13g2_decap_8 FILLER_139_198 ();
 sg13g2_decap_8 FILLER_139_205 ();
 sg13g2_decap_8 FILLER_139_212 ();
 sg13g2_decap_4 FILLER_139_219 ();
 sg13g2_decap_8 FILLER_139_235 ();
 sg13g2_decap_8 FILLER_139_242 ();
 sg13g2_decap_8 FILLER_139_249 ();
 sg13g2_decap_8 FILLER_139_256 ();
 sg13g2_decap_4 FILLER_139_263 ();
 sg13g2_decap_8 FILLER_139_271 ();
 sg13g2_decap_8 FILLER_139_278 ();
 sg13g2_fill_2 FILLER_139_285 ();
 sg13g2_decap_8 FILLER_139_296 ();
 sg13g2_decap_8 FILLER_139_303 ();
 sg13g2_decap_8 FILLER_139_310 ();
 sg13g2_decap_8 FILLER_139_317 ();
 sg13g2_fill_2 FILLER_139_324 ();
 sg13g2_decap_8 FILLER_139_335 ();
 sg13g2_decap_8 FILLER_139_342 ();
 sg13g2_decap_8 FILLER_139_349 ();
 sg13g2_decap_8 FILLER_139_356 ();
 sg13g2_decap_8 FILLER_139_363 ();
 sg13g2_decap_8 FILLER_139_370 ();
 sg13g2_decap_8 FILLER_139_377 ();
 sg13g2_fill_1 FILLER_139_384 ();
 sg13g2_fill_2 FILLER_139_398 ();
 sg13g2_decap_8 FILLER_139_408 ();
 sg13g2_decap_8 FILLER_139_420 ();
 sg13g2_decap_8 FILLER_139_427 ();
 sg13g2_decap_8 FILLER_139_434 ();
 sg13g2_decap_8 FILLER_139_441 ();
 sg13g2_decap_8 FILLER_139_448 ();
 sg13g2_decap_8 FILLER_139_455 ();
 sg13g2_decap_8 FILLER_139_462 ();
 sg13g2_fill_2 FILLER_139_469 ();
 sg13g2_decap_8 FILLER_139_479 ();
 sg13g2_decap_8 FILLER_139_486 ();
 sg13g2_decap_8 FILLER_139_493 ();
 sg13g2_decap_8 FILLER_139_500 ();
 sg13g2_decap_8 FILLER_139_507 ();
 sg13g2_decap_8 FILLER_139_514 ();
 sg13g2_decap_4 FILLER_139_521 ();
 sg13g2_fill_2 FILLER_139_530 ();
 sg13g2_fill_1 FILLER_139_532 ();
 sg13g2_fill_2 FILLER_139_543 ();
 sg13g2_fill_1 FILLER_139_545 ();
 sg13g2_decap_8 FILLER_139_568 ();
 sg13g2_decap_8 FILLER_139_575 ();
 sg13g2_decap_8 FILLER_139_582 ();
 sg13g2_fill_2 FILLER_139_605 ();
 sg13g2_fill_1 FILLER_139_607 ();
 sg13g2_decap_8 FILLER_139_613 ();
 sg13g2_decap_8 FILLER_139_620 ();
 sg13g2_decap_8 FILLER_139_627 ();
 sg13g2_fill_2 FILLER_139_634 ();
 sg13g2_decap_8 FILLER_139_644 ();
 sg13g2_decap_4 FILLER_139_651 ();
 sg13g2_decap_8 FILLER_139_665 ();
 sg13g2_decap_8 FILLER_139_672 ();
 sg13g2_decap_4 FILLER_139_679 ();
 sg13g2_fill_2 FILLER_139_683 ();
 sg13g2_fill_2 FILLER_139_693 ();
 sg13g2_fill_1 FILLER_139_695 ();
 sg13g2_decap_4 FILLER_139_704 ();
 sg13g2_decap_4 FILLER_139_713 ();
 sg13g2_fill_2 FILLER_139_717 ();
 sg13g2_decap_8 FILLER_139_723 ();
 sg13g2_decap_8 FILLER_139_730 ();
 sg13g2_decap_8 FILLER_139_737 ();
 sg13g2_decap_8 FILLER_139_744 ();
 sg13g2_decap_4 FILLER_139_751 ();
 sg13g2_decap_8 FILLER_139_767 ();
 sg13g2_decap_8 FILLER_139_774 ();
 sg13g2_decap_8 FILLER_139_781 ();
 sg13g2_decap_8 FILLER_139_788 ();
 sg13g2_decap_8 FILLER_139_795 ();
 sg13g2_decap_4 FILLER_139_802 ();
 sg13g2_fill_1 FILLER_139_806 ();
 sg13g2_decap_8 FILLER_139_811 ();
 sg13g2_decap_8 FILLER_139_821 ();
 sg13g2_decap_8 FILLER_139_828 ();
 sg13g2_decap_4 FILLER_139_835 ();
 sg13g2_fill_1 FILLER_139_839 ();
 sg13g2_decap_8 FILLER_139_851 ();
 sg13g2_decap_4 FILLER_139_858 ();
 sg13g2_fill_2 FILLER_139_862 ();
 sg13g2_decap_8 FILLER_139_896 ();
 sg13g2_decap_8 FILLER_139_903 ();
 sg13g2_decap_8 FILLER_139_923 ();
 sg13g2_decap_4 FILLER_139_930 ();
 sg13g2_decap_8 FILLER_139_942 ();
 sg13g2_decap_8 FILLER_139_949 ();
 sg13g2_decap_8 FILLER_139_965 ();
 sg13g2_decap_4 FILLER_139_972 ();
 sg13g2_fill_1 FILLER_139_976 ();
 sg13g2_fill_2 FILLER_139_982 ();
 sg13g2_fill_2 FILLER_139_989 ();
 sg13g2_fill_1 FILLER_139_991 ();
 sg13g2_decap_8 FILLER_139_1002 ();
 sg13g2_decap_8 FILLER_139_1009 ();
 sg13g2_decap_8 FILLER_139_1016 ();
 sg13g2_decap_8 FILLER_139_1023 ();
 sg13g2_decap_8 FILLER_139_1030 ();
 sg13g2_decap_8 FILLER_139_1054 ();
 sg13g2_decap_8 FILLER_139_1061 ();
 sg13g2_decap_8 FILLER_139_1068 ();
 sg13g2_decap_8 FILLER_139_1075 ();
 sg13g2_decap_8 FILLER_139_1082 ();
 sg13g2_decap_8 FILLER_139_1089 ();
 sg13g2_fill_2 FILLER_139_1096 ();
 sg13g2_decap_8 FILLER_139_1114 ();
 sg13g2_decap_8 FILLER_139_1121 ();
 sg13g2_decap_4 FILLER_139_1128 ();
 sg13g2_decap_8 FILLER_139_1142 ();
 sg13g2_decap_8 FILLER_139_1149 ();
 sg13g2_fill_1 FILLER_139_1156 ();
 sg13g2_decap_8 FILLER_139_1166 ();
 sg13g2_decap_8 FILLER_139_1173 ();
 sg13g2_decap_8 FILLER_139_1180 ();
 sg13g2_decap_8 FILLER_139_1187 ();
 sg13g2_decap_8 FILLER_139_1194 ();
 sg13g2_decap_8 FILLER_139_1201 ();
 sg13g2_decap_8 FILLER_139_1208 ();
 sg13g2_decap_8 FILLER_139_1215 ();
 sg13g2_decap_8 FILLER_139_1230 ();
 sg13g2_decap_8 FILLER_139_1237 ();
 sg13g2_decap_4 FILLER_139_1244 ();
 sg13g2_fill_1 FILLER_139_1248 ();
 sg13g2_decap_8 FILLER_139_1258 ();
 sg13g2_decap_8 FILLER_139_1265 ();
 sg13g2_decap_8 FILLER_139_1272 ();
 sg13g2_decap_8 FILLER_139_1279 ();
 sg13g2_fill_2 FILLER_139_1286 ();
 sg13g2_fill_1 FILLER_139_1288 ();
 sg13g2_decap_8 FILLER_139_1297 ();
 sg13g2_decap_8 FILLER_139_1304 ();
 sg13g2_decap_8 FILLER_139_1311 ();
 sg13g2_decap_8 FILLER_139_1318 ();
 sg13g2_decap_4 FILLER_139_1325 ();
 sg13g2_fill_2 FILLER_139_1333 ();
 sg13g2_fill_1 FILLER_139_1335 ();
 sg13g2_decap_8 FILLER_139_1354 ();
 sg13g2_decap_8 FILLER_139_1361 ();
 sg13g2_decap_8 FILLER_139_1368 ();
 sg13g2_decap_8 FILLER_139_1375 ();
 sg13g2_decap_8 FILLER_139_1382 ();
 sg13g2_fill_2 FILLER_139_1394 ();
 sg13g2_decap_4 FILLER_139_1409 ();
 sg13g2_fill_1 FILLER_139_1413 ();
 sg13g2_decap_8 FILLER_139_1422 ();
 sg13g2_decap_4 FILLER_139_1429 ();
 sg13g2_decap_8 FILLER_139_1436 ();
 sg13g2_decap_8 FILLER_139_1443 ();
 sg13g2_decap_8 FILLER_139_1450 ();
 sg13g2_decap_8 FILLER_139_1457 ();
 sg13g2_decap_8 FILLER_139_1464 ();
 sg13g2_fill_2 FILLER_139_1471 ();
 sg13g2_decap_8 FILLER_139_1491 ();
 sg13g2_decap_8 FILLER_139_1498 ();
 sg13g2_decap_8 FILLER_139_1505 ();
 sg13g2_decap_8 FILLER_139_1512 ();
 sg13g2_decap_8 FILLER_139_1519 ();
 sg13g2_decap_4 FILLER_139_1526 ();
 sg13g2_fill_1 FILLER_139_1530 ();
 sg13g2_decap_8 FILLER_139_1539 ();
 sg13g2_decap_8 FILLER_139_1546 ();
 sg13g2_decap_4 FILLER_139_1553 ();
 sg13g2_fill_2 FILLER_139_1557 ();
 sg13g2_decap_8 FILLER_139_1575 ();
 sg13g2_decap_8 FILLER_139_1582 ();
 sg13g2_decap_8 FILLER_139_1589 ();
 sg13g2_decap_8 FILLER_139_1596 ();
 sg13g2_decap_8 FILLER_139_1603 ();
 sg13g2_fill_2 FILLER_139_1610 ();
 sg13g2_decap_8 FILLER_139_1637 ();
 sg13g2_decap_8 FILLER_139_1644 ();
 sg13g2_decap_8 FILLER_139_1651 ();
 sg13g2_fill_1 FILLER_139_1658 ();
 sg13g2_decap_4 FILLER_139_1676 ();
 sg13g2_fill_1 FILLER_139_1680 ();
 sg13g2_decap_8 FILLER_139_1689 ();
 sg13g2_decap_8 FILLER_139_1696 ();
 sg13g2_decap_8 FILLER_139_1703 ();
 sg13g2_decap_8 FILLER_139_1710 ();
 sg13g2_decap_8 FILLER_139_1717 ();
 sg13g2_decap_8 FILLER_139_1724 ();
 sg13g2_decap_8 FILLER_139_1731 ();
 sg13g2_decap_8 FILLER_139_1738 ();
 sg13g2_decap_8 FILLER_139_1745 ();
 sg13g2_decap_8 FILLER_139_1752 ();
 sg13g2_decap_8 FILLER_139_1759 ();
 sg13g2_fill_2 FILLER_139_1766 ();
 sg13g2_decap_8 FILLER_140_0 ();
 sg13g2_decap_8 FILLER_140_7 ();
 sg13g2_decap_8 FILLER_140_14 ();
 sg13g2_decap_8 FILLER_140_64 ();
 sg13g2_decap_8 FILLER_140_71 ();
 sg13g2_decap_8 FILLER_140_78 ();
 sg13g2_decap_8 FILLER_140_85 ();
 sg13g2_decap_8 FILLER_140_92 ();
 sg13g2_decap_8 FILLER_140_99 ();
 sg13g2_fill_2 FILLER_140_106 ();
 sg13g2_decap_4 FILLER_140_113 ();
 sg13g2_fill_1 FILLER_140_117 ();
 sg13g2_decap_8 FILLER_140_127 ();
 sg13g2_decap_8 FILLER_140_134 ();
 sg13g2_decap_8 FILLER_140_141 ();
 sg13g2_decap_8 FILLER_140_148 ();
 sg13g2_decap_8 FILLER_140_155 ();
 sg13g2_decap_8 FILLER_140_162 ();
 sg13g2_decap_8 FILLER_140_169 ();
 sg13g2_decap_8 FILLER_140_176 ();
 sg13g2_fill_2 FILLER_140_183 ();
 sg13g2_fill_2 FILLER_140_193 ();
 sg13g2_decap_8 FILLER_140_203 ();
 sg13g2_decap_8 FILLER_140_210 ();
 sg13g2_decap_4 FILLER_140_217 ();
 sg13g2_fill_2 FILLER_140_221 ();
 sg13g2_decap_4 FILLER_140_239 ();
 sg13g2_decap_8 FILLER_140_247 ();
 sg13g2_decap_8 FILLER_140_263 ();
 sg13g2_decap_8 FILLER_140_270 ();
 sg13g2_decap_8 FILLER_140_277 ();
 sg13g2_decap_8 FILLER_140_284 ();
 sg13g2_decap_8 FILLER_140_291 ();
 sg13g2_decap_8 FILLER_140_298 ();
 sg13g2_decap_8 FILLER_140_305 ();
 sg13g2_decap_8 FILLER_140_312 ();
 sg13g2_fill_2 FILLER_140_319 ();
 sg13g2_decap_8 FILLER_140_372 ();
 sg13g2_fill_2 FILLER_140_379 ();
 sg13g2_fill_1 FILLER_140_381 ();
 sg13g2_decap_8 FILLER_140_391 ();
 sg13g2_decap_8 FILLER_140_398 ();
 sg13g2_decap_8 FILLER_140_405 ();
 sg13g2_decap_8 FILLER_140_412 ();
 sg13g2_decap_8 FILLER_140_419 ();
 sg13g2_decap_8 FILLER_140_426 ();
 sg13g2_decap_8 FILLER_140_433 ();
 sg13g2_decap_8 FILLER_140_440 ();
 sg13g2_decap_8 FILLER_140_447 ();
 sg13g2_decap_8 FILLER_140_454 ();
 sg13g2_decap_8 FILLER_140_461 ();
 sg13g2_decap_8 FILLER_140_468 ();
 sg13g2_decap_4 FILLER_140_475 ();
 sg13g2_fill_2 FILLER_140_479 ();
 sg13g2_decap_8 FILLER_140_494 ();
 sg13g2_decap_8 FILLER_140_501 ();
 sg13g2_decap_4 FILLER_140_508 ();
 sg13g2_fill_2 FILLER_140_512 ();
 sg13g2_fill_1 FILLER_140_543 ();
 sg13g2_decap_8 FILLER_140_548 ();
 sg13g2_decap_8 FILLER_140_555 ();
 sg13g2_decap_8 FILLER_140_562 ();
 sg13g2_decap_8 FILLER_140_569 ();
 sg13g2_decap_8 FILLER_140_576 ();
 sg13g2_fill_1 FILLER_140_583 ();
 sg13g2_decap_4 FILLER_140_589 ();
 sg13g2_fill_1 FILLER_140_593 ();
 sg13g2_decap_8 FILLER_140_602 ();
 sg13g2_decap_8 FILLER_140_609 ();
 sg13g2_decap_8 FILLER_140_616 ();
 sg13g2_decap_8 FILLER_140_623 ();
 sg13g2_decap_4 FILLER_140_634 ();
 sg13g2_fill_1 FILLER_140_638 ();
 sg13g2_decap_8 FILLER_140_658 ();
 sg13g2_decap_4 FILLER_140_665 ();
 sg13g2_fill_2 FILLER_140_669 ();
 sg13g2_decap_8 FILLER_140_679 ();
 sg13g2_decap_8 FILLER_140_686 ();
 sg13g2_fill_2 FILLER_140_703 ();
 sg13g2_fill_1 FILLER_140_713 ();
 sg13g2_decap_8 FILLER_140_718 ();
 sg13g2_decap_8 FILLER_140_725 ();
 sg13g2_decap_8 FILLER_140_732 ();
 sg13g2_decap_8 FILLER_140_739 ();
 sg13g2_decap_4 FILLER_140_746 ();
 sg13g2_fill_2 FILLER_140_750 ();
 sg13g2_decap_8 FILLER_140_777 ();
 sg13g2_decap_8 FILLER_140_784 ();
 sg13g2_decap_8 FILLER_140_791 ();
 sg13g2_decap_8 FILLER_140_798 ();
 sg13g2_decap_8 FILLER_140_805 ();
 sg13g2_fill_2 FILLER_140_812 ();
 sg13g2_fill_1 FILLER_140_814 ();
 sg13g2_decap_8 FILLER_140_822 ();
 sg13g2_fill_2 FILLER_140_829 ();
 sg13g2_fill_1 FILLER_140_831 ();
 sg13g2_decap_8 FILLER_140_840 ();
 sg13g2_decap_8 FILLER_140_847 ();
 sg13g2_decap_8 FILLER_140_854 ();
 sg13g2_decap_8 FILLER_140_861 ();
 sg13g2_decap_4 FILLER_140_868 ();
 sg13g2_fill_2 FILLER_140_876 ();
 sg13g2_decap_8 FILLER_140_887 ();
 sg13g2_decap_8 FILLER_140_894 ();
 sg13g2_decap_8 FILLER_140_901 ();
 sg13g2_decap_8 FILLER_140_908 ();
 sg13g2_decap_8 FILLER_140_915 ();
 sg13g2_decap_8 FILLER_140_922 ();
 sg13g2_decap_8 FILLER_140_929 ();
 sg13g2_decap_8 FILLER_140_936 ();
 sg13g2_fill_2 FILLER_140_943 ();
 sg13g2_fill_1 FILLER_140_945 ();
 sg13g2_fill_2 FILLER_140_949 ();
 sg13g2_fill_1 FILLER_140_951 ();
 sg13g2_decap_4 FILLER_140_957 ();
 sg13g2_fill_1 FILLER_140_966 ();
 sg13g2_fill_2 FILLER_140_992 ();
 sg13g2_fill_1 FILLER_140_994 ();
 sg13g2_decap_8 FILLER_140_1015 ();
 sg13g2_decap_8 FILLER_140_1022 ();
 sg13g2_fill_1 FILLER_140_1037 ();
 sg13g2_decap_8 FILLER_140_1041 ();
 sg13g2_decap_8 FILLER_140_1052 ();
 sg13g2_decap_8 FILLER_140_1059 ();
 sg13g2_decap_8 FILLER_140_1066 ();
 sg13g2_decap_8 FILLER_140_1073 ();
 sg13g2_decap_8 FILLER_140_1080 ();
 sg13g2_decap_8 FILLER_140_1087 ();
 sg13g2_decap_8 FILLER_140_1094 ();
 sg13g2_decap_8 FILLER_140_1101 ();
 sg13g2_decap_8 FILLER_140_1108 ();
 sg13g2_decap_8 FILLER_140_1115 ();
 sg13g2_decap_8 FILLER_140_1122 ();
 sg13g2_decap_8 FILLER_140_1129 ();
 sg13g2_decap_8 FILLER_140_1136 ();
 sg13g2_decap_8 FILLER_140_1143 ();
 sg13g2_decap_8 FILLER_140_1150 ();
 sg13g2_decap_8 FILLER_140_1162 ();
 sg13g2_decap_8 FILLER_140_1169 ();
 sg13g2_decap_8 FILLER_140_1176 ();
 sg13g2_decap_8 FILLER_140_1183 ();
 sg13g2_decap_8 FILLER_140_1190 ();
 sg13g2_decap_8 FILLER_140_1197 ();
 sg13g2_decap_8 FILLER_140_1204 ();
 sg13g2_decap_8 FILLER_140_1211 ();
 sg13g2_decap_8 FILLER_140_1218 ();
 sg13g2_decap_8 FILLER_140_1225 ();
 sg13g2_decap_4 FILLER_140_1232 ();
 sg13g2_fill_2 FILLER_140_1236 ();
 sg13g2_decap_8 FILLER_140_1243 ();
 sg13g2_decap_4 FILLER_140_1250 ();
 sg13g2_fill_1 FILLER_140_1254 ();
 sg13g2_decap_8 FILLER_140_1263 ();
 sg13g2_fill_2 FILLER_140_1270 ();
 sg13g2_fill_1 FILLER_140_1284 ();
 sg13g2_decap_8 FILLER_140_1293 ();
 sg13g2_decap_4 FILLER_140_1300 ();
 sg13g2_fill_2 FILLER_140_1304 ();
 sg13g2_decap_8 FILLER_140_1309 ();
 sg13g2_decap_8 FILLER_140_1316 ();
 sg13g2_decap_8 FILLER_140_1323 ();
 sg13g2_decap_8 FILLER_140_1330 ();
 sg13g2_fill_2 FILLER_140_1337 ();
 sg13g2_fill_1 FILLER_140_1339 ();
 sg13g2_decap_4 FILLER_140_1348 ();
 sg13g2_decap_8 FILLER_140_1364 ();
 sg13g2_decap_8 FILLER_140_1371 ();
 sg13g2_decap_4 FILLER_140_1378 ();
 sg13g2_fill_1 FILLER_140_1395 ();
 sg13g2_decap_8 FILLER_140_1416 ();
 sg13g2_decap_8 FILLER_140_1423 ();
 sg13g2_decap_8 FILLER_140_1430 ();
 sg13g2_decap_8 FILLER_140_1437 ();
 sg13g2_decap_8 FILLER_140_1444 ();
 sg13g2_decap_8 FILLER_140_1451 ();
 sg13g2_decap_8 FILLER_140_1458 ();
 sg13g2_decap_8 FILLER_140_1465 ();
 sg13g2_decap_4 FILLER_140_1472 ();
 sg13g2_decap_8 FILLER_140_1498 ();
 sg13g2_decap_4 FILLER_140_1505 ();
 sg13g2_decap_8 FILLER_140_1518 ();
 sg13g2_decap_8 FILLER_140_1525 ();
 sg13g2_decap_8 FILLER_140_1532 ();
 sg13g2_decap_8 FILLER_140_1539 ();
 sg13g2_decap_8 FILLER_140_1546 ();
 sg13g2_decap_8 FILLER_140_1553 ();
 sg13g2_decap_8 FILLER_140_1560 ();
 sg13g2_decap_4 FILLER_140_1576 ();
 sg13g2_decap_8 FILLER_140_1587 ();
 sg13g2_decap_8 FILLER_140_1594 ();
 sg13g2_decap_8 FILLER_140_1601 ();
 sg13g2_decap_8 FILLER_140_1608 ();
 sg13g2_decap_8 FILLER_140_1615 ();
 sg13g2_decap_8 FILLER_140_1622 ();
 sg13g2_decap_8 FILLER_140_1629 ();
 sg13g2_decap_8 FILLER_140_1636 ();
 sg13g2_decap_8 FILLER_140_1643 ();
 sg13g2_decap_8 FILLER_140_1650 ();
 sg13g2_decap_8 FILLER_140_1657 ();
 sg13g2_fill_1 FILLER_140_1664 ();
 sg13g2_decap_8 FILLER_140_1685 ();
 sg13g2_decap_8 FILLER_140_1692 ();
 sg13g2_decap_8 FILLER_140_1699 ();
 sg13g2_decap_8 FILLER_140_1706 ();
 sg13g2_decap_8 FILLER_140_1713 ();
 sg13g2_decap_8 FILLER_140_1720 ();
 sg13g2_decap_8 FILLER_140_1727 ();
 sg13g2_decap_8 FILLER_140_1734 ();
 sg13g2_decap_8 FILLER_140_1741 ();
 sg13g2_decap_8 FILLER_140_1748 ();
 sg13g2_decap_8 FILLER_140_1755 ();
 sg13g2_decap_4 FILLER_140_1762 ();
 sg13g2_fill_2 FILLER_140_1766 ();
 sg13g2_decap_8 FILLER_141_0 ();
 sg13g2_decap_8 FILLER_141_7 ();
 sg13g2_decap_8 FILLER_141_14 ();
 sg13g2_fill_2 FILLER_141_21 ();
 sg13g2_fill_2 FILLER_141_48 ();
 sg13g2_fill_1 FILLER_141_50 ();
 sg13g2_decap_8 FILLER_141_64 ();
 sg13g2_decap_8 FILLER_141_71 ();
 sg13g2_decap_8 FILLER_141_78 ();
 sg13g2_decap_8 FILLER_141_93 ();
 sg13g2_decap_4 FILLER_141_100 ();
 sg13g2_fill_1 FILLER_141_104 ();
 sg13g2_decap_8 FILLER_141_133 ();
 sg13g2_decap_8 FILLER_141_140 ();
 sg13g2_decap_8 FILLER_141_147 ();
 sg13g2_decap_8 FILLER_141_154 ();
 sg13g2_decap_8 FILLER_141_161 ();
 sg13g2_decap_8 FILLER_141_168 ();
 sg13g2_decap_8 FILLER_141_175 ();
 sg13g2_decap_4 FILLER_141_182 ();
 sg13g2_fill_2 FILLER_141_196 ();
 sg13g2_fill_1 FILLER_141_198 ();
 sg13g2_fill_2 FILLER_141_207 ();
 sg13g2_fill_2 FILLER_141_218 ();
 sg13g2_decap_8 FILLER_141_248 ();
 sg13g2_decap_4 FILLER_141_255 ();
 sg13g2_fill_2 FILLER_141_259 ();
 sg13g2_decap_8 FILLER_141_279 ();
 sg13g2_decap_8 FILLER_141_286 ();
 sg13g2_decap_8 FILLER_141_293 ();
 sg13g2_fill_1 FILLER_141_300 ();
 sg13g2_decap_8 FILLER_141_349 ();
 sg13g2_decap_8 FILLER_141_356 ();
 sg13g2_decap_8 FILLER_141_363 ();
 sg13g2_decap_8 FILLER_141_370 ();
 sg13g2_decap_8 FILLER_141_377 ();
 sg13g2_decap_8 FILLER_141_384 ();
 sg13g2_fill_1 FILLER_141_391 ();
 sg13g2_decap_8 FILLER_141_396 ();
 sg13g2_decap_8 FILLER_141_403 ();
 sg13g2_decap_8 FILLER_141_410 ();
 sg13g2_decap_8 FILLER_141_417 ();
 sg13g2_decap_8 FILLER_141_424 ();
 sg13g2_decap_8 FILLER_141_431 ();
 sg13g2_decap_8 FILLER_141_438 ();
 sg13g2_decap_8 FILLER_141_445 ();
 sg13g2_decap_8 FILLER_141_452 ();
 sg13g2_decap_4 FILLER_141_459 ();
 sg13g2_fill_2 FILLER_141_463 ();
 sg13g2_decap_8 FILLER_141_483 ();
 sg13g2_decap_8 FILLER_141_490 ();
 sg13g2_decap_8 FILLER_141_497 ();
 sg13g2_decap_8 FILLER_141_504 ();
 sg13g2_fill_1 FILLER_141_511 ();
 sg13g2_decap_8 FILLER_141_533 ();
 sg13g2_decap_8 FILLER_141_540 ();
 sg13g2_decap_8 FILLER_141_547 ();
 sg13g2_decap_8 FILLER_141_554 ();
 sg13g2_decap_8 FILLER_141_561 ();
 sg13g2_decap_8 FILLER_141_568 ();
 sg13g2_decap_4 FILLER_141_575 ();
 sg13g2_fill_1 FILLER_141_579 ();
 sg13g2_decap_8 FILLER_141_601 ();
 sg13g2_decap_8 FILLER_141_608 ();
 sg13g2_decap_4 FILLER_141_615 ();
 sg13g2_fill_2 FILLER_141_623 ();
 sg13g2_decap_4 FILLER_141_629 ();
 sg13g2_fill_1 FILLER_141_633 ();
 sg13g2_decap_8 FILLER_141_648 ();
 sg13g2_decap_8 FILLER_141_655 ();
 sg13g2_decap_4 FILLER_141_662 ();
 sg13g2_fill_1 FILLER_141_666 ();
 sg13g2_decap_8 FILLER_141_680 ();
 sg13g2_decap_8 FILLER_141_692 ();
 sg13g2_fill_2 FILLER_141_699 ();
 sg13g2_fill_1 FILLER_141_701 ();
 sg13g2_fill_2 FILLER_141_706 ();
 sg13g2_fill_2 FILLER_141_719 ();
 sg13g2_fill_1 FILLER_141_721 ();
 sg13g2_decap_8 FILLER_141_730 ();
 sg13g2_decap_8 FILLER_141_737 ();
 sg13g2_decap_8 FILLER_141_744 ();
 sg13g2_fill_2 FILLER_141_751 ();
 sg13g2_fill_1 FILLER_141_753 ();
 sg13g2_decap_8 FILLER_141_765 ();
 sg13g2_decap_8 FILLER_141_772 ();
 sg13g2_decap_8 FILLER_141_779 ();
 sg13g2_decap_8 FILLER_141_786 ();
 sg13g2_decap_8 FILLER_141_793 ();
 sg13g2_decap_8 FILLER_141_800 ();
 sg13g2_decap_8 FILLER_141_807 ();
 sg13g2_decap_4 FILLER_141_814 ();
 sg13g2_decap_8 FILLER_141_846 ();
 sg13g2_decap_4 FILLER_141_853 ();
 sg13g2_fill_1 FILLER_141_857 ();
 sg13g2_decap_4 FILLER_141_863 ();
 sg13g2_fill_1 FILLER_141_867 ();
 sg13g2_fill_1 FILLER_141_880 ();
 sg13g2_decap_8 FILLER_141_894 ();
 sg13g2_decap_8 FILLER_141_901 ();
 sg13g2_decap_8 FILLER_141_908 ();
 sg13g2_fill_2 FILLER_141_915 ();
 sg13g2_fill_1 FILLER_141_917 ();
 sg13g2_decap_8 FILLER_141_927 ();
 sg13g2_decap_8 FILLER_141_934 ();
 sg13g2_decap_4 FILLER_141_941 ();
 sg13g2_fill_1 FILLER_141_945 ();
 sg13g2_fill_2 FILLER_141_961 ();
 sg13g2_fill_1 FILLER_141_963 ();
 sg13g2_decap_8 FILLER_141_975 ();
 sg13g2_decap_8 FILLER_141_982 ();
 sg13g2_fill_1 FILLER_141_989 ();
 sg13g2_decap_8 FILLER_141_995 ();
 sg13g2_decap_8 FILLER_141_1002 ();
 sg13g2_decap_4 FILLER_141_1009 ();
 sg13g2_fill_1 FILLER_141_1013 ();
 sg13g2_decap_4 FILLER_141_1027 ();
 sg13g2_fill_2 FILLER_141_1031 ();
 sg13g2_decap_8 FILLER_141_1062 ();
 sg13g2_fill_2 FILLER_141_1069 ();
 sg13g2_fill_1 FILLER_141_1071 ();
 sg13g2_decap_8 FILLER_141_1081 ();
 sg13g2_decap_8 FILLER_141_1088 ();
 sg13g2_decap_8 FILLER_141_1095 ();
 sg13g2_decap_8 FILLER_141_1102 ();
 sg13g2_decap_8 FILLER_141_1109 ();
 sg13g2_decap_8 FILLER_141_1116 ();
 sg13g2_decap_4 FILLER_141_1123 ();
 sg13g2_fill_1 FILLER_141_1127 ();
 sg13g2_decap_8 FILLER_141_1145 ();
 sg13g2_fill_2 FILLER_141_1152 ();
 sg13g2_fill_1 FILLER_141_1154 ();
 sg13g2_decap_8 FILLER_141_1159 ();
 sg13g2_decap_8 FILLER_141_1166 ();
 sg13g2_decap_8 FILLER_141_1173 ();
 sg13g2_decap_8 FILLER_141_1180 ();
 sg13g2_decap_8 FILLER_141_1187 ();
 sg13g2_decap_8 FILLER_141_1202 ();
 sg13g2_decap_8 FILLER_141_1209 ();
 sg13g2_decap_4 FILLER_141_1216 ();
 sg13g2_fill_1 FILLER_141_1220 ();
 sg13g2_decap_4 FILLER_141_1232 ();
 sg13g2_fill_1 FILLER_141_1236 ();
 sg13g2_decap_8 FILLER_141_1245 ();
 sg13g2_decap_8 FILLER_141_1252 ();
 sg13g2_decap_8 FILLER_141_1259 ();
 sg13g2_decap_8 FILLER_141_1266 ();
 sg13g2_decap_4 FILLER_141_1273 ();
 sg13g2_decap_8 FILLER_141_1298 ();
 sg13g2_fill_1 FILLER_141_1305 ();
 sg13g2_decap_4 FILLER_141_1314 ();
 sg13g2_decap_8 FILLER_141_1322 ();
 sg13g2_decap_8 FILLER_141_1329 ();
 sg13g2_fill_1 FILLER_141_1336 ();
 sg13g2_decap_4 FILLER_141_1342 ();
 sg13g2_fill_1 FILLER_141_1346 ();
 sg13g2_decap_8 FILLER_141_1355 ();
 sg13g2_decap_8 FILLER_141_1362 ();
 sg13g2_decap_8 FILLER_141_1369 ();
 sg13g2_decap_8 FILLER_141_1376 ();
 sg13g2_fill_1 FILLER_141_1383 ();
 sg13g2_decap_8 FILLER_141_1387 ();
 sg13g2_decap_8 FILLER_141_1399 ();
 sg13g2_decap_8 FILLER_141_1406 ();
 sg13g2_decap_8 FILLER_141_1413 ();
 sg13g2_decap_8 FILLER_141_1420 ();
 sg13g2_decap_4 FILLER_141_1427 ();
 sg13g2_fill_1 FILLER_141_1431 ();
 sg13g2_decap_4 FILLER_141_1440 ();
 sg13g2_fill_1 FILLER_141_1444 ();
 sg13g2_decap_8 FILLER_141_1454 ();
 sg13g2_decap_8 FILLER_141_1461 ();
 sg13g2_decap_4 FILLER_141_1468 ();
 sg13g2_fill_2 FILLER_141_1472 ();
 sg13g2_decap_8 FILLER_141_1485 ();
 sg13g2_decap_8 FILLER_141_1492 ();
 sg13g2_decap_8 FILLER_141_1499 ();
 sg13g2_fill_1 FILLER_141_1506 ();
 sg13g2_decap_8 FILLER_141_1527 ();
 sg13g2_decap_8 FILLER_141_1534 ();
 sg13g2_decap_8 FILLER_141_1541 ();
 sg13g2_decap_8 FILLER_141_1548 ();
 sg13g2_decap_8 FILLER_141_1555 ();
 sg13g2_fill_1 FILLER_141_1562 ();
 sg13g2_decap_8 FILLER_141_1592 ();
 sg13g2_decap_8 FILLER_141_1599 ();
 sg13g2_decap_8 FILLER_141_1606 ();
 sg13g2_decap_8 FILLER_141_1613 ();
 sg13g2_decap_8 FILLER_141_1620 ();
 sg13g2_decap_8 FILLER_141_1627 ();
 sg13g2_decap_8 FILLER_141_1634 ();
 sg13g2_decap_8 FILLER_141_1641 ();
 sg13g2_decap_8 FILLER_141_1648 ();
 sg13g2_decap_8 FILLER_141_1655 ();
 sg13g2_decap_8 FILLER_141_1662 ();
 sg13g2_decap_8 FILLER_141_1669 ();
 sg13g2_decap_8 FILLER_141_1676 ();
 sg13g2_decap_8 FILLER_141_1683 ();
 sg13g2_decap_8 FILLER_141_1690 ();
 sg13g2_decap_8 FILLER_141_1697 ();
 sg13g2_decap_8 FILLER_141_1704 ();
 sg13g2_decap_8 FILLER_141_1711 ();
 sg13g2_decap_8 FILLER_141_1718 ();
 sg13g2_decap_8 FILLER_141_1725 ();
 sg13g2_decap_8 FILLER_141_1732 ();
 sg13g2_decap_8 FILLER_141_1739 ();
 sg13g2_decap_8 FILLER_141_1746 ();
 sg13g2_decap_8 FILLER_141_1753 ();
 sg13g2_decap_8 FILLER_141_1760 ();
 sg13g2_fill_1 FILLER_141_1767 ();
 sg13g2_decap_8 FILLER_142_0 ();
 sg13g2_decap_8 FILLER_142_7 ();
 sg13g2_decap_8 FILLER_142_14 ();
 sg13g2_fill_2 FILLER_142_21 ();
 sg13g2_fill_1 FILLER_142_23 ();
 sg13g2_decap_8 FILLER_142_32 ();
 sg13g2_fill_2 FILLER_142_39 ();
 sg13g2_fill_1 FILLER_142_41 ();
 sg13g2_fill_2 FILLER_142_47 ();
 sg13g2_decap_8 FILLER_142_57 ();
 sg13g2_decap_8 FILLER_142_64 ();
 sg13g2_decap_4 FILLER_142_71 ();
 sg13g2_fill_1 FILLER_142_75 ();
 sg13g2_decap_4 FILLER_142_89 ();
 sg13g2_fill_1 FILLER_142_93 ();
 sg13g2_fill_1 FILLER_142_102 ();
 sg13g2_fill_2 FILLER_142_108 ();
 sg13g2_decap_4 FILLER_142_115 ();
 sg13g2_fill_1 FILLER_142_119 ();
 sg13g2_decap_8 FILLER_142_124 ();
 sg13g2_decap_8 FILLER_142_131 ();
 sg13g2_decap_4 FILLER_142_138 ();
 sg13g2_fill_2 FILLER_142_142 ();
 sg13g2_decap_8 FILLER_142_163 ();
 sg13g2_decap_8 FILLER_142_170 ();
 sg13g2_decap_4 FILLER_142_177 ();
 sg13g2_fill_1 FILLER_142_181 ();
 sg13g2_decap_8 FILLER_142_187 ();
 sg13g2_decap_4 FILLER_142_194 ();
 sg13g2_fill_2 FILLER_142_198 ();
 sg13g2_decap_8 FILLER_142_204 ();
 sg13g2_fill_2 FILLER_142_211 ();
 sg13g2_decap_8 FILLER_142_221 ();
 sg13g2_decap_4 FILLER_142_228 ();
 sg13g2_decap_8 FILLER_142_237 ();
 sg13g2_decap_8 FILLER_142_244 ();
 sg13g2_decap_8 FILLER_142_251 ();
 sg13g2_decap_8 FILLER_142_258 ();
 sg13g2_fill_1 FILLER_142_265 ();
 sg13g2_fill_2 FILLER_142_283 ();
 sg13g2_decap_8 FILLER_142_289 ();
 sg13g2_decap_8 FILLER_142_336 ();
 sg13g2_decap_8 FILLER_142_343 ();
 sg13g2_decap_8 FILLER_142_350 ();
 sg13g2_decap_8 FILLER_142_357 ();
 sg13g2_fill_2 FILLER_142_364 ();
 sg13g2_fill_1 FILLER_142_366 ();
 sg13g2_decap_8 FILLER_142_380 ();
 sg13g2_decap_8 FILLER_142_387 ();
 sg13g2_decap_8 FILLER_142_394 ();
 sg13g2_decap_8 FILLER_142_401 ();
 sg13g2_decap_8 FILLER_142_408 ();
 sg13g2_decap_8 FILLER_142_432 ();
 sg13g2_decap_8 FILLER_142_439 ();
 sg13g2_decap_8 FILLER_142_446 ();
 sg13g2_decap_8 FILLER_142_453 ();
 sg13g2_decap_8 FILLER_142_460 ();
 sg13g2_decap_8 FILLER_142_480 ();
 sg13g2_decap_8 FILLER_142_487 ();
 sg13g2_decap_8 FILLER_142_494 ();
 sg13g2_decap_8 FILLER_142_501 ();
 sg13g2_decap_8 FILLER_142_508 ();
 sg13g2_decap_8 FILLER_142_515 ();
 sg13g2_decap_8 FILLER_142_522 ();
 sg13g2_decap_8 FILLER_142_529 ();
 sg13g2_decap_8 FILLER_142_536 ();
 sg13g2_decap_8 FILLER_142_543 ();
 sg13g2_fill_2 FILLER_142_550 ();
 sg13g2_decap_8 FILLER_142_556 ();
 sg13g2_decap_8 FILLER_142_563 ();
 sg13g2_decap_8 FILLER_142_570 ();
 sg13g2_decap_8 FILLER_142_577 ();
 sg13g2_decap_4 FILLER_142_584 ();
 sg13g2_fill_2 FILLER_142_588 ();
 sg13g2_decap_8 FILLER_142_593 ();
 sg13g2_decap_8 FILLER_142_600 ();
 sg13g2_decap_8 FILLER_142_607 ();
 sg13g2_decap_8 FILLER_142_661 ();
 sg13g2_decap_8 FILLER_142_668 ();
 sg13g2_fill_2 FILLER_142_675 ();
 sg13g2_fill_1 FILLER_142_677 ();
 sg13g2_decap_8 FILLER_142_698 ();
 sg13g2_decap_8 FILLER_142_705 ();
 sg13g2_fill_1 FILLER_142_712 ();
 sg13g2_decap_4 FILLER_142_722 ();
 sg13g2_decap_8 FILLER_142_730 ();
 sg13g2_decap_8 FILLER_142_737 ();
 sg13g2_decap_8 FILLER_142_744 ();
 sg13g2_decap_8 FILLER_142_751 ();
 sg13g2_decap_4 FILLER_142_758 ();
 sg13g2_fill_2 FILLER_142_762 ();
 sg13g2_decap_8 FILLER_142_767 ();
 sg13g2_decap_8 FILLER_142_774 ();
 sg13g2_decap_8 FILLER_142_781 ();
 sg13g2_decap_8 FILLER_142_788 ();
 sg13g2_decap_8 FILLER_142_795 ();
 sg13g2_decap_8 FILLER_142_802 ();
 sg13g2_fill_2 FILLER_142_809 ();
 sg13g2_fill_1 FILLER_142_811 ();
 sg13g2_decap_8 FILLER_142_833 ();
 sg13g2_decap_8 FILLER_142_840 ();
 sg13g2_decap_4 FILLER_142_847 ();
 sg13g2_fill_2 FILLER_142_851 ();
 sg13g2_fill_2 FILLER_142_873 ();
 sg13g2_fill_1 FILLER_142_875 ();
 sg13g2_decap_8 FILLER_142_884 ();
 sg13g2_fill_1 FILLER_142_891 ();
 sg13g2_fill_2 FILLER_142_931 ();
 sg13g2_fill_1 FILLER_142_933 ();
 sg13g2_decap_8 FILLER_142_942 ();
 sg13g2_decap_8 FILLER_142_949 ();
 sg13g2_decap_4 FILLER_142_956 ();
 sg13g2_fill_2 FILLER_142_960 ();
 sg13g2_decap_8 FILLER_142_966 ();
 sg13g2_decap_8 FILLER_142_973 ();
 sg13g2_decap_8 FILLER_142_980 ();
 sg13g2_decap_8 FILLER_142_987 ();
 sg13g2_fill_1 FILLER_142_994 ();
 sg13g2_decap_8 FILLER_142_1003 ();
 sg13g2_decap_8 FILLER_142_1010 ();
 sg13g2_decap_8 FILLER_142_1017 ();
 sg13g2_decap_8 FILLER_142_1024 ();
 sg13g2_decap_8 FILLER_142_1031 ();
 sg13g2_fill_1 FILLER_142_1038 ();
 sg13g2_decap_8 FILLER_142_1047 ();
 sg13g2_decap_8 FILLER_142_1054 ();
 sg13g2_fill_1 FILLER_142_1061 ();
 sg13g2_fill_1 FILLER_142_1070 ();
 sg13g2_decap_8 FILLER_142_1083 ();
 sg13g2_decap_4 FILLER_142_1090 ();
 sg13g2_decap_8 FILLER_142_1116 ();
 sg13g2_decap_4 FILLER_142_1123 ();
 sg13g2_fill_1 FILLER_142_1127 ();
 sg13g2_decap_8 FILLER_142_1136 ();
 sg13g2_decap_4 FILLER_142_1143 ();
 sg13g2_fill_2 FILLER_142_1147 ();
 sg13g2_decap_8 FILLER_142_1175 ();
 sg13g2_decap_8 FILLER_142_1182 ();
 sg13g2_decap_8 FILLER_142_1189 ();
 sg13g2_fill_2 FILLER_142_1196 ();
 sg13g2_fill_1 FILLER_142_1198 ();
 sg13g2_decap_4 FILLER_142_1215 ();
 sg13g2_decap_4 FILLER_142_1228 ();
 sg13g2_fill_2 FILLER_142_1232 ();
 sg13g2_decap_8 FILLER_142_1242 ();
 sg13g2_decap_8 FILLER_142_1249 ();
 sg13g2_decap_8 FILLER_142_1256 ();
 sg13g2_decap_8 FILLER_142_1263 ();
 sg13g2_decap_4 FILLER_142_1270 ();
 sg13g2_decap_8 FILLER_142_1278 ();
 sg13g2_decap_8 FILLER_142_1289 ();
 sg13g2_decap_8 FILLER_142_1296 ();
 sg13g2_decap_4 FILLER_142_1303 ();
 sg13g2_fill_1 FILLER_142_1307 ();
 sg13g2_decap_8 FILLER_142_1315 ();
 sg13g2_decap_8 FILLER_142_1322 ();
 sg13g2_fill_2 FILLER_142_1329 ();
 sg13g2_decap_8 FILLER_142_1341 ();
 sg13g2_decap_8 FILLER_142_1348 ();
 sg13g2_fill_2 FILLER_142_1355 ();
 sg13g2_decap_8 FILLER_142_1365 ();
 sg13g2_fill_2 FILLER_142_1372 ();
 sg13g2_fill_1 FILLER_142_1374 ();
 sg13g2_decap_8 FILLER_142_1379 ();
 sg13g2_decap_8 FILLER_142_1386 ();
 sg13g2_decap_8 FILLER_142_1393 ();
 sg13g2_decap_8 FILLER_142_1400 ();
 sg13g2_decap_8 FILLER_142_1407 ();
 sg13g2_decap_8 FILLER_142_1414 ();
 sg13g2_decap_8 FILLER_142_1421 ();
 sg13g2_fill_1 FILLER_142_1428 ();
 sg13g2_fill_2 FILLER_142_1434 ();
 sg13g2_fill_1 FILLER_142_1436 ();
 sg13g2_decap_8 FILLER_142_1442 ();
 sg13g2_decap_8 FILLER_142_1449 ();
 sg13g2_decap_4 FILLER_142_1456 ();
 sg13g2_fill_2 FILLER_142_1460 ();
 sg13g2_fill_1 FILLER_142_1469 ();
 sg13g2_decap_4 FILLER_142_1478 ();
 sg13g2_fill_1 FILLER_142_1482 ();
 sg13g2_fill_2 FILLER_142_1491 ();
 sg13g2_decap_8 FILLER_142_1503 ();
 sg13g2_decap_4 FILLER_142_1510 ();
 sg13g2_fill_1 FILLER_142_1518 ();
 sg13g2_decap_8 FILLER_142_1527 ();
 sg13g2_decap_8 FILLER_142_1534 ();
 sg13g2_decap_8 FILLER_142_1541 ();
 sg13g2_decap_8 FILLER_142_1548 ();
 sg13g2_decap_8 FILLER_142_1555 ();
 sg13g2_fill_1 FILLER_142_1562 ();
 sg13g2_decap_8 FILLER_142_1591 ();
 sg13g2_decap_8 FILLER_142_1598 ();
 sg13g2_fill_1 FILLER_142_1605 ();
 sg13g2_decap_8 FILLER_142_1645 ();
 sg13g2_decap_8 FILLER_142_1652 ();
 sg13g2_decap_8 FILLER_142_1675 ();
 sg13g2_decap_8 FILLER_142_1682 ();
 sg13g2_decap_8 FILLER_142_1689 ();
 sg13g2_decap_8 FILLER_142_1696 ();
 sg13g2_decap_8 FILLER_142_1703 ();
 sg13g2_decap_8 FILLER_142_1710 ();
 sg13g2_decap_8 FILLER_142_1717 ();
 sg13g2_decap_8 FILLER_142_1724 ();
 sg13g2_decap_8 FILLER_142_1731 ();
 sg13g2_decap_8 FILLER_142_1738 ();
 sg13g2_decap_8 FILLER_142_1745 ();
 sg13g2_decap_8 FILLER_142_1752 ();
 sg13g2_decap_8 FILLER_142_1759 ();
 sg13g2_fill_2 FILLER_142_1766 ();
 sg13g2_decap_8 FILLER_143_0 ();
 sg13g2_decap_8 FILLER_143_7 ();
 sg13g2_decap_8 FILLER_143_14 ();
 sg13g2_decap_8 FILLER_143_21 ();
 sg13g2_decap_8 FILLER_143_28 ();
 sg13g2_fill_1 FILLER_143_35 ();
 sg13g2_decap_4 FILLER_143_44 ();
 sg13g2_decap_8 FILLER_143_52 ();
 sg13g2_decap_8 FILLER_143_59 ();
 sg13g2_decap_8 FILLER_143_66 ();
 sg13g2_decap_8 FILLER_143_73 ();
 sg13g2_decap_8 FILLER_143_80 ();
 sg13g2_decap_8 FILLER_143_87 ();
 sg13g2_decap_4 FILLER_143_94 ();
 sg13g2_fill_1 FILLER_143_98 ();
 sg13g2_decap_8 FILLER_143_104 ();
 sg13g2_decap_8 FILLER_143_111 ();
 sg13g2_decap_8 FILLER_143_118 ();
 sg13g2_decap_8 FILLER_143_125 ();
 sg13g2_fill_2 FILLER_143_132 ();
 sg13g2_fill_1 FILLER_143_134 ();
 sg13g2_fill_2 FILLER_143_139 ();
 sg13g2_fill_1 FILLER_143_141 ();
 sg13g2_decap_8 FILLER_143_160 ();
 sg13g2_decap_8 FILLER_143_167 ();
 sg13g2_fill_2 FILLER_143_174 ();
 sg13g2_fill_1 FILLER_143_176 ();
 sg13g2_decap_8 FILLER_143_190 ();
 sg13g2_decap_8 FILLER_143_197 ();
 sg13g2_decap_8 FILLER_143_204 ();
 sg13g2_decap_8 FILLER_143_211 ();
 sg13g2_decap_8 FILLER_143_222 ();
 sg13g2_decap_8 FILLER_143_229 ();
 sg13g2_decap_8 FILLER_143_236 ();
 sg13g2_decap_8 FILLER_143_243 ();
 sg13g2_decap_8 FILLER_143_250 ();
 sg13g2_fill_2 FILLER_143_257 ();
 sg13g2_fill_1 FILLER_143_267 ();
 sg13g2_decap_8 FILLER_143_289 ();
 sg13g2_decap_8 FILLER_143_296 ();
 sg13g2_decap_8 FILLER_143_303 ();
 sg13g2_decap_4 FILLER_143_310 ();
 sg13g2_fill_1 FILLER_143_314 ();
 sg13g2_decap_8 FILLER_143_328 ();
 sg13g2_decap_8 FILLER_143_335 ();
 sg13g2_decap_8 FILLER_143_342 ();
 sg13g2_decap_8 FILLER_143_349 ();
 sg13g2_decap_8 FILLER_143_356 ();
 sg13g2_decap_8 FILLER_143_363 ();
 sg13g2_decap_8 FILLER_143_370 ();
 sg13g2_decap_8 FILLER_143_377 ();
 sg13g2_decap_4 FILLER_143_384 ();
 sg13g2_fill_1 FILLER_143_388 ();
 sg13g2_decap_8 FILLER_143_405 ();
 sg13g2_decap_4 FILLER_143_412 ();
 sg13g2_decap_8 FILLER_143_432 ();
 sg13g2_decap_8 FILLER_143_439 ();
 sg13g2_decap_8 FILLER_143_454 ();
 sg13g2_decap_8 FILLER_143_461 ();
 sg13g2_fill_2 FILLER_143_468 ();
 sg13g2_fill_1 FILLER_143_470 ();
 sg13g2_fill_2 FILLER_143_479 ();
 sg13g2_fill_1 FILLER_143_481 ();
 sg13g2_fill_1 FILLER_143_485 ();
 sg13g2_decap_8 FILLER_143_490 ();
 sg13g2_decap_8 FILLER_143_497 ();
 sg13g2_decap_8 FILLER_143_504 ();
 sg13g2_decap_8 FILLER_143_511 ();
 sg13g2_decap_8 FILLER_143_518 ();
 sg13g2_fill_2 FILLER_143_525 ();
 sg13g2_decap_8 FILLER_143_536 ();
 sg13g2_decap_4 FILLER_143_543 ();
 sg13g2_fill_1 FILLER_143_547 ();
 sg13g2_decap_8 FILLER_143_557 ();
 sg13g2_decap_8 FILLER_143_564 ();
 sg13g2_decap_4 FILLER_143_571 ();
 sg13g2_fill_2 FILLER_143_575 ();
 sg13g2_decap_8 FILLER_143_603 ();
 sg13g2_decap_8 FILLER_143_610 ();
 sg13g2_decap_8 FILLER_143_617 ();
 sg13g2_decap_8 FILLER_143_624 ();
 sg13g2_decap_8 FILLER_143_631 ();
 sg13g2_decap_8 FILLER_143_638 ();
 sg13g2_decap_8 FILLER_143_645 ();
 sg13g2_decap_8 FILLER_143_652 ();
 sg13g2_decap_8 FILLER_143_659 ();
 sg13g2_decap_4 FILLER_143_666 ();
 sg13g2_fill_1 FILLER_143_670 ();
 sg13g2_decap_8 FILLER_143_675 ();
 sg13g2_fill_2 FILLER_143_682 ();
 sg13g2_fill_1 FILLER_143_684 ();
 sg13g2_decap_8 FILLER_143_689 ();
 sg13g2_decap_8 FILLER_143_696 ();
 sg13g2_decap_8 FILLER_143_703 ();
 sg13g2_decap_4 FILLER_143_710 ();
 sg13g2_fill_2 FILLER_143_714 ();
 sg13g2_decap_4 FILLER_143_719 ();
 sg13g2_fill_2 FILLER_143_723 ();
 sg13g2_decap_8 FILLER_143_737 ();
 sg13g2_decap_8 FILLER_143_744 ();
 sg13g2_decap_8 FILLER_143_751 ();
 sg13g2_fill_2 FILLER_143_770 ();
 sg13g2_decap_8 FILLER_143_784 ();
 sg13g2_decap_8 FILLER_143_791 ();
 sg13g2_decap_8 FILLER_143_798 ();
 sg13g2_fill_2 FILLER_143_805 ();
 sg13g2_fill_1 FILLER_143_807 ();
 sg13g2_decap_4 FILLER_143_816 ();
 sg13g2_decap_8 FILLER_143_828 ();
 sg13g2_decap_8 FILLER_143_835 ();
 sg13g2_decap_8 FILLER_143_842 ();
 sg13g2_fill_2 FILLER_143_849 ();
 sg13g2_decap_8 FILLER_143_857 ();
 sg13g2_decap_8 FILLER_143_864 ();
 sg13g2_decap_8 FILLER_143_871 ();
 sg13g2_fill_2 FILLER_143_878 ();
 sg13g2_decap_8 FILLER_143_883 ();
 sg13g2_decap_8 FILLER_143_890 ();
 sg13g2_decap_4 FILLER_143_897 ();
 sg13g2_fill_2 FILLER_143_901 ();
 sg13g2_decap_8 FILLER_143_907 ();
 sg13g2_decap_8 FILLER_143_914 ();
 sg13g2_decap_8 FILLER_143_921 ();
 sg13g2_decap_8 FILLER_143_928 ();
 sg13g2_decap_8 FILLER_143_935 ();
 sg13g2_decap_8 FILLER_143_942 ();
 sg13g2_decap_8 FILLER_143_949 ();
 sg13g2_fill_2 FILLER_143_956 ();
 sg13g2_decap_8 FILLER_143_961 ();
 sg13g2_decap_8 FILLER_143_968 ();
 sg13g2_decap_8 FILLER_143_975 ();
 sg13g2_fill_2 FILLER_143_982 ();
 sg13g2_decap_8 FILLER_143_1002 ();
 sg13g2_decap_8 FILLER_143_1009 ();
 sg13g2_decap_8 FILLER_143_1016 ();
 sg13g2_decap_8 FILLER_143_1023 ();
 sg13g2_decap_8 FILLER_143_1030 ();
 sg13g2_decap_8 FILLER_143_1037 ();
 sg13g2_decap_8 FILLER_143_1044 ();
 sg13g2_decap_8 FILLER_143_1051 ();
 sg13g2_decap_8 FILLER_143_1058 ();
 sg13g2_decap_4 FILLER_143_1065 ();
 sg13g2_fill_1 FILLER_143_1069 ();
 sg13g2_decap_8 FILLER_143_1078 ();
 sg13g2_decap_8 FILLER_143_1085 ();
 sg13g2_decap_8 FILLER_143_1092 ();
 sg13g2_fill_2 FILLER_143_1099 ();
 sg13g2_decap_8 FILLER_143_1118 ();
 sg13g2_decap_8 FILLER_143_1125 ();
 sg13g2_decap_8 FILLER_143_1132 ();
 sg13g2_decap_8 FILLER_143_1139 ();
 sg13g2_decap_8 FILLER_143_1146 ();
 sg13g2_fill_2 FILLER_143_1153 ();
 sg13g2_decap_8 FILLER_143_1161 ();
 sg13g2_decap_4 FILLER_143_1168 ();
 sg13g2_decap_4 FILLER_143_1177 ();
 sg13g2_decap_8 FILLER_143_1185 ();
 sg13g2_decap_8 FILLER_143_1192 ();
 sg13g2_decap_8 FILLER_143_1199 ();
 sg13g2_fill_2 FILLER_143_1222 ();
 sg13g2_decap_8 FILLER_143_1232 ();
 sg13g2_decap_8 FILLER_143_1239 ();
 sg13g2_decap_8 FILLER_143_1246 ();
 sg13g2_decap_8 FILLER_143_1253 ();
 sg13g2_decap_8 FILLER_143_1260 ();
 sg13g2_fill_2 FILLER_143_1267 ();
 sg13g2_fill_2 FILLER_143_1281 ();
 sg13g2_fill_1 FILLER_143_1283 ();
 sg13g2_decap_8 FILLER_143_1289 ();
 sg13g2_decap_8 FILLER_143_1296 ();
 sg13g2_decap_4 FILLER_143_1303 ();
 sg13g2_fill_1 FILLER_143_1307 ();
 sg13g2_fill_2 FILLER_143_1314 ();
 sg13g2_fill_1 FILLER_143_1316 ();
 sg13g2_decap_8 FILLER_143_1321 ();
 sg13g2_decap_8 FILLER_143_1328 ();
 sg13g2_decap_8 FILLER_143_1335 ();
 sg13g2_decap_8 FILLER_143_1342 ();
 sg13g2_decap_8 FILLER_143_1349 ();
 sg13g2_decap_8 FILLER_143_1356 ();
 sg13g2_decap_4 FILLER_143_1363 ();
 sg13g2_decap_8 FILLER_143_1387 ();
 sg13g2_decap_8 FILLER_143_1394 ();
 sg13g2_decap_8 FILLER_143_1401 ();
 sg13g2_decap_8 FILLER_143_1408 ();
 sg13g2_decap_4 FILLER_143_1415 ();
 sg13g2_fill_1 FILLER_143_1419 ();
 sg13g2_decap_4 FILLER_143_1425 ();
 sg13g2_fill_1 FILLER_143_1429 ();
 sg13g2_decap_8 FILLER_143_1438 ();
 sg13g2_fill_2 FILLER_143_1445 ();
 sg13g2_decap_8 FILLER_143_1451 ();
 sg13g2_fill_1 FILLER_143_1458 ();
 sg13g2_decap_8 FILLER_143_1475 ();
 sg13g2_decap_8 FILLER_143_1482 ();
 sg13g2_decap_8 FILLER_143_1489 ();
 sg13g2_decap_4 FILLER_143_1496 ();
 sg13g2_fill_2 FILLER_143_1500 ();
 sg13g2_decap_8 FILLER_143_1510 ();
 sg13g2_decap_8 FILLER_143_1517 ();
 sg13g2_decap_8 FILLER_143_1524 ();
 sg13g2_decap_8 FILLER_143_1531 ();
 sg13g2_decap_8 FILLER_143_1538 ();
 sg13g2_decap_8 FILLER_143_1545 ();
 sg13g2_decap_8 FILLER_143_1552 ();
 sg13g2_decap_8 FILLER_143_1559 ();
 sg13g2_decap_4 FILLER_143_1566 ();
 sg13g2_decap_8 FILLER_143_1586 ();
 sg13g2_decap_8 FILLER_143_1593 ();
 sg13g2_decap_8 FILLER_143_1600 ();
 sg13g2_decap_8 FILLER_143_1607 ();
 sg13g2_fill_2 FILLER_143_1614 ();
 sg13g2_decap_8 FILLER_143_1620 ();
 sg13g2_decap_8 FILLER_143_1627 ();
 sg13g2_decap_8 FILLER_143_1634 ();
 sg13g2_decap_8 FILLER_143_1641 ();
 sg13g2_decap_8 FILLER_143_1648 ();
 sg13g2_decap_8 FILLER_143_1675 ();
 sg13g2_decap_8 FILLER_143_1682 ();
 sg13g2_decap_8 FILLER_143_1689 ();
 sg13g2_decap_8 FILLER_143_1696 ();
 sg13g2_decap_8 FILLER_143_1703 ();
 sg13g2_decap_8 FILLER_143_1710 ();
 sg13g2_decap_8 FILLER_143_1717 ();
 sg13g2_decap_8 FILLER_143_1724 ();
 sg13g2_decap_8 FILLER_143_1731 ();
 sg13g2_decap_8 FILLER_143_1738 ();
 sg13g2_decap_8 FILLER_143_1745 ();
 sg13g2_decap_8 FILLER_143_1752 ();
 sg13g2_decap_8 FILLER_143_1759 ();
 sg13g2_fill_2 FILLER_143_1766 ();
 sg13g2_decap_8 FILLER_144_0 ();
 sg13g2_decap_8 FILLER_144_7 ();
 sg13g2_fill_2 FILLER_144_14 ();
 sg13g2_fill_1 FILLER_144_16 ();
 sg13g2_decap_8 FILLER_144_33 ();
 sg13g2_decap_8 FILLER_144_40 ();
 sg13g2_decap_8 FILLER_144_47 ();
 sg13g2_decap_8 FILLER_144_54 ();
 sg13g2_decap_8 FILLER_144_61 ();
 sg13g2_decap_8 FILLER_144_68 ();
 sg13g2_decap_8 FILLER_144_75 ();
 sg13g2_decap_8 FILLER_144_82 ();
 sg13g2_decap_8 FILLER_144_89 ();
 sg13g2_decap_4 FILLER_144_96 ();
 sg13g2_fill_1 FILLER_144_100 ();
 sg13g2_decap_8 FILLER_144_105 ();
 sg13g2_decap_8 FILLER_144_112 ();
 sg13g2_decap_8 FILLER_144_119 ();
 sg13g2_fill_2 FILLER_144_126 ();
 sg13g2_fill_1 FILLER_144_128 ();
 sg13g2_decap_8 FILLER_144_142 ();
 sg13g2_decap_8 FILLER_144_149 ();
 sg13g2_decap_8 FILLER_144_156 ();
 sg13g2_fill_2 FILLER_144_163 ();
 sg13g2_decap_8 FILLER_144_173 ();
 sg13g2_decap_8 FILLER_144_180 ();
 sg13g2_decap_8 FILLER_144_187 ();
 sg13g2_decap_8 FILLER_144_194 ();
 sg13g2_decap_8 FILLER_144_201 ();
 sg13g2_decap_8 FILLER_144_208 ();
 sg13g2_fill_1 FILLER_144_215 ();
 sg13g2_decap_8 FILLER_144_224 ();
 sg13g2_decap_8 FILLER_144_231 ();
 sg13g2_decap_8 FILLER_144_238 ();
 sg13g2_decap_8 FILLER_144_245 ();
 sg13g2_decap_4 FILLER_144_252 ();
 sg13g2_decap_8 FILLER_144_282 ();
 sg13g2_decap_8 FILLER_144_289 ();
 sg13g2_decap_8 FILLER_144_296 ();
 sg13g2_decap_8 FILLER_144_303 ();
 sg13g2_fill_1 FILLER_144_310 ();
 sg13g2_decap_8 FILLER_144_324 ();
 sg13g2_decap_4 FILLER_144_331 ();
 sg13g2_fill_1 FILLER_144_335 ();
 sg13g2_decap_8 FILLER_144_349 ();
 sg13g2_fill_2 FILLER_144_356 ();
 sg13g2_fill_1 FILLER_144_358 ();
 sg13g2_decap_8 FILLER_144_372 ();
 sg13g2_decap_8 FILLER_144_379 ();
 sg13g2_decap_8 FILLER_144_386 ();
 sg13g2_decap_8 FILLER_144_393 ();
 sg13g2_decap_8 FILLER_144_408 ();
 sg13g2_decap_8 FILLER_144_415 ();
 sg13g2_decap_8 FILLER_144_430 ();
 sg13g2_decap_8 FILLER_144_437 ();
 sg13g2_decap_8 FILLER_144_444 ();
 sg13g2_fill_2 FILLER_144_451 ();
 sg13g2_decap_8 FILLER_144_468 ();
 sg13g2_decap_4 FILLER_144_475 ();
 sg13g2_fill_2 FILLER_144_479 ();
 sg13g2_decap_8 FILLER_144_498 ();
 sg13g2_fill_1 FILLER_144_505 ();
 sg13g2_fill_2 FILLER_144_517 ();
 sg13g2_decap_8 FILLER_144_527 ();
 sg13g2_decap_8 FILLER_144_534 ();
 sg13g2_decap_8 FILLER_144_562 ();
 sg13g2_fill_2 FILLER_144_569 ();
 sg13g2_decap_8 FILLER_144_575 ();
 sg13g2_decap_8 FILLER_144_582 ();
 sg13g2_decap_8 FILLER_144_589 ();
 sg13g2_decap_8 FILLER_144_596 ();
 sg13g2_decap_8 FILLER_144_603 ();
 sg13g2_decap_8 FILLER_144_610 ();
 sg13g2_decap_8 FILLER_144_629 ();
 sg13g2_decap_8 FILLER_144_636 ();
 sg13g2_decap_8 FILLER_144_643 ();
 sg13g2_decap_4 FILLER_144_650 ();
 sg13g2_decap_8 FILLER_144_662 ();
 sg13g2_decap_8 FILLER_144_669 ();
 sg13g2_decap_8 FILLER_144_676 ();
 sg13g2_decap_8 FILLER_144_683 ();
 sg13g2_decap_8 FILLER_144_690 ();
 sg13g2_decap_8 FILLER_144_746 ();
 sg13g2_decap_8 FILLER_144_753 ();
 sg13g2_fill_1 FILLER_144_776 ();
 sg13g2_decap_8 FILLER_144_786 ();
 sg13g2_decap_8 FILLER_144_793 ();
 sg13g2_decap_4 FILLER_144_800 ();
 sg13g2_fill_1 FILLER_144_804 ();
 sg13g2_decap_8 FILLER_144_813 ();
 sg13g2_decap_8 FILLER_144_820 ();
 sg13g2_fill_1 FILLER_144_827 ();
 sg13g2_decap_8 FILLER_144_845 ();
 sg13g2_decap_8 FILLER_144_852 ();
 sg13g2_decap_8 FILLER_144_859 ();
 sg13g2_decap_8 FILLER_144_866 ();
 sg13g2_decap_8 FILLER_144_873 ();
 sg13g2_decap_8 FILLER_144_888 ();
 sg13g2_decap_8 FILLER_144_895 ();
 sg13g2_decap_8 FILLER_144_902 ();
 sg13g2_decap_8 FILLER_144_909 ();
 sg13g2_decap_8 FILLER_144_916 ();
 sg13g2_decap_8 FILLER_144_923 ();
 sg13g2_decap_8 FILLER_144_930 ();
 sg13g2_decap_8 FILLER_144_937 ();
 sg13g2_decap_4 FILLER_144_944 ();
 sg13g2_fill_2 FILLER_144_948 ();
 sg13g2_decap_8 FILLER_144_962 ();
 sg13g2_decap_8 FILLER_144_974 ();
 sg13g2_decap_8 FILLER_144_981 ();
 sg13g2_fill_2 FILLER_144_988 ();
 sg13g2_decap_4 FILLER_144_1009 ();
 sg13g2_decap_8 FILLER_144_1021 ();
 sg13g2_decap_8 FILLER_144_1028 ();
 sg13g2_decap_8 FILLER_144_1035 ();
 sg13g2_decap_8 FILLER_144_1042 ();
 sg13g2_decap_8 FILLER_144_1049 ();
 sg13g2_decap_8 FILLER_144_1056 ();
 sg13g2_decap_8 FILLER_144_1063 ();
 sg13g2_decap_8 FILLER_144_1070 ();
 sg13g2_decap_8 FILLER_144_1077 ();
 sg13g2_fill_1 FILLER_144_1089 ();
 sg13g2_decap_4 FILLER_144_1095 ();
 sg13g2_fill_1 FILLER_144_1099 ();
 sg13g2_decap_8 FILLER_144_1108 ();
 sg13g2_decap_8 FILLER_144_1119 ();
 sg13g2_fill_2 FILLER_144_1126 ();
 sg13g2_decap_4 FILLER_144_1132 ();
 sg13g2_fill_2 FILLER_144_1141 ();
 sg13g2_fill_1 FILLER_144_1143 ();
 sg13g2_decap_8 FILLER_144_1160 ();
 sg13g2_decap_8 FILLER_144_1167 ();
 sg13g2_decap_8 FILLER_144_1174 ();
 sg13g2_decap_8 FILLER_144_1197 ();
 sg13g2_decap_8 FILLER_144_1204 ();
 sg13g2_decap_8 FILLER_144_1211 ();
 sg13g2_fill_1 FILLER_144_1218 ();
 sg13g2_fill_1 FILLER_144_1224 ();
 sg13g2_decap_8 FILLER_144_1238 ();
 sg13g2_decap_8 FILLER_144_1245 ();
 sg13g2_decap_8 FILLER_144_1252 ();
 sg13g2_decap_8 FILLER_144_1259 ();
 sg13g2_fill_2 FILLER_144_1266 ();
 sg13g2_fill_1 FILLER_144_1268 ();
 sg13g2_decap_4 FILLER_144_1278 ();
 sg13g2_decap_8 FILLER_144_1298 ();
 sg13g2_decap_8 FILLER_144_1336 ();
 sg13g2_decap_8 FILLER_144_1353 ();
 sg13g2_decap_8 FILLER_144_1360 ();
 sg13g2_fill_2 FILLER_144_1367 ();
 sg13g2_fill_1 FILLER_144_1369 ();
 sg13g2_decap_8 FILLER_144_1378 ();
 sg13g2_decap_8 FILLER_144_1391 ();
 sg13g2_decap_8 FILLER_144_1398 ();
 sg13g2_decap_8 FILLER_144_1405 ();
 sg13g2_fill_2 FILLER_144_1412 ();
 sg13g2_fill_1 FILLER_144_1414 ();
 sg13g2_decap_8 FILLER_144_1426 ();
 sg13g2_decap_8 FILLER_144_1433 ();
 sg13g2_decap_8 FILLER_144_1440 ();
 sg13g2_decap_8 FILLER_144_1447 ();
 sg13g2_decap_8 FILLER_144_1454 ();
 sg13g2_decap_8 FILLER_144_1461 ();
 sg13g2_decap_8 FILLER_144_1468 ();
 sg13g2_decap_8 FILLER_144_1475 ();
 sg13g2_decap_8 FILLER_144_1482 ();
 sg13g2_decap_8 FILLER_144_1489 ();
 sg13g2_decap_8 FILLER_144_1496 ();
 sg13g2_decap_8 FILLER_144_1503 ();
 sg13g2_fill_2 FILLER_144_1510 ();
 sg13g2_decap_8 FILLER_144_1515 ();
 sg13g2_decap_8 FILLER_144_1522 ();
 sg13g2_decap_8 FILLER_144_1529 ();
 sg13g2_fill_2 FILLER_144_1536 ();
 sg13g2_fill_1 FILLER_144_1538 ();
 sg13g2_decap_8 FILLER_144_1555 ();
 sg13g2_decap_8 FILLER_144_1562 ();
 sg13g2_decap_4 FILLER_144_1569 ();
 sg13g2_fill_1 FILLER_144_1573 ();
 sg13g2_decap_8 FILLER_144_1579 ();
 sg13g2_decap_8 FILLER_144_1586 ();
 sg13g2_decap_8 FILLER_144_1593 ();
 sg13g2_decap_8 FILLER_144_1600 ();
 sg13g2_decap_8 FILLER_144_1607 ();
 sg13g2_decap_8 FILLER_144_1614 ();
 sg13g2_decap_8 FILLER_144_1621 ();
 sg13g2_decap_8 FILLER_144_1628 ();
 sg13g2_decap_8 FILLER_144_1635 ();
 sg13g2_fill_1 FILLER_144_1642 ();
 sg13g2_fill_1 FILLER_144_1659 ();
 sg13g2_decap_8 FILLER_144_1670 ();
 sg13g2_decap_8 FILLER_144_1677 ();
 sg13g2_decap_8 FILLER_144_1684 ();
 sg13g2_decap_8 FILLER_144_1691 ();
 sg13g2_decap_8 FILLER_144_1698 ();
 sg13g2_decap_8 FILLER_144_1705 ();
 sg13g2_decap_8 FILLER_144_1712 ();
 sg13g2_decap_8 FILLER_144_1719 ();
 sg13g2_decap_8 FILLER_144_1726 ();
 sg13g2_decap_8 FILLER_144_1733 ();
 sg13g2_decap_8 FILLER_144_1740 ();
 sg13g2_decap_8 FILLER_144_1747 ();
 sg13g2_decap_8 FILLER_144_1754 ();
 sg13g2_decap_8 FILLER_144_1761 ();
 sg13g2_decap_8 FILLER_145_0 ();
 sg13g2_decap_8 FILLER_145_7 ();
 sg13g2_fill_2 FILLER_145_14 ();
 sg13g2_fill_2 FILLER_145_24 ();
 sg13g2_fill_1 FILLER_145_26 ();
 sg13g2_fill_1 FILLER_145_32 ();
 sg13g2_decap_4 FILLER_145_36 ();
 sg13g2_fill_2 FILLER_145_40 ();
 sg13g2_decap_8 FILLER_145_47 ();
 sg13g2_decap_8 FILLER_145_54 ();
 sg13g2_decap_8 FILLER_145_61 ();
 sg13g2_decap_8 FILLER_145_68 ();
 sg13g2_fill_2 FILLER_145_75 ();
 sg13g2_decap_4 FILLER_145_85 ();
 sg13g2_fill_1 FILLER_145_89 ();
 sg13g2_fill_1 FILLER_145_98 ();
 sg13g2_fill_1 FILLER_145_103 ();
 sg13g2_fill_1 FILLER_145_109 ();
 sg13g2_decap_8 FILLER_145_114 ();
 sg13g2_decap_8 FILLER_145_121 ();
 sg13g2_decap_8 FILLER_145_128 ();
 sg13g2_decap_8 FILLER_145_135 ();
 sg13g2_fill_2 FILLER_145_142 ();
 sg13g2_fill_1 FILLER_145_144 ();
 sg13g2_fill_1 FILLER_145_157 ();
 sg13g2_decap_8 FILLER_145_182 ();
 sg13g2_decap_8 FILLER_145_189 ();
 sg13g2_decap_8 FILLER_145_196 ();
 sg13g2_fill_2 FILLER_145_203 ();
 sg13g2_fill_1 FILLER_145_205 ();
 sg13g2_decap_8 FILLER_145_210 ();
 sg13g2_decap_8 FILLER_145_217 ();
 sg13g2_fill_2 FILLER_145_224 ();
 sg13g2_fill_1 FILLER_145_226 ();
 sg13g2_decap_8 FILLER_145_235 ();
 sg13g2_decap_8 FILLER_145_242 ();
 sg13g2_decap_8 FILLER_145_249 ();
 sg13g2_decap_8 FILLER_145_256 ();
 sg13g2_decap_8 FILLER_145_263 ();
 sg13g2_decap_8 FILLER_145_270 ();
 sg13g2_decap_8 FILLER_145_277 ();
 sg13g2_decap_8 FILLER_145_284 ();
 sg13g2_decap_8 FILLER_145_291 ();
 sg13g2_decap_8 FILLER_145_298 ();
 sg13g2_decap_8 FILLER_145_305 ();
 sg13g2_decap_8 FILLER_145_312 ();
 sg13g2_decap_8 FILLER_145_319 ();
 sg13g2_decap_8 FILLER_145_326 ();
 sg13g2_decap_8 FILLER_145_333 ();
 sg13g2_decap_8 FILLER_145_340 ();
 sg13g2_decap_4 FILLER_145_347 ();
 sg13g2_fill_1 FILLER_145_351 ();
 sg13g2_decap_4 FILLER_145_366 ();
 sg13g2_decap_8 FILLER_145_378 ();
 sg13g2_decap_8 FILLER_145_385 ();
 sg13g2_decap_8 FILLER_145_392 ();
 sg13g2_fill_1 FILLER_145_399 ();
 sg13g2_decap_8 FILLER_145_416 ();
 sg13g2_fill_1 FILLER_145_423 ();
 sg13g2_decap_4 FILLER_145_436 ();
 sg13g2_fill_2 FILLER_145_440 ();
 sg13g2_decap_8 FILLER_145_447 ();
 sg13g2_fill_2 FILLER_145_454 ();
 sg13g2_fill_1 FILLER_145_456 ();
 sg13g2_fill_1 FILLER_145_462 ();
 sg13g2_decap_8 FILLER_145_475 ();
 sg13g2_decap_8 FILLER_145_482 ();
 sg13g2_decap_8 FILLER_145_489 ();
 sg13g2_decap_8 FILLER_145_496 ();
 sg13g2_fill_2 FILLER_145_511 ();
 sg13g2_fill_1 FILLER_145_513 ();
 sg13g2_decap_8 FILLER_145_526 ();
 sg13g2_decap_4 FILLER_145_533 ();
 sg13g2_fill_2 FILLER_145_537 ();
 sg13g2_decap_8 FILLER_145_555 ();
 sg13g2_decap_8 FILLER_145_562 ();
 sg13g2_decap_8 FILLER_145_569 ();
 sg13g2_decap_4 FILLER_145_576 ();
 sg13g2_decap_8 FILLER_145_601 ();
 sg13g2_fill_2 FILLER_145_608 ();
 sg13g2_fill_1 FILLER_145_610 ();
 sg13g2_decap_8 FILLER_145_619 ();
 sg13g2_decap_8 FILLER_145_626 ();
 sg13g2_fill_1 FILLER_145_633 ();
 sg13g2_fill_2 FILLER_145_642 ();
 sg13g2_decap_8 FILLER_145_652 ();
 sg13g2_decap_8 FILLER_145_659 ();
 sg13g2_fill_2 FILLER_145_666 ();
 sg13g2_fill_1 FILLER_145_668 ();
 sg13g2_decap_8 FILLER_145_677 ();
 sg13g2_decap_8 FILLER_145_684 ();
 sg13g2_decap_8 FILLER_145_691 ();
 sg13g2_decap_8 FILLER_145_706 ();
 sg13g2_decap_8 FILLER_145_713 ();
 sg13g2_decap_8 FILLER_145_720 ();
 sg13g2_decap_8 FILLER_145_727 ();
 sg13g2_decap_8 FILLER_145_734 ();
 sg13g2_decap_8 FILLER_145_741 ();
 sg13g2_decap_8 FILLER_145_748 ();
 sg13g2_decap_8 FILLER_145_755 ();
 sg13g2_decap_4 FILLER_145_762 ();
 sg13g2_fill_1 FILLER_145_766 ();
 sg13g2_decap_8 FILLER_145_791 ();
 sg13g2_decap_8 FILLER_145_798 ();
 sg13g2_decap_8 FILLER_145_805 ();
 sg13g2_decap_8 FILLER_145_812 ();
 sg13g2_decap_8 FILLER_145_819 ();
 sg13g2_fill_1 FILLER_145_826 ();
 sg13g2_decap_8 FILLER_145_841 ();
 sg13g2_decap_8 FILLER_145_848 ();
 sg13g2_decap_8 FILLER_145_855 ();
 sg13g2_decap_8 FILLER_145_862 ();
 sg13g2_fill_2 FILLER_145_869 ();
 sg13g2_fill_1 FILLER_145_871 ();
 sg13g2_decap_4 FILLER_145_877 ();
 sg13g2_fill_2 FILLER_145_881 ();
 sg13g2_decap_8 FILLER_145_887 ();
 sg13g2_decap_8 FILLER_145_894 ();
 sg13g2_decap_8 FILLER_145_901 ();
 sg13g2_decap_8 FILLER_145_908 ();
 sg13g2_decap_8 FILLER_145_915 ();
 sg13g2_decap_8 FILLER_145_922 ();
 sg13g2_decap_4 FILLER_145_929 ();
 sg13g2_fill_1 FILLER_145_933 ();
 sg13g2_fill_2 FILLER_145_942 ();
 sg13g2_fill_1 FILLER_145_944 ();
 sg13g2_decap_4 FILLER_145_950 ();
 sg13g2_fill_2 FILLER_145_954 ();
 sg13g2_decap_8 FILLER_145_962 ();
 sg13g2_decap_8 FILLER_145_969 ();
 sg13g2_decap_8 FILLER_145_976 ();
 sg13g2_decap_4 FILLER_145_983 ();
 sg13g2_fill_1 FILLER_145_987 ();
 sg13g2_decap_4 FILLER_145_993 ();
 sg13g2_fill_2 FILLER_145_997 ();
 sg13g2_decap_4 FILLER_145_1007 ();
 sg13g2_fill_2 FILLER_145_1011 ();
 sg13g2_decap_8 FILLER_145_1018 ();
 sg13g2_decap_8 FILLER_145_1025 ();
 sg13g2_decap_8 FILLER_145_1032 ();
 sg13g2_decap_8 FILLER_145_1039 ();
 sg13g2_decap_4 FILLER_145_1046 ();
 sg13g2_decap_8 FILLER_145_1064 ();
 sg13g2_decap_8 FILLER_145_1071 ();
 sg13g2_decap_8 FILLER_145_1078 ();
 sg13g2_fill_2 FILLER_145_1085 ();
 sg13g2_fill_2 FILLER_145_1091 ();
 sg13g2_decap_8 FILLER_145_1097 ();
 sg13g2_decap_8 FILLER_145_1104 ();
 sg13g2_decap_8 FILLER_145_1111 ();
 sg13g2_decap_8 FILLER_145_1118 ();
 sg13g2_decap_8 FILLER_145_1125 ();
 sg13g2_decap_8 FILLER_145_1132 ();
 sg13g2_decap_4 FILLER_145_1139 ();
 sg13g2_decap_8 FILLER_145_1157 ();
 sg13g2_fill_2 FILLER_145_1164 ();
 sg13g2_decap_8 FILLER_145_1183 ();
 sg13g2_fill_2 FILLER_145_1190 ();
 sg13g2_decap_8 FILLER_145_1199 ();
 sg13g2_decap_8 FILLER_145_1206 ();
 sg13g2_decap_8 FILLER_145_1213 ();
 sg13g2_decap_8 FILLER_145_1220 ();
 sg13g2_decap_8 FILLER_145_1227 ();
 sg13g2_decap_8 FILLER_145_1234 ();
 sg13g2_decap_8 FILLER_145_1241 ();
 sg13g2_decap_8 FILLER_145_1248 ();
 sg13g2_decap_8 FILLER_145_1255 ();
 sg13g2_decap_4 FILLER_145_1262 ();
 sg13g2_fill_2 FILLER_145_1266 ();
 sg13g2_decap_8 FILLER_145_1281 ();
 sg13g2_decap_8 FILLER_145_1288 ();
 sg13g2_decap_8 FILLER_145_1295 ();
 sg13g2_decap_4 FILLER_145_1302 ();
 sg13g2_fill_2 FILLER_145_1306 ();
 sg13g2_decap_8 FILLER_145_1311 ();
 sg13g2_fill_1 FILLER_145_1318 ();
 sg13g2_fill_2 FILLER_145_1323 ();
 sg13g2_decap_8 FILLER_145_1333 ();
 sg13g2_decap_8 FILLER_145_1360 ();
 sg13g2_decap_8 FILLER_145_1367 ();
 sg13g2_decap_8 FILLER_145_1374 ();
 sg13g2_decap_8 FILLER_145_1381 ();
 sg13g2_fill_2 FILLER_145_1388 ();
 sg13g2_decap_8 FILLER_145_1404 ();
 sg13g2_fill_2 FILLER_145_1411 ();
 sg13g2_decap_8 FILLER_145_1435 ();
 sg13g2_decap_4 FILLER_145_1442 ();
 sg13g2_decap_4 FILLER_145_1454 ();
 sg13g2_fill_2 FILLER_145_1458 ();
 sg13g2_decap_8 FILLER_145_1470 ();
 sg13g2_decap_8 FILLER_145_1477 ();
 sg13g2_decap_8 FILLER_145_1484 ();
 sg13g2_decap_8 FILLER_145_1491 ();
 sg13g2_decap_8 FILLER_145_1498 ();
 sg13g2_decap_4 FILLER_145_1505 ();
 sg13g2_fill_1 FILLER_145_1509 ();
 sg13g2_decap_8 FILLER_145_1531 ();
 sg13g2_decap_8 FILLER_145_1538 ();
 sg13g2_decap_4 FILLER_145_1545 ();
 sg13g2_fill_2 FILLER_145_1554 ();
 sg13g2_fill_1 FILLER_145_1556 ();
 sg13g2_decap_8 FILLER_145_1565 ();
 sg13g2_decap_8 FILLER_145_1572 ();
 sg13g2_decap_8 FILLER_145_1579 ();
 sg13g2_decap_8 FILLER_145_1586 ();
 sg13g2_decap_8 FILLER_145_1593 ();
 sg13g2_decap_8 FILLER_145_1600 ();
 sg13g2_decap_8 FILLER_145_1607 ();
 sg13g2_decap_8 FILLER_145_1614 ();
 sg13g2_decap_8 FILLER_145_1621 ();
 sg13g2_decap_8 FILLER_145_1628 ();
 sg13g2_decap_4 FILLER_145_1635 ();
 sg13g2_fill_1 FILLER_145_1639 ();
 sg13g2_decap_8 FILLER_145_1663 ();
 sg13g2_decap_8 FILLER_145_1670 ();
 sg13g2_decap_8 FILLER_145_1677 ();
 sg13g2_decap_8 FILLER_145_1684 ();
 sg13g2_decap_8 FILLER_145_1691 ();
 sg13g2_decap_8 FILLER_145_1698 ();
 sg13g2_decap_8 FILLER_145_1705 ();
 sg13g2_decap_8 FILLER_145_1712 ();
 sg13g2_decap_8 FILLER_145_1719 ();
 sg13g2_decap_8 FILLER_145_1726 ();
 sg13g2_decap_8 FILLER_145_1733 ();
 sg13g2_decap_8 FILLER_145_1740 ();
 sg13g2_decap_8 FILLER_145_1747 ();
 sg13g2_decap_8 FILLER_145_1754 ();
 sg13g2_decap_8 FILLER_145_1761 ();
 sg13g2_decap_8 FILLER_146_0 ();
 sg13g2_decap_8 FILLER_146_7 ();
 sg13g2_decap_4 FILLER_146_14 ();
 sg13g2_decap_8 FILLER_146_22 ();
 sg13g2_fill_2 FILLER_146_37 ();
 sg13g2_fill_1 FILLER_146_39 ();
 sg13g2_fill_2 FILLER_146_44 ();
 sg13g2_decap_8 FILLER_146_50 ();
 sg13g2_fill_2 FILLER_146_57 ();
 sg13g2_fill_1 FILLER_146_59 ();
 sg13g2_decap_4 FILLER_146_85 ();
 sg13g2_fill_2 FILLER_146_89 ();
 sg13g2_decap_8 FILLER_146_111 ();
 sg13g2_decap_8 FILLER_146_118 ();
 sg13g2_decap_8 FILLER_146_125 ();
 sg13g2_decap_8 FILLER_146_132 ();
 sg13g2_decap_8 FILLER_146_139 ();
 sg13g2_decap_8 FILLER_146_146 ();
 sg13g2_fill_2 FILLER_146_153 ();
 sg13g2_fill_2 FILLER_146_163 ();
 sg13g2_decap_8 FILLER_146_170 ();
 sg13g2_decap_8 FILLER_146_177 ();
 sg13g2_fill_2 FILLER_146_184 ();
 sg13g2_fill_1 FILLER_146_186 ();
 sg13g2_fill_1 FILLER_146_196 ();
 sg13g2_decap_8 FILLER_146_217 ();
 sg13g2_decap_8 FILLER_146_224 ();
 sg13g2_decap_8 FILLER_146_231 ();
 sg13g2_decap_8 FILLER_146_238 ();
 sg13g2_decap_8 FILLER_146_245 ();
 sg13g2_decap_8 FILLER_146_252 ();
 sg13g2_decap_8 FILLER_146_259 ();
 sg13g2_decap_8 FILLER_146_266 ();
 sg13g2_decap_8 FILLER_146_273 ();
 sg13g2_decap_8 FILLER_146_280 ();
 sg13g2_decap_8 FILLER_146_287 ();
 sg13g2_decap_8 FILLER_146_294 ();
 sg13g2_decap_8 FILLER_146_301 ();
 sg13g2_decap_8 FILLER_146_308 ();
 sg13g2_decap_8 FILLER_146_315 ();
 sg13g2_decap_8 FILLER_146_322 ();
 sg13g2_decap_8 FILLER_146_329 ();
 sg13g2_decap_8 FILLER_146_336 ();
 sg13g2_decap_8 FILLER_146_343 ();
 sg13g2_decap_8 FILLER_146_350 ();
 sg13g2_decap_4 FILLER_146_357 ();
 sg13g2_fill_2 FILLER_146_361 ();
 sg13g2_decap_8 FILLER_146_371 ();
 sg13g2_decap_8 FILLER_146_378 ();
 sg13g2_decap_8 FILLER_146_385 ();
 sg13g2_decap_8 FILLER_146_392 ();
 sg13g2_decap_8 FILLER_146_399 ();
 sg13g2_decap_8 FILLER_146_406 ();
 sg13g2_decap_8 FILLER_146_431 ();
 sg13g2_decap_4 FILLER_146_438 ();
 sg13g2_decap_8 FILLER_146_455 ();
 sg13g2_decap_8 FILLER_146_462 ();
 sg13g2_decap_8 FILLER_146_469 ();
 sg13g2_decap_8 FILLER_146_476 ();
 sg13g2_decap_8 FILLER_146_483 ();
 sg13g2_decap_8 FILLER_146_490 ();
 sg13g2_decap_8 FILLER_146_497 ();
 sg13g2_decap_4 FILLER_146_504 ();
 sg13g2_fill_2 FILLER_146_508 ();
 sg13g2_fill_1 FILLER_146_515 ();
 sg13g2_decap_8 FILLER_146_519 ();
 sg13g2_decap_8 FILLER_146_526 ();
 sg13g2_decap_8 FILLER_146_533 ();
 sg13g2_decap_8 FILLER_146_540 ();
 sg13g2_decap_8 FILLER_146_547 ();
 sg13g2_decap_8 FILLER_146_554 ();
 sg13g2_decap_8 FILLER_146_561 ();
 sg13g2_decap_8 FILLER_146_568 ();
 sg13g2_decap_8 FILLER_146_575 ();
 sg13g2_decap_8 FILLER_146_582 ();
 sg13g2_decap_4 FILLER_146_589 ();
 sg13g2_decap_8 FILLER_146_606 ();
 sg13g2_decap_8 FILLER_146_613 ();
 sg13g2_decap_8 FILLER_146_620 ();
 sg13g2_decap_8 FILLER_146_627 ();
 sg13g2_fill_1 FILLER_146_634 ();
 sg13g2_fill_1 FILLER_146_643 ();
 sg13g2_decap_8 FILLER_146_656 ();
 sg13g2_decap_8 FILLER_146_663 ();
 sg13g2_decap_8 FILLER_146_670 ();
 sg13g2_decap_8 FILLER_146_677 ();
 sg13g2_decap_8 FILLER_146_684 ();
 sg13g2_decap_8 FILLER_146_691 ();
 sg13g2_decap_8 FILLER_146_698 ();
 sg13g2_decap_8 FILLER_146_705 ();
 sg13g2_decap_8 FILLER_146_712 ();
 sg13g2_decap_8 FILLER_146_719 ();
 sg13g2_decap_8 FILLER_146_736 ();
 sg13g2_decap_8 FILLER_146_743 ();
 sg13g2_decap_8 FILLER_146_750 ();
 sg13g2_decap_8 FILLER_146_757 ();
 sg13g2_decap_8 FILLER_146_764 ();
 sg13g2_decap_8 FILLER_146_771 ();
 sg13g2_decap_8 FILLER_146_778 ();
 sg13g2_fill_1 FILLER_146_785 ();
 sg13g2_decap_8 FILLER_146_801 ();
 sg13g2_decap_4 FILLER_146_808 ();
 sg13g2_decap_8 FILLER_146_828 ();
 sg13g2_decap_8 FILLER_146_835 ();
 sg13g2_decap_8 FILLER_146_842 ();
 sg13g2_decap_8 FILLER_146_849 ();
 sg13g2_decap_8 FILLER_146_856 ();
 sg13g2_decap_4 FILLER_146_863 ();
 sg13g2_fill_2 FILLER_146_867 ();
 sg13g2_decap_8 FILLER_146_885 ();
 sg13g2_decap_8 FILLER_146_892 ();
 sg13g2_decap_8 FILLER_146_899 ();
 sg13g2_fill_2 FILLER_146_906 ();
 sg13g2_fill_1 FILLER_146_908 ();
 sg13g2_decap_8 FILLER_146_917 ();
 sg13g2_decap_8 FILLER_146_924 ();
 sg13g2_decap_4 FILLER_146_931 ();
 sg13g2_fill_2 FILLER_146_935 ();
 sg13g2_fill_2 FILLER_146_962 ();
 sg13g2_fill_1 FILLER_146_964 ();
 sg13g2_decap_8 FILLER_146_969 ();
 sg13g2_fill_2 FILLER_146_984 ();
 sg13g2_decap_8 FILLER_146_1005 ();
 sg13g2_decap_8 FILLER_146_1012 ();
 sg13g2_decap_8 FILLER_146_1019 ();
 sg13g2_decap_8 FILLER_146_1026 ();
 sg13g2_decap_4 FILLER_146_1033 ();
 sg13g2_fill_1 FILLER_146_1037 ();
 sg13g2_fill_2 FILLER_146_1047 ();
 sg13g2_fill_1 FILLER_146_1049 ();
 sg13g2_decap_8 FILLER_146_1062 ();
 sg13g2_decap_4 FILLER_146_1069 ();
 sg13g2_fill_2 FILLER_146_1073 ();
 sg13g2_decap_4 FILLER_146_1088 ();
 sg13g2_fill_2 FILLER_146_1092 ();
 sg13g2_decap_4 FILLER_146_1108 ();
 sg13g2_fill_1 FILLER_146_1112 ();
 sg13g2_decap_8 FILLER_146_1117 ();
 sg13g2_decap_8 FILLER_146_1124 ();
 sg13g2_decap_8 FILLER_146_1131 ();
 sg13g2_decap_8 FILLER_146_1138 ();
 sg13g2_decap_8 FILLER_146_1145 ();
 sg13g2_decap_8 FILLER_146_1152 ();
 sg13g2_decap_8 FILLER_146_1159 ();
 sg13g2_decap_8 FILLER_146_1174 ();
 sg13g2_decap_8 FILLER_146_1185 ();
 sg13g2_decap_4 FILLER_146_1192 ();
 sg13g2_fill_1 FILLER_146_1196 ();
 sg13g2_decap_8 FILLER_146_1202 ();
 sg13g2_decap_8 FILLER_146_1209 ();
 sg13g2_decap_8 FILLER_146_1216 ();
 sg13g2_decap_8 FILLER_146_1223 ();
 sg13g2_decap_4 FILLER_146_1230 ();
 sg13g2_decap_8 FILLER_146_1239 ();
 sg13g2_decap_8 FILLER_146_1246 ();
 sg13g2_decap_4 FILLER_146_1253 ();
 sg13g2_decap_8 FILLER_146_1265 ();
 sg13g2_fill_2 FILLER_146_1272 ();
 sg13g2_decap_8 FILLER_146_1282 ();
 sg13g2_decap_8 FILLER_146_1289 ();
 sg13g2_decap_8 FILLER_146_1296 ();
 sg13g2_decap_4 FILLER_146_1303 ();
 sg13g2_fill_1 FILLER_146_1307 ();
 sg13g2_decap_8 FILLER_146_1311 ();
 sg13g2_decap_8 FILLER_146_1318 ();
 sg13g2_decap_8 FILLER_146_1325 ();
 sg13g2_decap_8 FILLER_146_1332 ();
 sg13g2_decap_8 FILLER_146_1339 ();
 sg13g2_decap_8 FILLER_146_1346 ();
 sg13g2_decap_8 FILLER_146_1353 ();
 sg13g2_decap_8 FILLER_146_1360 ();
 sg13g2_decap_8 FILLER_146_1367 ();
 sg13g2_decap_8 FILLER_146_1374 ();
 sg13g2_decap_8 FILLER_146_1381 ();
 sg13g2_fill_2 FILLER_146_1388 ();
 sg13g2_fill_1 FILLER_146_1390 ();
 sg13g2_decap_4 FILLER_146_1396 ();
 sg13g2_fill_2 FILLER_146_1400 ();
 sg13g2_decap_8 FILLER_146_1409 ();
 sg13g2_decap_8 FILLER_146_1416 ();
 sg13g2_decap_8 FILLER_146_1423 ();
 sg13g2_decap_8 FILLER_146_1430 ();
 sg13g2_decap_8 FILLER_146_1437 ();
 sg13g2_decap_8 FILLER_146_1444 ();
 sg13g2_decap_8 FILLER_146_1451 ();
 sg13g2_decap_8 FILLER_146_1458 ();
 sg13g2_decap_4 FILLER_146_1465 ();
 sg13g2_fill_1 FILLER_146_1469 ();
 sg13g2_decap_8 FILLER_146_1479 ();
 sg13g2_decap_8 FILLER_146_1486 ();
 sg13g2_decap_8 FILLER_146_1493 ();
 sg13g2_decap_8 FILLER_146_1500 ();
 sg13g2_fill_1 FILLER_146_1507 ();
 sg13g2_fill_2 FILLER_146_1517 ();
 sg13g2_fill_1 FILLER_146_1519 ();
 sg13g2_decap_4 FILLER_146_1525 ();
 sg13g2_fill_1 FILLER_146_1529 ();
 sg13g2_decap_8 FILLER_146_1538 ();
 sg13g2_decap_8 FILLER_146_1545 ();
 sg13g2_decap_8 FILLER_146_1552 ();
 sg13g2_decap_8 FILLER_146_1559 ();
 sg13g2_decap_4 FILLER_146_1566 ();
 sg13g2_fill_2 FILLER_146_1570 ();
 sg13g2_fill_2 FILLER_146_1576 ();
 sg13g2_decap_8 FILLER_146_1591 ();
 sg13g2_decap_8 FILLER_146_1598 ();
 sg13g2_decap_8 FILLER_146_1605 ();
 sg13g2_decap_8 FILLER_146_1612 ();
 sg13g2_decap_8 FILLER_146_1619 ();
 sg13g2_decap_8 FILLER_146_1626 ();
 sg13g2_fill_2 FILLER_146_1633 ();
 sg13g2_fill_1 FILLER_146_1635 ();
 sg13g2_decap_8 FILLER_146_1660 ();
 sg13g2_decap_8 FILLER_146_1667 ();
 sg13g2_decap_8 FILLER_146_1674 ();
 sg13g2_decap_8 FILLER_146_1681 ();
 sg13g2_decap_8 FILLER_146_1688 ();
 sg13g2_decap_8 FILLER_146_1695 ();
 sg13g2_decap_8 FILLER_146_1702 ();
 sg13g2_decap_8 FILLER_146_1709 ();
 sg13g2_decap_8 FILLER_146_1716 ();
 sg13g2_decap_8 FILLER_146_1723 ();
 sg13g2_decap_8 FILLER_146_1730 ();
 sg13g2_decap_8 FILLER_146_1737 ();
 sg13g2_decap_8 FILLER_146_1744 ();
 sg13g2_decap_8 FILLER_146_1751 ();
 sg13g2_decap_8 FILLER_146_1758 ();
 sg13g2_fill_2 FILLER_146_1765 ();
 sg13g2_fill_1 FILLER_146_1767 ();
 sg13g2_decap_8 FILLER_147_0 ();
 sg13g2_fill_2 FILLER_147_7 ();
 sg13g2_fill_1 FILLER_147_9 ();
 sg13g2_fill_1 FILLER_147_38 ();
 sg13g2_decap_8 FILLER_147_44 ();
 sg13g2_decap_4 FILLER_147_51 ();
 sg13g2_fill_2 FILLER_147_55 ();
 sg13g2_decap_8 FILLER_147_67 ();
 sg13g2_decap_8 FILLER_147_78 ();
 sg13g2_decap_4 FILLER_147_85 ();
 sg13g2_decap_4 FILLER_147_92 ();
 sg13g2_fill_1 FILLER_147_96 ();
 sg13g2_decap_8 FILLER_147_105 ();
 sg13g2_decap_8 FILLER_147_112 ();
 sg13g2_decap_8 FILLER_147_119 ();
 sg13g2_decap_8 FILLER_147_126 ();
 sg13g2_decap_8 FILLER_147_133 ();
 sg13g2_decap_8 FILLER_147_140 ();
 sg13g2_decap_8 FILLER_147_147 ();
 sg13g2_decap_8 FILLER_147_154 ();
 sg13g2_decap_8 FILLER_147_161 ();
 sg13g2_fill_2 FILLER_147_168 ();
 sg13g2_fill_1 FILLER_147_170 ();
 sg13g2_decap_8 FILLER_147_181 ();
 sg13g2_decap_8 FILLER_147_188 ();
 sg13g2_decap_8 FILLER_147_195 ();
 sg13g2_fill_1 FILLER_147_202 ();
 sg13g2_decap_8 FILLER_147_219 ();
 sg13g2_decap_8 FILLER_147_226 ();
 sg13g2_decap_8 FILLER_147_233 ();
 sg13g2_decap_4 FILLER_147_240 ();
 sg13g2_decap_8 FILLER_147_249 ();
 sg13g2_decap_8 FILLER_147_256 ();
 sg13g2_decap_8 FILLER_147_263 ();
 sg13g2_decap_8 FILLER_147_270 ();
 sg13g2_decap_8 FILLER_147_277 ();
 sg13g2_decap_8 FILLER_147_284 ();
 sg13g2_decap_8 FILLER_147_291 ();
 sg13g2_decap_8 FILLER_147_298 ();
 sg13g2_fill_1 FILLER_147_322 ();
 sg13g2_fill_2 FILLER_147_327 ();
 sg13g2_decap_8 FILLER_147_337 ();
 sg13g2_decap_8 FILLER_147_348 ();
 sg13g2_decap_8 FILLER_147_355 ();
 sg13g2_decap_8 FILLER_147_362 ();
 sg13g2_decap_8 FILLER_147_369 ();
 sg13g2_fill_1 FILLER_147_376 ();
 sg13g2_decap_4 FILLER_147_386 ();
 sg13g2_fill_2 FILLER_147_390 ();
 sg13g2_fill_2 FILLER_147_400 ();
 sg13g2_decap_8 FILLER_147_406 ();
 sg13g2_decap_8 FILLER_147_413 ();
 sg13g2_fill_2 FILLER_147_420 ();
 sg13g2_fill_1 FILLER_147_422 ();
 sg13g2_decap_8 FILLER_147_431 ();
 sg13g2_decap_8 FILLER_147_438 ();
 sg13g2_fill_2 FILLER_147_445 ();
 sg13g2_fill_1 FILLER_147_447 ();
 sg13g2_decap_8 FILLER_147_453 ();
 sg13g2_decap_8 FILLER_147_460 ();
 sg13g2_fill_1 FILLER_147_467 ();
 sg13g2_decap_8 FILLER_147_473 ();
 sg13g2_decap_8 FILLER_147_480 ();
 sg13g2_decap_8 FILLER_147_487 ();
 sg13g2_decap_8 FILLER_147_494 ();
 sg13g2_decap_8 FILLER_147_501 ();
 sg13g2_fill_1 FILLER_147_508 ();
 sg13g2_decap_8 FILLER_147_526 ();
 sg13g2_decap_8 FILLER_147_533 ();
 sg13g2_decap_8 FILLER_147_540 ();
 sg13g2_decap_8 FILLER_147_547 ();
 sg13g2_decap_8 FILLER_147_554 ();
 sg13g2_decap_8 FILLER_147_561 ();
 sg13g2_fill_2 FILLER_147_568 ();
 sg13g2_fill_2 FILLER_147_582 ();
 sg13g2_fill_1 FILLER_147_584 ();
 sg13g2_decap_8 FILLER_147_601 ();
 sg13g2_decap_8 FILLER_147_608 ();
 sg13g2_decap_8 FILLER_147_615 ();
 sg13g2_decap_8 FILLER_147_622 ();
 sg13g2_decap_8 FILLER_147_629 ();
 sg13g2_fill_1 FILLER_147_636 ();
 sg13g2_fill_1 FILLER_147_651 ();
 sg13g2_decap_8 FILLER_147_660 ();
 sg13g2_decap_8 FILLER_147_667 ();
 sg13g2_decap_4 FILLER_147_674 ();
 sg13g2_fill_1 FILLER_147_678 ();
 sg13g2_decap_8 FILLER_147_692 ();
 sg13g2_decap_8 FILLER_147_699 ();
 sg13g2_decap_8 FILLER_147_706 ();
 sg13g2_decap_8 FILLER_147_713 ();
 sg13g2_decap_8 FILLER_147_745 ();
 sg13g2_decap_8 FILLER_147_752 ();
 sg13g2_decap_8 FILLER_147_759 ();
 sg13g2_decap_8 FILLER_147_766 ();
 sg13g2_decap_8 FILLER_147_773 ();
 sg13g2_decap_8 FILLER_147_785 ();
 sg13g2_fill_2 FILLER_147_792 ();
 sg13g2_fill_1 FILLER_147_794 ();
 sg13g2_decap_8 FILLER_147_802 ();
 sg13g2_decap_4 FILLER_147_809 ();
 sg13g2_fill_1 FILLER_147_813 ();
 sg13g2_decap_8 FILLER_147_830 ();
 sg13g2_decap_8 FILLER_147_837 ();
 sg13g2_decap_8 FILLER_147_844 ();
 sg13g2_decap_8 FILLER_147_851 ();
 sg13g2_decap_8 FILLER_147_858 ();
 sg13g2_decap_8 FILLER_147_865 ();
 sg13g2_fill_2 FILLER_147_872 ();
 sg13g2_fill_1 FILLER_147_874 ();
 sg13g2_decap_8 FILLER_147_898 ();
 sg13g2_decap_8 FILLER_147_905 ();
 sg13g2_decap_8 FILLER_147_912 ();
 sg13g2_decap_8 FILLER_147_926 ();
 sg13g2_fill_2 FILLER_147_933 ();
 sg13g2_fill_1 FILLER_147_935 ();
 sg13g2_fill_1 FILLER_147_944 ();
 sg13g2_decap_8 FILLER_147_969 ();
 sg13g2_decap_8 FILLER_147_976 ();
 sg13g2_decap_4 FILLER_147_983 ();
 sg13g2_fill_1 FILLER_147_987 ();
 sg13g2_decap_4 FILLER_147_1004 ();
 sg13g2_decap_8 FILLER_147_1013 ();
 sg13g2_decap_8 FILLER_147_1020 ();
 sg13g2_decap_8 FILLER_147_1027 ();
 sg13g2_decap_4 FILLER_147_1034 ();
 sg13g2_fill_1 FILLER_147_1038 ();
 sg13g2_decap_8 FILLER_147_1043 ();
 sg13g2_decap_8 FILLER_147_1050 ();
 sg13g2_decap_8 FILLER_147_1057 ();
 sg13g2_decap_8 FILLER_147_1064 ();
 sg13g2_decap_8 FILLER_147_1071 ();
 sg13g2_decap_8 FILLER_147_1078 ();
 sg13g2_decap_8 FILLER_147_1093 ();
 sg13g2_decap_8 FILLER_147_1100 ();
 sg13g2_decap_8 FILLER_147_1107 ();
 sg13g2_decap_8 FILLER_147_1114 ();
 sg13g2_fill_2 FILLER_147_1121 ();
 sg13g2_decap_8 FILLER_147_1131 ();
 sg13g2_decap_8 FILLER_147_1138 ();
 sg13g2_decap_8 FILLER_147_1145 ();
 sg13g2_decap_8 FILLER_147_1152 ();
 sg13g2_decap_8 FILLER_147_1159 ();
 sg13g2_decap_4 FILLER_147_1166 ();
 sg13g2_fill_1 FILLER_147_1170 ();
 sg13g2_decap_8 FILLER_147_1176 ();
 sg13g2_decap_8 FILLER_147_1183 ();
 sg13g2_fill_1 FILLER_147_1190 ();
 sg13g2_decap_4 FILLER_147_1206 ();
 sg13g2_decap_8 FILLER_147_1216 ();
 sg13g2_decap_4 FILLER_147_1223 ();
 sg13g2_fill_2 FILLER_147_1227 ();
 sg13g2_decap_8 FILLER_147_1245 ();
 sg13g2_decap_8 FILLER_147_1252 ();
 sg13g2_decap_8 FILLER_147_1259 ();
 sg13g2_decap_8 FILLER_147_1266 ();
 sg13g2_fill_2 FILLER_147_1273 ();
 sg13g2_decap_8 FILLER_147_1283 ();
 sg13g2_decap_8 FILLER_147_1290 ();
 sg13g2_decap_8 FILLER_147_1297 ();
 sg13g2_fill_2 FILLER_147_1304 ();
 sg13g2_decap_8 FILLER_147_1319 ();
 sg13g2_decap_8 FILLER_147_1326 ();
 sg13g2_fill_2 FILLER_147_1333 ();
 sg13g2_decap_8 FILLER_147_1340 ();
 sg13g2_decap_4 FILLER_147_1347 ();
 sg13g2_fill_2 FILLER_147_1351 ();
 sg13g2_decap_8 FILLER_147_1361 ();
 sg13g2_decap_8 FILLER_147_1368 ();
 sg13g2_decap_8 FILLER_147_1375 ();
 sg13g2_decap_8 FILLER_147_1382 ();
 sg13g2_fill_2 FILLER_147_1389 ();
 sg13g2_fill_1 FILLER_147_1391 ();
 sg13g2_decap_8 FILLER_147_1395 ();
 sg13g2_decap_8 FILLER_147_1402 ();
 sg13g2_decap_8 FILLER_147_1409 ();
 sg13g2_decap_8 FILLER_147_1416 ();
 sg13g2_fill_2 FILLER_147_1423 ();
 sg13g2_fill_1 FILLER_147_1425 ();
 sg13g2_fill_1 FILLER_147_1430 ();
 sg13g2_decap_8 FILLER_147_1436 ();
 sg13g2_decap_8 FILLER_147_1443 ();
 sg13g2_decap_8 FILLER_147_1450 ();
 sg13g2_decap_8 FILLER_147_1457 ();
 sg13g2_decap_4 FILLER_147_1464 ();
 sg13g2_fill_1 FILLER_147_1468 ();
 sg13g2_decap_8 FILLER_147_1487 ();
 sg13g2_decap_8 FILLER_147_1494 ();
 sg13g2_decap_8 FILLER_147_1501 ();
 sg13g2_decap_8 FILLER_147_1508 ();
 sg13g2_fill_2 FILLER_147_1515 ();
 sg13g2_fill_1 FILLER_147_1529 ();
 sg13g2_decap_8 FILLER_147_1538 ();
 sg13g2_decap_8 FILLER_147_1545 ();
 sg13g2_decap_8 FILLER_147_1552 ();
 sg13g2_decap_8 FILLER_147_1559 ();
 sg13g2_decap_4 FILLER_147_1566 ();
 sg13g2_fill_1 FILLER_147_1570 ();
 sg13g2_decap_4 FILLER_147_1575 ();
 sg13g2_fill_1 FILLER_147_1579 ();
 sg13g2_decap_8 FILLER_147_1592 ();
 sg13g2_decap_8 FILLER_147_1599 ();
 sg13g2_decap_8 FILLER_147_1606 ();
 sg13g2_decap_8 FILLER_147_1613 ();
 sg13g2_decap_8 FILLER_147_1620 ();
 sg13g2_decap_8 FILLER_147_1627 ();
 sg13g2_fill_1 FILLER_147_1634 ();
 sg13g2_decap_8 FILLER_147_1651 ();
 sg13g2_decap_8 FILLER_147_1658 ();
 sg13g2_decap_8 FILLER_147_1665 ();
 sg13g2_decap_8 FILLER_147_1672 ();
 sg13g2_decap_8 FILLER_147_1679 ();
 sg13g2_decap_8 FILLER_147_1686 ();
 sg13g2_decap_8 FILLER_147_1693 ();
 sg13g2_decap_8 FILLER_147_1700 ();
 sg13g2_decap_8 FILLER_147_1707 ();
 sg13g2_decap_8 FILLER_147_1714 ();
 sg13g2_decap_8 FILLER_147_1721 ();
 sg13g2_decap_8 FILLER_147_1728 ();
 sg13g2_decap_8 FILLER_147_1735 ();
 sg13g2_decap_8 FILLER_147_1742 ();
 sg13g2_decap_8 FILLER_147_1749 ();
 sg13g2_decap_8 FILLER_147_1756 ();
 sg13g2_decap_4 FILLER_147_1763 ();
 sg13g2_fill_1 FILLER_147_1767 ();
 sg13g2_decap_8 FILLER_148_0 ();
 sg13g2_decap_8 FILLER_148_7 ();
 sg13g2_decap_8 FILLER_148_14 ();
 sg13g2_decap_8 FILLER_148_21 ();
 sg13g2_decap_8 FILLER_148_28 ();
 sg13g2_decap_8 FILLER_148_35 ();
 sg13g2_decap_8 FILLER_148_42 ();
 sg13g2_decap_8 FILLER_148_49 ();
 sg13g2_decap_8 FILLER_148_56 ();
 sg13g2_decap_4 FILLER_148_63 ();
 sg13g2_decap_8 FILLER_148_75 ();
 sg13g2_decap_4 FILLER_148_82 ();
 sg13g2_fill_1 FILLER_148_86 ();
 sg13g2_decap_8 FILLER_148_96 ();
 sg13g2_decap_8 FILLER_148_103 ();
 sg13g2_decap_8 FILLER_148_110 ();
 sg13g2_decap_8 FILLER_148_117 ();
 sg13g2_decap_8 FILLER_148_124 ();
 sg13g2_decap_8 FILLER_148_131 ();
 sg13g2_decap_8 FILLER_148_138 ();
 sg13g2_decap_8 FILLER_148_145 ();
 sg13g2_decap_8 FILLER_148_152 ();
 sg13g2_fill_2 FILLER_148_159 ();
 sg13g2_fill_1 FILLER_148_161 ();
 sg13g2_fill_1 FILLER_148_166 ();
 sg13g2_decap_8 FILLER_148_172 ();
 sg13g2_decap_4 FILLER_148_179 ();
 sg13g2_fill_1 FILLER_148_183 ();
 sg13g2_fill_2 FILLER_148_189 ();
 sg13g2_decap_4 FILLER_148_196 ();
 sg13g2_fill_2 FILLER_148_200 ();
 sg13g2_decap_8 FILLER_148_222 ();
 sg13g2_decap_8 FILLER_148_229 ();
 sg13g2_fill_2 FILLER_148_236 ();
 sg13g2_fill_2 FILLER_148_269 ();
 sg13g2_fill_1 FILLER_148_271 ();
 sg13g2_decap_8 FILLER_148_285 ();
 sg13g2_decap_8 FILLER_148_292 ();
 sg13g2_fill_2 FILLER_148_299 ();
 sg13g2_fill_1 FILLER_148_301 ();
 sg13g2_fill_1 FILLER_148_332 ();
 sg13g2_decap_8 FILLER_148_359 ();
 sg13g2_decap_8 FILLER_148_366 ();
 sg13g2_decap_8 FILLER_148_373 ();
 sg13g2_decap_4 FILLER_148_380 ();
 sg13g2_fill_2 FILLER_148_384 ();
 sg13g2_decap_8 FILLER_148_391 ();
 sg13g2_decap_8 FILLER_148_398 ();
 sg13g2_decap_8 FILLER_148_405 ();
 sg13g2_decap_8 FILLER_148_412 ();
 sg13g2_decap_8 FILLER_148_419 ();
 sg13g2_decap_8 FILLER_148_426 ();
 sg13g2_decap_8 FILLER_148_433 ();
 sg13g2_decap_8 FILLER_148_440 ();
 sg13g2_decap_8 FILLER_148_447 ();
 sg13g2_decap_8 FILLER_148_454 ();
 sg13g2_decap_4 FILLER_148_461 ();
 sg13g2_decap_8 FILLER_148_485 ();
 sg13g2_decap_4 FILLER_148_492 ();
 sg13g2_fill_1 FILLER_148_528 ();
 sg13g2_decap_8 FILLER_148_545 ();
 sg13g2_decap_8 FILLER_148_552 ();
 sg13g2_decap_8 FILLER_148_559 ();
 sg13g2_decap_8 FILLER_148_566 ();
 sg13g2_decap_8 FILLER_148_573 ();
 sg13g2_fill_2 FILLER_148_593 ();
 sg13g2_decap_8 FILLER_148_603 ();
 sg13g2_decap_4 FILLER_148_610 ();
 sg13g2_decap_8 FILLER_148_622 ();
 sg13g2_decap_8 FILLER_148_629 ();
 sg13g2_decap_8 FILLER_148_636 ();
 sg13g2_decap_8 FILLER_148_643 ();
 sg13g2_fill_2 FILLER_148_650 ();
 sg13g2_fill_1 FILLER_148_652 ();
 sg13g2_decap_8 FILLER_148_665 ();
 sg13g2_decap_8 FILLER_148_672 ();
 sg13g2_decap_4 FILLER_148_679 ();
 sg13g2_fill_1 FILLER_148_683 ();
 sg13g2_fill_2 FILLER_148_689 ();
 sg13g2_fill_1 FILLER_148_691 ();
 sg13g2_decap_8 FILLER_148_704 ();
 sg13g2_decap_8 FILLER_148_711 ();
 sg13g2_decap_8 FILLER_148_718 ();
 sg13g2_decap_8 FILLER_148_725 ();
 sg13g2_decap_8 FILLER_148_732 ();
 sg13g2_fill_2 FILLER_148_739 ();
 sg13g2_fill_1 FILLER_148_741 ();
 sg13g2_decap_8 FILLER_148_762 ();
 sg13g2_decap_4 FILLER_148_769 ();
 sg13g2_fill_2 FILLER_148_773 ();
 sg13g2_decap_8 FILLER_148_787 ();
 sg13g2_decap_8 FILLER_148_794 ();
 sg13g2_decap_8 FILLER_148_801 ();
 sg13g2_decap_8 FILLER_148_808 ();
 sg13g2_decap_8 FILLER_148_815 ();
 sg13g2_decap_8 FILLER_148_822 ();
 sg13g2_decap_8 FILLER_148_829 ();
 sg13g2_decap_8 FILLER_148_836 ();
 sg13g2_decap_8 FILLER_148_843 ();
 sg13g2_decap_4 FILLER_148_850 ();
 sg13g2_fill_2 FILLER_148_854 ();
 sg13g2_decap_8 FILLER_148_860 ();
 sg13g2_decap_8 FILLER_148_867 ();
 sg13g2_decap_4 FILLER_148_874 ();
 sg13g2_fill_2 FILLER_148_878 ();
 sg13g2_decap_8 FILLER_148_886 ();
 sg13g2_decap_8 FILLER_148_893 ();
 sg13g2_decap_4 FILLER_148_900 ();
 sg13g2_fill_1 FILLER_148_904 ();
 sg13g2_decap_8 FILLER_148_912 ();
 sg13g2_decap_8 FILLER_148_919 ();
 sg13g2_decap_8 FILLER_148_926 ();
 sg13g2_decap_8 FILLER_148_933 ();
 sg13g2_decap_8 FILLER_148_940 ();
 sg13g2_decap_8 FILLER_148_947 ();
 sg13g2_decap_8 FILLER_148_954 ();
 sg13g2_decap_8 FILLER_148_961 ();
 sg13g2_decap_8 FILLER_148_968 ();
 sg13g2_decap_8 FILLER_148_975 ();
 sg13g2_decap_8 FILLER_148_982 ();
 sg13g2_decap_8 FILLER_148_989 ();
 sg13g2_decap_8 FILLER_148_996 ();
 sg13g2_fill_2 FILLER_148_1019 ();
 sg13g2_fill_1 FILLER_148_1021 ();
 sg13g2_decap_8 FILLER_148_1049 ();
 sg13g2_decap_8 FILLER_148_1060 ();
 sg13g2_fill_1 FILLER_148_1067 ();
 sg13g2_decap_8 FILLER_148_1073 ();
 sg13g2_decap_4 FILLER_148_1080 ();
 sg13g2_fill_1 FILLER_148_1084 ();
 sg13g2_decap_8 FILLER_148_1089 ();
 sg13g2_decap_8 FILLER_148_1096 ();
 sg13g2_decap_8 FILLER_148_1103 ();
 sg13g2_decap_4 FILLER_148_1110 ();
 sg13g2_fill_2 FILLER_148_1114 ();
 sg13g2_decap_8 FILLER_148_1137 ();
 sg13g2_decap_8 FILLER_148_1144 ();
 sg13g2_decap_8 FILLER_148_1151 ();
 sg13g2_decap_8 FILLER_148_1158 ();
 sg13g2_fill_2 FILLER_148_1165 ();
 sg13g2_decap_4 FILLER_148_1186 ();
 sg13g2_decap_8 FILLER_148_1199 ();
 sg13g2_decap_4 FILLER_148_1206 ();
 sg13g2_decap_8 FILLER_148_1218 ();
 sg13g2_decap_8 FILLER_148_1225 ();
 sg13g2_fill_2 FILLER_148_1232 ();
 sg13g2_fill_1 FILLER_148_1234 ();
 sg13g2_decap_4 FILLER_148_1251 ();
 sg13g2_fill_2 FILLER_148_1268 ();
 sg13g2_decap_8 FILLER_148_1278 ();
 sg13g2_decap_8 FILLER_148_1285 ();
 sg13g2_decap_8 FILLER_148_1292 ();
 sg13g2_fill_1 FILLER_148_1299 ();
 sg13g2_decap_8 FILLER_148_1324 ();
 sg13g2_decap_8 FILLER_148_1349 ();
 sg13g2_decap_4 FILLER_148_1356 ();
 sg13g2_fill_1 FILLER_148_1360 ();
 sg13g2_decap_4 FILLER_148_1365 ();
 sg13g2_decap_8 FILLER_148_1381 ();
 sg13g2_decap_4 FILLER_148_1388 ();
 sg13g2_decap_8 FILLER_148_1409 ();
 sg13g2_decap_4 FILLER_148_1416 ();
 sg13g2_decap_8 FILLER_148_1437 ();
 sg13g2_decap_8 FILLER_148_1444 ();
 sg13g2_decap_4 FILLER_148_1451 ();
 sg13g2_decap_8 FILLER_148_1480 ();
 sg13g2_decap_8 FILLER_148_1503 ();
 sg13g2_decap_8 FILLER_148_1510 ();
 sg13g2_decap_4 FILLER_148_1517 ();
 sg13g2_decap_8 FILLER_148_1525 ();
 sg13g2_decap_8 FILLER_148_1532 ();
 sg13g2_decap_8 FILLER_148_1539 ();
 sg13g2_fill_2 FILLER_148_1546 ();
 sg13g2_fill_1 FILLER_148_1548 ();
 sg13g2_decap_8 FILLER_148_1558 ();
 sg13g2_fill_2 FILLER_148_1565 ();
 sg13g2_decap_8 FILLER_148_1594 ();
 sg13g2_decap_8 FILLER_148_1601 ();
 sg13g2_decap_8 FILLER_148_1608 ();
 sg13g2_decap_8 FILLER_148_1615 ();
 sg13g2_decap_8 FILLER_148_1622 ();
 sg13g2_decap_8 FILLER_148_1629 ();
 sg13g2_decap_8 FILLER_148_1636 ();
 sg13g2_decap_8 FILLER_148_1643 ();
 sg13g2_decap_8 FILLER_148_1650 ();
 sg13g2_decap_8 FILLER_148_1657 ();
 sg13g2_decap_8 FILLER_148_1664 ();
 sg13g2_decap_8 FILLER_148_1671 ();
 sg13g2_decap_8 FILLER_148_1678 ();
 sg13g2_decap_8 FILLER_148_1685 ();
 sg13g2_decap_8 FILLER_148_1692 ();
 sg13g2_decap_8 FILLER_148_1699 ();
 sg13g2_decap_8 FILLER_148_1706 ();
 sg13g2_decap_8 FILLER_148_1713 ();
 sg13g2_decap_8 FILLER_148_1720 ();
 sg13g2_decap_8 FILLER_148_1727 ();
 sg13g2_decap_8 FILLER_148_1734 ();
 sg13g2_decap_8 FILLER_148_1741 ();
 sg13g2_decap_8 FILLER_148_1748 ();
 sg13g2_decap_8 FILLER_148_1755 ();
 sg13g2_decap_4 FILLER_148_1762 ();
 sg13g2_fill_2 FILLER_148_1766 ();
 sg13g2_decap_8 FILLER_149_0 ();
 sg13g2_decap_8 FILLER_149_7 ();
 sg13g2_decap_8 FILLER_149_14 ();
 sg13g2_decap_8 FILLER_149_21 ();
 sg13g2_decap_8 FILLER_149_28 ();
 sg13g2_decap_8 FILLER_149_39 ();
 sg13g2_decap_4 FILLER_149_46 ();
 sg13g2_fill_1 FILLER_149_66 ();
 sg13g2_decap_8 FILLER_149_71 ();
 sg13g2_decap_8 FILLER_149_78 ();
 sg13g2_fill_2 FILLER_149_85 ();
 sg13g2_fill_1 FILLER_149_87 ();
 sg13g2_decap_8 FILLER_149_97 ();
 sg13g2_decap_8 FILLER_149_104 ();
 sg13g2_decap_8 FILLER_149_111 ();
 sg13g2_decap_8 FILLER_149_118 ();
 sg13g2_decap_8 FILLER_149_125 ();
 sg13g2_decap_8 FILLER_149_132 ();
 sg13g2_decap_8 FILLER_149_139 ();
 sg13g2_decap_8 FILLER_149_146 ();
 sg13g2_decap_4 FILLER_149_153 ();
 sg13g2_fill_2 FILLER_149_157 ();
 sg13g2_decap_8 FILLER_149_168 ();
 sg13g2_fill_2 FILLER_149_175 ();
 sg13g2_decap_8 FILLER_149_196 ();
 sg13g2_decap_8 FILLER_149_203 ();
 sg13g2_fill_1 FILLER_149_210 ();
 sg13g2_decap_8 FILLER_149_216 ();
 sg13g2_decap_8 FILLER_149_223 ();
 sg13g2_decap_8 FILLER_149_243 ();
 sg13g2_decap_4 FILLER_149_250 ();
 sg13g2_decap_8 FILLER_149_258 ();
 sg13g2_decap_8 FILLER_149_265 ();
 sg13g2_decap_8 FILLER_149_272 ();
 sg13g2_decap_8 FILLER_149_279 ();
 sg13g2_decap_4 FILLER_149_286 ();
 sg13g2_fill_1 FILLER_149_290 ();
 sg13g2_decap_8 FILLER_149_325 ();
 sg13g2_fill_1 FILLER_149_332 ();
 sg13g2_decap_8 FILLER_149_344 ();
 sg13g2_decap_8 FILLER_149_351 ();
 sg13g2_decap_8 FILLER_149_358 ();
 sg13g2_decap_8 FILLER_149_365 ();
 sg13g2_fill_1 FILLER_149_372 ();
 sg13g2_fill_1 FILLER_149_393 ();
 sg13g2_fill_1 FILLER_149_402 ();
 sg13g2_decap_8 FILLER_149_408 ();
 sg13g2_decap_8 FILLER_149_415 ();
 sg13g2_decap_8 FILLER_149_422 ();
 sg13g2_decap_8 FILLER_149_429 ();
 sg13g2_decap_8 FILLER_149_436 ();
 sg13g2_decap_8 FILLER_149_443 ();
 sg13g2_decap_8 FILLER_149_450 ();
 sg13g2_decap_4 FILLER_149_467 ();
 sg13g2_decap_8 FILLER_149_481 ();
 sg13g2_decap_8 FILLER_149_488 ();
 sg13g2_fill_2 FILLER_149_495 ();
 sg13g2_decap_4 FILLER_149_505 ();
 sg13g2_fill_2 FILLER_149_509 ();
 sg13g2_fill_2 FILLER_149_516 ();
 sg13g2_decap_8 FILLER_149_526 ();
 sg13g2_fill_2 FILLER_149_533 ();
 sg13g2_decap_8 FILLER_149_551 ();
 sg13g2_decap_8 FILLER_149_558 ();
 sg13g2_decap_8 FILLER_149_565 ();
 sg13g2_decap_8 FILLER_149_572 ();
 sg13g2_fill_2 FILLER_149_587 ();
 sg13g2_decap_8 FILLER_149_599 ();
 sg13g2_decap_8 FILLER_149_606 ();
 sg13g2_decap_8 FILLER_149_613 ();
 sg13g2_decap_8 FILLER_149_620 ();
 sg13g2_decap_8 FILLER_149_627 ();
 sg13g2_decap_8 FILLER_149_634 ();
 sg13g2_decap_8 FILLER_149_641 ();
 sg13g2_decap_8 FILLER_149_648 ();
 sg13g2_decap_8 FILLER_149_655 ();
 sg13g2_decap_8 FILLER_149_662 ();
 sg13g2_fill_2 FILLER_149_669 ();
 sg13g2_fill_1 FILLER_149_671 ();
 sg13g2_fill_2 FILLER_149_682 ();
 sg13g2_fill_1 FILLER_149_684 ();
 sg13g2_decap_8 FILLER_149_695 ();
 sg13g2_decap_4 FILLER_149_702 ();
 sg13g2_decap_8 FILLER_149_718 ();
 sg13g2_decap_8 FILLER_149_725 ();
 sg13g2_decap_8 FILLER_149_732 ();
 sg13g2_decap_8 FILLER_149_739 ();
 sg13g2_fill_2 FILLER_149_746 ();
 sg13g2_fill_1 FILLER_149_748 ();
 sg13g2_decap_8 FILLER_149_757 ();
 sg13g2_decap_8 FILLER_149_764 ();
 sg13g2_decap_8 FILLER_149_771 ();
 sg13g2_decap_8 FILLER_149_778 ();
 sg13g2_decap_4 FILLER_149_785 ();
 sg13g2_fill_1 FILLER_149_793 ();
 sg13g2_fill_1 FILLER_149_802 ();
 sg13g2_decap_8 FILLER_149_820 ();
 sg13g2_decap_8 FILLER_149_827 ();
 sg13g2_decap_8 FILLER_149_834 ();
 sg13g2_decap_8 FILLER_149_841 ();
 sg13g2_decap_4 FILLER_149_848 ();
 sg13g2_decap_8 FILLER_149_880 ();
 sg13g2_decap_8 FILLER_149_887 ();
 sg13g2_decap_4 FILLER_149_894 ();
 sg13g2_fill_1 FILLER_149_898 ();
 sg13g2_decap_8 FILLER_149_914 ();
 sg13g2_decap_8 FILLER_149_921 ();
 sg13g2_decap_8 FILLER_149_928 ();
 sg13g2_decap_8 FILLER_149_935 ();
 sg13g2_fill_2 FILLER_149_942 ();
 sg13g2_fill_1 FILLER_149_944 ();
 sg13g2_decap_8 FILLER_149_949 ();
 sg13g2_decap_8 FILLER_149_956 ();
 sg13g2_decap_4 FILLER_149_963 ();
 sg13g2_decap_8 FILLER_149_975 ();
 sg13g2_decap_8 FILLER_149_982 ();
 sg13g2_decap_8 FILLER_149_989 ();
 sg13g2_decap_8 FILLER_149_996 ();
 sg13g2_decap_4 FILLER_149_1003 ();
 sg13g2_decap_4 FILLER_149_1011 ();
 sg13g2_fill_1 FILLER_149_1015 ();
 sg13g2_fill_2 FILLER_149_1024 ();
 sg13g2_decap_8 FILLER_149_1044 ();
 sg13g2_decap_4 FILLER_149_1051 ();
 sg13g2_decap_8 FILLER_149_1060 ();
 sg13g2_decap_4 FILLER_149_1067 ();
 sg13g2_fill_1 FILLER_149_1071 ();
 sg13g2_decap_4 FILLER_149_1080 ();
 sg13g2_decap_8 FILLER_149_1096 ();
 sg13g2_decap_8 FILLER_149_1103 ();
 sg13g2_decap_8 FILLER_149_1110 ();
 sg13g2_decap_8 FILLER_149_1117 ();
 sg13g2_decap_4 FILLER_149_1124 ();
 sg13g2_fill_1 FILLER_149_1128 ();
 sg13g2_decap_8 FILLER_149_1137 ();
 sg13g2_decap_8 FILLER_149_1144 ();
 sg13g2_decap_8 FILLER_149_1151 ();
 sg13g2_decap_8 FILLER_149_1158 ();
 sg13g2_decap_4 FILLER_149_1165 ();
 sg13g2_fill_2 FILLER_149_1169 ();
 sg13g2_fill_2 FILLER_149_1175 ();
 sg13g2_fill_1 FILLER_149_1177 ();
 sg13g2_decap_8 FILLER_149_1192 ();
 sg13g2_decap_8 FILLER_149_1199 ();
 sg13g2_decap_8 FILLER_149_1206 ();
 sg13g2_fill_1 FILLER_149_1213 ();
 sg13g2_decap_8 FILLER_149_1222 ();
 sg13g2_decap_8 FILLER_149_1229 ();
 sg13g2_decap_8 FILLER_149_1236 ();
 sg13g2_fill_2 FILLER_149_1243 ();
 sg13g2_decap_8 FILLER_149_1250 ();
 sg13g2_fill_2 FILLER_149_1257 ();
 sg13g2_decap_8 FILLER_149_1271 ();
 sg13g2_decap_8 FILLER_149_1278 ();
 sg13g2_decap_4 FILLER_149_1285 ();
 sg13g2_decap_8 FILLER_149_1295 ();
 sg13g2_decap_4 FILLER_149_1302 ();
 sg13g2_fill_1 FILLER_149_1306 ();
 sg13g2_decap_8 FILLER_149_1320 ();
 sg13g2_decap_8 FILLER_149_1327 ();
 sg13g2_decap_8 FILLER_149_1334 ();
 sg13g2_fill_2 FILLER_149_1341 ();
 sg13g2_fill_1 FILLER_149_1343 ();
 sg13g2_decap_8 FILLER_149_1349 ();
 sg13g2_fill_1 FILLER_149_1356 ();
 sg13g2_fill_2 FILLER_149_1381 ();
 sg13g2_decap_8 FILLER_149_1388 ();
 sg13g2_decap_8 FILLER_149_1395 ();
 sg13g2_decap_8 FILLER_149_1402 ();
 sg13g2_decap_8 FILLER_149_1409 ();
 sg13g2_decap_8 FILLER_149_1416 ();
 sg13g2_decap_4 FILLER_149_1423 ();
 sg13g2_fill_1 FILLER_149_1427 ();
 sg13g2_decap_8 FILLER_149_1451 ();
 sg13g2_decap_8 FILLER_149_1458 ();
 sg13g2_decap_8 FILLER_149_1465 ();
 sg13g2_fill_1 FILLER_149_1472 ();
 sg13g2_decap_4 FILLER_149_1482 ();
 sg13g2_fill_2 FILLER_149_1486 ();
 sg13g2_decap_4 FILLER_149_1491 ();
 sg13g2_fill_2 FILLER_149_1495 ();
 sg13g2_fill_2 FILLER_149_1510 ();
 sg13g2_fill_2 FILLER_149_1517 ();
 sg13g2_fill_1 FILLER_149_1524 ();
 sg13g2_decap_8 FILLER_149_1529 ();
 sg13g2_decap_8 FILLER_149_1536 ();
 sg13g2_decap_8 FILLER_149_1543 ();
 sg13g2_decap_8 FILLER_149_1550 ();
 sg13g2_decap_8 FILLER_149_1557 ();
 sg13g2_decap_8 FILLER_149_1564 ();
 sg13g2_decap_4 FILLER_149_1571 ();
 sg13g2_fill_1 FILLER_149_1575 ();
 sg13g2_decap_8 FILLER_149_1589 ();
 sg13g2_decap_8 FILLER_149_1596 ();
 sg13g2_decap_8 FILLER_149_1603 ();
 sg13g2_decap_8 FILLER_149_1610 ();
 sg13g2_decap_8 FILLER_149_1617 ();
 sg13g2_decap_8 FILLER_149_1624 ();
 sg13g2_decap_8 FILLER_149_1631 ();
 sg13g2_decap_8 FILLER_149_1638 ();
 sg13g2_decap_8 FILLER_149_1645 ();
 sg13g2_decap_8 FILLER_149_1652 ();
 sg13g2_decap_8 FILLER_149_1659 ();
 sg13g2_decap_8 FILLER_149_1666 ();
 sg13g2_decap_8 FILLER_149_1673 ();
 sg13g2_decap_8 FILLER_149_1680 ();
 sg13g2_decap_8 FILLER_149_1687 ();
 sg13g2_decap_8 FILLER_149_1694 ();
 sg13g2_decap_8 FILLER_149_1701 ();
 sg13g2_decap_8 FILLER_149_1708 ();
 sg13g2_decap_8 FILLER_149_1715 ();
 sg13g2_decap_8 FILLER_149_1722 ();
 sg13g2_decap_8 FILLER_149_1729 ();
 sg13g2_decap_8 FILLER_149_1736 ();
 sg13g2_decap_8 FILLER_149_1743 ();
 sg13g2_decap_8 FILLER_149_1750 ();
 sg13g2_decap_8 FILLER_149_1757 ();
 sg13g2_decap_4 FILLER_149_1764 ();
 sg13g2_decap_8 FILLER_150_0 ();
 sg13g2_decap_8 FILLER_150_7 ();
 sg13g2_decap_8 FILLER_150_14 ();
 sg13g2_decap_8 FILLER_150_21 ();
 sg13g2_fill_2 FILLER_150_28 ();
 sg13g2_decap_8 FILLER_150_51 ();
 sg13g2_decap_8 FILLER_150_58 ();
 sg13g2_decap_8 FILLER_150_65 ();
 sg13g2_decap_8 FILLER_150_72 ();
 sg13g2_decap_8 FILLER_150_79 ();
 sg13g2_decap_8 FILLER_150_86 ();
 sg13g2_decap_4 FILLER_150_93 ();
 sg13g2_fill_1 FILLER_150_97 ();
 sg13g2_fill_2 FILLER_150_106 ();
 sg13g2_fill_1 FILLER_150_108 ();
 sg13g2_decap_8 FILLER_150_122 ();
 sg13g2_decap_8 FILLER_150_129 ();
 sg13g2_decap_8 FILLER_150_136 ();
 sg13g2_decap_4 FILLER_150_143 ();
 sg13g2_fill_1 FILLER_150_147 ();
 sg13g2_fill_2 FILLER_150_152 ();
 sg13g2_decap_8 FILLER_150_161 ();
 sg13g2_decap_8 FILLER_150_168 ();
 sg13g2_decap_8 FILLER_150_175 ();
 sg13g2_decap_8 FILLER_150_182 ();
 sg13g2_decap_8 FILLER_150_189 ();
 sg13g2_decap_8 FILLER_150_196 ();
 sg13g2_decap_8 FILLER_150_203 ();
 sg13g2_decap_8 FILLER_150_210 ();
 sg13g2_decap_8 FILLER_150_217 ();
 sg13g2_fill_1 FILLER_150_224 ();
 sg13g2_decap_8 FILLER_150_231 ();
 sg13g2_decap_8 FILLER_150_238 ();
 sg13g2_decap_8 FILLER_150_245 ();
 sg13g2_decap_8 FILLER_150_252 ();
 sg13g2_decap_8 FILLER_150_259 ();
 sg13g2_decap_8 FILLER_150_266 ();
 sg13g2_decap_8 FILLER_150_273 ();
 sg13g2_decap_8 FILLER_150_280 ();
 sg13g2_decap_8 FILLER_150_287 ();
 sg13g2_decap_8 FILLER_150_294 ();
 sg13g2_fill_1 FILLER_150_301 ();
 sg13g2_decap_8 FILLER_150_315 ();
 sg13g2_decap_8 FILLER_150_322 ();
 sg13g2_decap_8 FILLER_150_329 ();
 sg13g2_decap_8 FILLER_150_340 ();
 sg13g2_decap_8 FILLER_150_347 ();
 sg13g2_decap_8 FILLER_150_354 ();
 sg13g2_decap_8 FILLER_150_361 ();
 sg13g2_decap_8 FILLER_150_368 ();
 sg13g2_fill_2 FILLER_150_375 ();
 sg13g2_decap_8 FILLER_150_394 ();
 sg13g2_decap_4 FILLER_150_401 ();
 sg13g2_fill_2 FILLER_150_405 ();
 sg13g2_decap_8 FILLER_150_415 ();
 sg13g2_fill_2 FILLER_150_422 ();
 sg13g2_decap_4 FILLER_150_428 ();
 sg13g2_fill_1 FILLER_150_432 ();
 sg13g2_decap_8 FILLER_150_437 ();
 sg13g2_decap_4 FILLER_150_444 ();
 sg13g2_fill_2 FILLER_150_448 ();
 sg13g2_decap_8 FILLER_150_454 ();
 sg13g2_decap_8 FILLER_150_461 ();
 sg13g2_decap_8 FILLER_150_468 ();
 sg13g2_decap_8 FILLER_150_475 ();
 sg13g2_decap_8 FILLER_150_482 ();
 sg13g2_decap_8 FILLER_150_489 ();
 sg13g2_decap_8 FILLER_150_496 ();
 sg13g2_decap_8 FILLER_150_503 ();
 sg13g2_decap_8 FILLER_150_510 ();
 sg13g2_decap_8 FILLER_150_517 ();
 sg13g2_decap_8 FILLER_150_524 ();
 sg13g2_decap_8 FILLER_150_531 ();
 sg13g2_decap_8 FILLER_150_538 ();
 sg13g2_decap_8 FILLER_150_545 ();
 sg13g2_decap_8 FILLER_150_552 ();
 sg13g2_decap_8 FILLER_150_559 ();
 sg13g2_decap_4 FILLER_150_566 ();
 sg13g2_decap_8 FILLER_150_594 ();
 sg13g2_decap_8 FILLER_150_601 ();
 sg13g2_decap_8 FILLER_150_608 ();
 sg13g2_decap_8 FILLER_150_615 ();
 sg13g2_fill_2 FILLER_150_622 ();
 sg13g2_decap_8 FILLER_150_637 ();
 sg13g2_decap_8 FILLER_150_644 ();
 sg13g2_decap_8 FILLER_150_651 ();
 sg13g2_decap_8 FILLER_150_658 ();
 sg13g2_decap_8 FILLER_150_665 ();
 sg13g2_fill_2 FILLER_150_672 ();
 sg13g2_decap_8 FILLER_150_677 ();
 sg13g2_decap_8 FILLER_150_684 ();
 sg13g2_fill_2 FILLER_150_691 ();
 sg13g2_decap_4 FILLER_150_701 ();
 sg13g2_decap_8 FILLER_150_721 ();
 sg13g2_fill_2 FILLER_150_728 ();
 sg13g2_fill_1 FILLER_150_730 ();
 sg13g2_decap_8 FILLER_150_749 ();
 sg13g2_decap_8 FILLER_150_756 ();
 sg13g2_decap_8 FILLER_150_763 ();
 sg13g2_decap_8 FILLER_150_770 ();
 sg13g2_decap_8 FILLER_150_777 ();
 sg13g2_decap_8 FILLER_150_804 ();
 sg13g2_decap_8 FILLER_150_811 ();
 sg13g2_decap_8 FILLER_150_818 ();
 sg13g2_decap_4 FILLER_150_825 ();
 sg13g2_fill_2 FILLER_150_829 ();
 sg13g2_decap_8 FILLER_150_835 ();
 sg13g2_decap_4 FILLER_150_842 ();
 sg13g2_fill_1 FILLER_150_862 ();
 sg13g2_decap_8 FILLER_150_879 ();
 sg13g2_decap_8 FILLER_150_886 ();
 sg13g2_fill_2 FILLER_150_893 ();
 sg13g2_fill_1 FILLER_150_895 ();
 sg13g2_decap_8 FILLER_150_909 ();
 sg13g2_decap_8 FILLER_150_916 ();
 sg13g2_decap_8 FILLER_150_923 ();
 sg13g2_decap_4 FILLER_150_930 ();
 sg13g2_decap_8 FILLER_150_955 ();
 sg13g2_decap_8 FILLER_150_962 ();
 sg13g2_decap_8 FILLER_150_969 ();
 sg13g2_decap_8 FILLER_150_976 ();
 sg13g2_decap_8 FILLER_150_983 ();
 sg13g2_decap_8 FILLER_150_990 ();
 sg13g2_decap_8 FILLER_150_997 ();
 sg13g2_decap_8 FILLER_150_1004 ();
 sg13g2_decap_8 FILLER_150_1011 ();
 sg13g2_decap_8 FILLER_150_1018 ();
 sg13g2_decap_8 FILLER_150_1025 ();
 sg13g2_fill_2 FILLER_150_1032 ();
 sg13g2_fill_1 FILLER_150_1034 ();
 sg13g2_decap_8 FILLER_150_1040 ();
 sg13g2_decap_8 FILLER_150_1047 ();
 sg13g2_decap_8 FILLER_150_1054 ();
 sg13g2_decap_8 FILLER_150_1061 ();
 sg13g2_decap_8 FILLER_150_1068 ();
 sg13g2_decap_8 FILLER_150_1075 ();
 sg13g2_fill_1 FILLER_150_1090 ();
 sg13g2_decap_8 FILLER_150_1096 ();
 sg13g2_decap_8 FILLER_150_1103 ();
 sg13g2_decap_8 FILLER_150_1110 ();
 sg13g2_decap_8 FILLER_150_1117 ();
 sg13g2_decap_8 FILLER_150_1124 ();
 sg13g2_decap_8 FILLER_150_1131 ();
 sg13g2_decap_8 FILLER_150_1138 ();
 sg13g2_decap_8 FILLER_150_1145 ();
 sg13g2_decap_8 FILLER_150_1152 ();
 sg13g2_decap_8 FILLER_150_1159 ();
 sg13g2_decap_8 FILLER_150_1166 ();
 sg13g2_decap_8 FILLER_150_1189 ();
 sg13g2_decap_8 FILLER_150_1196 ();
 sg13g2_decap_4 FILLER_150_1203 ();
 sg13g2_fill_1 FILLER_150_1207 ();
 sg13g2_fill_2 FILLER_150_1216 ();
 sg13g2_decap_8 FILLER_150_1226 ();
 sg13g2_decap_8 FILLER_150_1233 ();
 sg13g2_fill_2 FILLER_150_1240 ();
 sg13g2_fill_1 FILLER_150_1242 ();
 sg13g2_decap_8 FILLER_150_1251 ();
 sg13g2_fill_2 FILLER_150_1258 ();
 sg13g2_fill_1 FILLER_150_1260 ();
 sg13g2_decap_4 FILLER_150_1277 ();
 sg13g2_fill_2 FILLER_150_1281 ();
 sg13g2_decap_8 FILLER_150_1291 ();
 sg13g2_decap_8 FILLER_150_1298 ();
 sg13g2_fill_1 FILLER_150_1305 ();
 sg13g2_fill_2 FILLER_150_1310 ();
 sg13g2_fill_1 FILLER_150_1312 ();
 sg13g2_fill_1 FILLER_150_1317 ();
 sg13g2_decap_8 FILLER_150_1331 ();
 sg13g2_fill_2 FILLER_150_1346 ();
 sg13g2_decap_8 FILLER_150_1356 ();
 sg13g2_decap_8 FILLER_150_1363 ();
 sg13g2_decap_8 FILLER_150_1370 ();
 sg13g2_fill_2 FILLER_150_1377 ();
 sg13g2_decap_8 FILLER_150_1394 ();
 sg13g2_decap_8 FILLER_150_1401 ();
 sg13g2_decap_8 FILLER_150_1408 ();
 sg13g2_decap_8 FILLER_150_1415 ();
 sg13g2_decap_8 FILLER_150_1432 ();
 sg13g2_decap_4 FILLER_150_1439 ();
 sg13g2_fill_1 FILLER_150_1443 ();
 sg13g2_decap_8 FILLER_150_1452 ();
 sg13g2_decap_8 FILLER_150_1459 ();
 sg13g2_decap_8 FILLER_150_1474 ();
 sg13g2_decap_8 FILLER_150_1481 ();
 sg13g2_decap_8 FILLER_150_1488 ();
 sg13g2_decap_8 FILLER_150_1495 ();
 sg13g2_decap_8 FILLER_150_1502 ();
 sg13g2_decap_4 FILLER_150_1509 ();
 sg13g2_fill_2 FILLER_150_1513 ();
 sg13g2_fill_2 FILLER_150_1523 ();
 sg13g2_fill_1 FILLER_150_1533 ();
 sg13g2_decap_8 FILLER_150_1558 ();
 sg13g2_decap_8 FILLER_150_1565 ();
 sg13g2_decap_4 FILLER_150_1572 ();
 sg13g2_fill_1 FILLER_150_1576 ();
 sg13g2_fill_2 FILLER_150_1582 ();
 sg13g2_fill_1 FILLER_150_1584 ();
 sg13g2_decap_8 FILLER_150_1603 ();
 sg13g2_decap_8 FILLER_150_1610 ();
 sg13g2_decap_8 FILLER_150_1617 ();
 sg13g2_decap_8 FILLER_150_1624 ();
 sg13g2_decap_8 FILLER_150_1631 ();
 sg13g2_decap_8 FILLER_150_1638 ();
 sg13g2_decap_8 FILLER_150_1645 ();
 sg13g2_decap_8 FILLER_150_1652 ();
 sg13g2_decap_8 FILLER_150_1659 ();
 sg13g2_decap_8 FILLER_150_1666 ();
 sg13g2_decap_8 FILLER_150_1673 ();
 sg13g2_decap_8 FILLER_150_1680 ();
 sg13g2_decap_8 FILLER_150_1687 ();
 sg13g2_decap_8 FILLER_150_1694 ();
 sg13g2_decap_8 FILLER_150_1701 ();
 sg13g2_decap_8 FILLER_150_1708 ();
 sg13g2_decap_8 FILLER_150_1715 ();
 sg13g2_decap_8 FILLER_150_1722 ();
 sg13g2_decap_8 FILLER_150_1729 ();
 sg13g2_decap_8 FILLER_150_1736 ();
 sg13g2_decap_8 FILLER_150_1743 ();
 sg13g2_decap_8 FILLER_150_1750 ();
 sg13g2_decap_8 FILLER_150_1757 ();
 sg13g2_decap_4 FILLER_150_1764 ();
 sg13g2_decap_8 FILLER_151_0 ();
 sg13g2_decap_8 FILLER_151_7 ();
 sg13g2_decap_8 FILLER_151_14 ();
 sg13g2_fill_2 FILLER_151_21 ();
 sg13g2_fill_2 FILLER_151_30 ();
 sg13g2_fill_1 FILLER_151_32 ();
 sg13g2_decap_8 FILLER_151_51 ();
 sg13g2_decap_8 FILLER_151_58 ();
 sg13g2_decap_8 FILLER_151_65 ();
 sg13g2_decap_8 FILLER_151_72 ();
 sg13g2_decap_8 FILLER_151_79 ();
 sg13g2_decap_8 FILLER_151_86 ();
 sg13g2_fill_2 FILLER_151_93 ();
 sg13g2_fill_1 FILLER_151_95 ();
 sg13g2_decap_8 FILLER_151_123 ();
 sg13g2_decap_8 FILLER_151_130 ();
 sg13g2_fill_1 FILLER_151_137 ();
 sg13g2_fill_2 FILLER_151_149 ();
 sg13g2_decap_8 FILLER_151_161 ();
 sg13g2_decap_8 FILLER_151_168 ();
 sg13g2_decap_8 FILLER_151_175 ();
 sg13g2_decap_8 FILLER_151_182 ();
 sg13g2_decap_8 FILLER_151_189 ();
 sg13g2_decap_8 FILLER_151_196 ();
 sg13g2_decap_8 FILLER_151_203 ();
 sg13g2_decap_8 FILLER_151_210 ();
 sg13g2_decap_8 FILLER_151_217 ();
 sg13g2_decap_8 FILLER_151_224 ();
 sg13g2_decap_8 FILLER_151_231 ();
 sg13g2_decap_8 FILLER_151_238 ();
 sg13g2_decap_8 FILLER_151_245 ();
 sg13g2_decap_8 FILLER_151_252 ();
 sg13g2_decap_8 FILLER_151_259 ();
 sg13g2_decap_8 FILLER_151_266 ();
 sg13g2_decap_4 FILLER_151_273 ();
 sg13g2_decap_8 FILLER_151_285 ();
 sg13g2_decap_8 FILLER_151_292 ();
 sg13g2_decap_8 FILLER_151_299 ();
 sg13g2_decap_8 FILLER_151_306 ();
 sg13g2_decap_8 FILLER_151_313 ();
 sg13g2_decap_4 FILLER_151_320 ();
 sg13g2_fill_2 FILLER_151_324 ();
 sg13g2_decap_8 FILLER_151_330 ();
 sg13g2_fill_2 FILLER_151_337 ();
 sg13g2_decap_8 FILLER_151_344 ();
 sg13g2_decap_8 FILLER_151_351 ();
 sg13g2_decap_8 FILLER_151_358 ();
 sg13g2_decap_8 FILLER_151_365 ();
 sg13g2_decap_8 FILLER_151_372 ();
 sg13g2_fill_1 FILLER_151_379 ();
 sg13g2_fill_1 FILLER_151_388 ();
 sg13g2_decap_8 FILLER_151_399 ();
 sg13g2_decap_8 FILLER_151_406 ();
 sg13g2_decap_8 FILLER_151_413 ();
 sg13g2_decap_8 FILLER_151_420 ();
 sg13g2_decap_8 FILLER_151_427 ();
 sg13g2_decap_4 FILLER_151_434 ();
 sg13g2_fill_2 FILLER_151_438 ();
 sg13g2_fill_2 FILLER_151_448 ();
 sg13g2_decap_8 FILLER_151_468 ();
 sg13g2_decap_8 FILLER_151_475 ();
 sg13g2_fill_1 FILLER_151_486 ();
 sg13g2_decap_8 FILLER_151_498 ();
 sg13g2_decap_8 FILLER_151_505 ();
 sg13g2_decap_8 FILLER_151_512 ();
 sg13g2_decap_8 FILLER_151_519 ();
 sg13g2_decap_8 FILLER_151_526 ();
 sg13g2_decap_8 FILLER_151_533 ();
 sg13g2_decap_8 FILLER_151_540 ();
 sg13g2_decap_8 FILLER_151_547 ();
 sg13g2_decap_8 FILLER_151_554 ();
 sg13g2_decap_8 FILLER_151_561 ();
 sg13g2_decap_8 FILLER_151_568 ();
 sg13g2_decap_8 FILLER_151_575 ();
 sg13g2_decap_8 FILLER_151_590 ();
 sg13g2_decap_8 FILLER_151_597 ();
 sg13g2_decap_8 FILLER_151_604 ();
 sg13g2_decap_8 FILLER_151_611 ();
 sg13g2_decap_8 FILLER_151_618 ();
 sg13g2_fill_2 FILLER_151_625 ();
 sg13g2_fill_1 FILLER_151_627 ();
 sg13g2_decap_4 FILLER_151_638 ();
 sg13g2_decap_4 FILLER_151_655 ();
 sg13g2_fill_1 FILLER_151_659 ();
 sg13g2_decap_8 FILLER_151_668 ();
 sg13g2_decap_8 FILLER_151_675 ();
 sg13g2_decap_8 FILLER_151_682 ();
 sg13g2_decap_8 FILLER_151_702 ();
 sg13g2_decap_8 FILLER_151_709 ();
 sg13g2_decap_8 FILLER_151_716 ();
 sg13g2_decap_8 FILLER_151_723 ();
 sg13g2_decap_8 FILLER_151_730 ();
 sg13g2_decap_8 FILLER_151_737 ();
 sg13g2_fill_2 FILLER_151_744 ();
 sg13g2_decap_8 FILLER_151_759 ();
 sg13g2_decap_8 FILLER_151_766 ();
 sg13g2_decap_8 FILLER_151_773 ();
 sg13g2_decap_8 FILLER_151_780 ();
 sg13g2_decap_4 FILLER_151_787 ();
 sg13g2_decap_8 FILLER_151_795 ();
 sg13g2_decap_8 FILLER_151_802 ();
 sg13g2_decap_8 FILLER_151_809 ();
 sg13g2_decap_8 FILLER_151_816 ();
 sg13g2_decap_8 FILLER_151_823 ();
 sg13g2_decap_4 FILLER_151_830 ();
 sg13g2_fill_2 FILLER_151_860 ();
 sg13g2_fill_1 FILLER_151_862 ();
 sg13g2_decap_8 FILLER_151_872 ();
 sg13g2_decap_8 FILLER_151_879 ();
 sg13g2_decap_8 FILLER_151_886 ();
 sg13g2_fill_2 FILLER_151_893 ();
 sg13g2_decap_8 FILLER_151_911 ();
 sg13g2_decap_8 FILLER_151_918 ();
 sg13g2_decap_8 FILLER_151_925 ();
 sg13g2_decap_4 FILLER_151_932 ();
 sg13g2_fill_1 FILLER_151_936 ();
 sg13g2_decap_8 FILLER_151_958 ();
 sg13g2_decap_4 FILLER_151_965 ();
 sg13g2_fill_1 FILLER_151_969 ();
 sg13g2_decap_8 FILLER_151_975 ();
 sg13g2_decap_8 FILLER_151_982 ();
 sg13g2_decap_8 FILLER_151_989 ();
 sg13g2_decap_8 FILLER_151_996 ();
 sg13g2_decap_8 FILLER_151_1003 ();
 sg13g2_fill_2 FILLER_151_1039 ();
 sg13g2_decap_8 FILLER_151_1049 ();
 sg13g2_decap_8 FILLER_151_1056 ();
 sg13g2_decap_8 FILLER_151_1063 ();
 sg13g2_fill_2 FILLER_151_1070 ();
 sg13g2_decap_8 FILLER_151_1103 ();
 sg13g2_fill_2 FILLER_151_1110 ();
 sg13g2_decap_4 FILLER_151_1124 ();
 sg13g2_fill_1 FILLER_151_1128 ();
 sg13g2_fill_1 FILLER_151_1134 ();
 sg13g2_decap_8 FILLER_151_1143 ();
 sg13g2_decap_8 FILLER_151_1150 ();
 sg13g2_decap_8 FILLER_151_1157 ();
 sg13g2_decap_8 FILLER_151_1164 ();
 sg13g2_fill_1 FILLER_151_1171 ();
 sg13g2_decap_8 FILLER_151_1186 ();
 sg13g2_decap_8 FILLER_151_1193 ();
 sg13g2_decap_4 FILLER_151_1200 ();
 sg13g2_fill_2 FILLER_151_1204 ();
 sg13g2_decap_8 FILLER_151_1214 ();
 sg13g2_decap_8 FILLER_151_1221 ();
 sg13g2_decap_8 FILLER_151_1228 ();
 sg13g2_decap_8 FILLER_151_1235 ();
 sg13g2_decap_8 FILLER_151_1242 ();
 sg13g2_decap_8 FILLER_151_1249 ();
 sg13g2_decap_8 FILLER_151_1256 ();
 sg13g2_decap_8 FILLER_151_1263 ();
 sg13g2_decap_8 FILLER_151_1270 ();
 sg13g2_decap_8 FILLER_151_1277 ();
 sg13g2_decap_8 FILLER_151_1284 ();
 sg13g2_decap_8 FILLER_151_1291 ();
 sg13g2_decap_8 FILLER_151_1298 ();
 sg13g2_fill_2 FILLER_151_1305 ();
 sg13g2_fill_2 FILLER_151_1319 ();
 sg13g2_decap_8 FILLER_151_1329 ();
 sg13g2_decap_8 FILLER_151_1336 ();
 sg13g2_fill_1 FILLER_151_1343 ();
 sg13g2_decap_8 FILLER_151_1349 ();
 sg13g2_decap_8 FILLER_151_1356 ();
 sg13g2_decap_8 FILLER_151_1363 ();
 sg13g2_decap_8 FILLER_151_1370 ();
 sg13g2_decap_8 FILLER_151_1377 ();
 sg13g2_decap_8 FILLER_151_1384 ();
 sg13g2_decap_8 FILLER_151_1391 ();
 sg13g2_decap_8 FILLER_151_1398 ();
 sg13g2_decap_8 FILLER_151_1405 ();
 sg13g2_decap_8 FILLER_151_1412 ();
 sg13g2_decap_4 FILLER_151_1419 ();
 sg13g2_fill_2 FILLER_151_1423 ();
 sg13g2_decap_8 FILLER_151_1438 ();
 sg13g2_decap_8 FILLER_151_1445 ();
 sg13g2_decap_8 FILLER_151_1452 ();
 sg13g2_decap_4 FILLER_151_1459 ();
 sg13g2_fill_1 FILLER_151_1463 ();
 sg13g2_decap_8 FILLER_151_1472 ();
 sg13g2_decap_8 FILLER_151_1479 ();
 sg13g2_decap_8 FILLER_151_1486 ();
 sg13g2_decap_8 FILLER_151_1493 ();
 sg13g2_decap_4 FILLER_151_1500 ();
 sg13g2_fill_1 FILLER_151_1504 ();
 sg13g2_fill_1 FILLER_151_1510 ();
 sg13g2_decap_8 FILLER_151_1515 ();
 sg13g2_fill_2 FILLER_151_1522 ();
 sg13g2_fill_1 FILLER_151_1524 ();
 sg13g2_fill_2 FILLER_151_1529 ();
 sg13g2_decap_8 FILLER_151_1536 ();
 sg13g2_decap_8 FILLER_151_1543 ();
 sg13g2_fill_2 FILLER_151_1550 ();
 sg13g2_decap_8 FILLER_151_1556 ();
 sg13g2_decap_8 FILLER_151_1563 ();
 sg13g2_fill_2 FILLER_151_1570 ();
 sg13g2_fill_1 FILLER_151_1588 ();
 sg13g2_decap_8 FILLER_151_1604 ();
 sg13g2_decap_8 FILLER_151_1611 ();
 sg13g2_decap_8 FILLER_151_1618 ();
 sg13g2_decap_8 FILLER_151_1625 ();
 sg13g2_decap_8 FILLER_151_1632 ();
 sg13g2_decap_8 FILLER_151_1639 ();
 sg13g2_decap_8 FILLER_151_1646 ();
 sg13g2_decap_8 FILLER_151_1653 ();
 sg13g2_decap_8 FILLER_151_1660 ();
 sg13g2_decap_8 FILLER_151_1667 ();
 sg13g2_decap_8 FILLER_151_1674 ();
 sg13g2_decap_8 FILLER_151_1681 ();
 sg13g2_decap_8 FILLER_151_1688 ();
 sg13g2_decap_8 FILLER_151_1695 ();
 sg13g2_decap_8 FILLER_151_1702 ();
 sg13g2_decap_8 FILLER_151_1709 ();
 sg13g2_decap_8 FILLER_151_1716 ();
 sg13g2_decap_8 FILLER_151_1723 ();
 sg13g2_decap_8 FILLER_151_1730 ();
 sg13g2_decap_8 FILLER_151_1737 ();
 sg13g2_decap_8 FILLER_151_1744 ();
 sg13g2_decap_8 FILLER_151_1751 ();
 sg13g2_decap_8 FILLER_151_1758 ();
 sg13g2_fill_2 FILLER_151_1765 ();
 sg13g2_fill_1 FILLER_151_1767 ();
 sg13g2_decap_8 FILLER_152_0 ();
 sg13g2_decap_8 FILLER_152_7 ();
 sg13g2_decap_8 FILLER_152_14 ();
 sg13g2_decap_8 FILLER_152_21 ();
 sg13g2_decap_4 FILLER_152_28 ();
 sg13g2_fill_2 FILLER_152_37 ();
 sg13g2_decap_8 FILLER_152_55 ();
 sg13g2_decap_8 FILLER_152_62 ();
 sg13g2_decap_8 FILLER_152_69 ();
 sg13g2_decap_4 FILLER_152_76 ();
 sg13g2_fill_2 FILLER_152_80 ();
 sg13g2_decap_8 FILLER_152_91 ();
 sg13g2_decap_8 FILLER_152_98 ();
 sg13g2_decap_8 FILLER_152_105 ();
 sg13g2_decap_8 FILLER_152_112 ();
 sg13g2_decap_8 FILLER_152_119 ();
 sg13g2_fill_2 FILLER_152_140 ();
 sg13g2_decap_8 FILLER_152_154 ();
 sg13g2_decap_8 FILLER_152_161 ();
 sg13g2_fill_2 FILLER_152_168 ();
 sg13g2_decap_8 FILLER_152_180 ();
 sg13g2_decap_4 FILLER_152_187 ();
 sg13g2_fill_1 FILLER_152_191 ();
 sg13g2_decap_8 FILLER_152_205 ();
 sg13g2_decap_8 FILLER_152_248 ();
 sg13g2_decap_8 FILLER_152_255 ();
 sg13g2_fill_2 FILLER_152_262 ();
 sg13g2_fill_1 FILLER_152_264 ();
 sg13g2_decap_8 FILLER_152_278 ();
 sg13g2_decap_8 FILLER_152_285 ();
 sg13g2_decap_8 FILLER_152_292 ();
 sg13g2_decap_4 FILLER_152_299 ();
 sg13g2_fill_1 FILLER_152_303 ();
 sg13g2_decap_8 FILLER_152_309 ();
 sg13g2_decap_8 FILLER_152_316 ();
 sg13g2_decap_8 FILLER_152_328 ();
 sg13g2_decap_8 FILLER_152_335 ();
 sg13g2_decap_8 FILLER_152_342 ();
 sg13g2_decap_8 FILLER_152_349 ();
 sg13g2_decap_8 FILLER_152_356 ();
 sg13g2_decap_8 FILLER_152_363 ();
 sg13g2_decap_8 FILLER_152_370 ();
 sg13g2_decap_8 FILLER_152_377 ();
 sg13g2_fill_2 FILLER_152_384 ();
 sg13g2_decap_8 FILLER_152_394 ();
 sg13g2_fill_2 FILLER_152_401 ();
 sg13g2_fill_1 FILLER_152_407 ();
 sg13g2_fill_1 FILLER_152_411 ();
 sg13g2_decap_8 FILLER_152_429 ();
 sg13g2_decap_8 FILLER_152_436 ();
 sg13g2_fill_2 FILLER_152_443 ();
 sg13g2_fill_1 FILLER_152_445 ();
 sg13g2_decap_8 FILLER_152_463 ();
 sg13g2_decap_8 FILLER_152_470 ();
 sg13g2_decap_8 FILLER_152_477 ();
 sg13g2_decap_8 FILLER_152_484 ();
 sg13g2_fill_2 FILLER_152_491 ();
 sg13g2_fill_1 FILLER_152_493 ();
 sg13g2_decap_8 FILLER_152_511 ();
 sg13g2_decap_8 FILLER_152_518 ();
 sg13g2_fill_1 FILLER_152_525 ();
 sg13g2_decap_8 FILLER_152_535 ();
 sg13g2_decap_8 FILLER_152_542 ();
 sg13g2_decap_8 FILLER_152_549 ();
 sg13g2_decap_8 FILLER_152_556 ();
 sg13g2_decap_8 FILLER_152_563 ();
 sg13g2_decap_8 FILLER_152_570 ();
 sg13g2_decap_8 FILLER_152_577 ();
 sg13g2_decap_8 FILLER_152_584 ();
 sg13g2_decap_8 FILLER_152_591 ();
 sg13g2_decap_8 FILLER_152_602 ();
 sg13g2_decap_8 FILLER_152_609 ();
 sg13g2_decap_8 FILLER_152_616 ();
 sg13g2_decap_8 FILLER_152_623 ();
 sg13g2_decap_8 FILLER_152_630 ();
 sg13g2_decap_8 FILLER_152_637 ();
 sg13g2_decap_8 FILLER_152_644 ();
 sg13g2_fill_2 FILLER_152_651 ();
 sg13g2_fill_1 FILLER_152_653 ();
 sg13g2_decap_8 FILLER_152_659 ();
 sg13g2_decap_8 FILLER_152_666 ();
 sg13g2_decap_8 FILLER_152_673 ();
 sg13g2_decap_8 FILLER_152_680 ();
 sg13g2_decap_8 FILLER_152_695 ();
 sg13g2_decap_8 FILLER_152_702 ();
 sg13g2_decap_8 FILLER_152_709 ();
 sg13g2_decap_8 FILLER_152_716 ();
 sg13g2_decap_8 FILLER_152_723 ();
 sg13g2_decap_8 FILLER_152_730 ();
 sg13g2_decap_8 FILLER_152_737 ();
 sg13g2_decap_8 FILLER_152_744 ();
 sg13g2_decap_8 FILLER_152_751 ();
 sg13g2_decap_8 FILLER_152_758 ();
 sg13g2_decap_8 FILLER_152_765 ();
 sg13g2_decap_8 FILLER_152_772 ();
 sg13g2_fill_2 FILLER_152_779 ();
 sg13g2_fill_1 FILLER_152_781 ();
 sg13g2_decap_8 FILLER_152_786 ();
 sg13g2_decap_8 FILLER_152_793 ();
 sg13g2_decap_8 FILLER_152_800 ();
 sg13g2_decap_4 FILLER_152_807 ();
 sg13g2_decap_8 FILLER_152_819 ();
 sg13g2_decap_8 FILLER_152_826 ();
 sg13g2_decap_8 FILLER_152_833 ();
 sg13g2_fill_1 FILLER_152_840 ();
 sg13g2_decap_8 FILLER_152_846 ();
 sg13g2_decap_8 FILLER_152_853 ();
 sg13g2_decap_8 FILLER_152_860 ();
 sg13g2_decap_8 FILLER_152_867 ();
 sg13g2_decap_8 FILLER_152_874 ();
 sg13g2_decap_8 FILLER_152_881 ();
 sg13g2_decap_8 FILLER_152_888 ();
 sg13g2_decap_8 FILLER_152_895 ();
 sg13g2_decap_8 FILLER_152_902 ();
 sg13g2_fill_2 FILLER_152_909 ();
 sg13g2_decap_8 FILLER_152_923 ();
 sg13g2_fill_2 FILLER_152_930 ();
 sg13g2_decap_8 FILLER_152_939 ();
 sg13g2_decap_8 FILLER_152_946 ();
 sg13g2_decap_8 FILLER_152_953 ();
 sg13g2_decap_8 FILLER_152_960 ();
 sg13g2_decap_4 FILLER_152_967 ();
 sg13g2_fill_2 FILLER_152_971 ();
 sg13g2_decap_8 FILLER_152_981 ();
 sg13g2_decap_8 FILLER_152_988 ();
 sg13g2_decap_8 FILLER_152_995 ();
 sg13g2_fill_1 FILLER_152_1002 ();
 sg13g2_decap_8 FILLER_152_1012 ();
 sg13g2_decap_8 FILLER_152_1019 ();
 sg13g2_decap_8 FILLER_152_1026 ();
 sg13g2_decap_8 FILLER_152_1033 ();
 sg13g2_decap_8 FILLER_152_1040 ();
 sg13g2_decap_8 FILLER_152_1047 ();
 sg13g2_decap_8 FILLER_152_1054 ();
 sg13g2_decap_8 FILLER_152_1061 ();
 sg13g2_decap_8 FILLER_152_1068 ();
 sg13g2_decap_4 FILLER_152_1075 ();
 sg13g2_fill_1 FILLER_152_1084 ();
 sg13g2_fill_2 FILLER_152_1092 ();
 sg13g2_fill_1 FILLER_152_1094 ();
 sg13g2_decap_8 FILLER_152_1108 ();
 sg13g2_decap_8 FILLER_152_1115 ();
 sg13g2_decap_4 FILLER_152_1122 ();
 sg13g2_fill_2 FILLER_152_1131 ();
 sg13g2_decap_8 FILLER_152_1149 ();
 sg13g2_decap_8 FILLER_152_1156 ();
 sg13g2_decap_8 FILLER_152_1163 ();
 sg13g2_decap_8 FILLER_152_1170 ();
 sg13g2_fill_2 FILLER_152_1177 ();
 sg13g2_decap_8 FILLER_152_1187 ();
 sg13g2_decap_8 FILLER_152_1194 ();
 sg13g2_decap_4 FILLER_152_1201 ();
 sg13g2_fill_2 FILLER_152_1205 ();
 sg13g2_decap_8 FILLER_152_1215 ();
 sg13g2_decap_8 FILLER_152_1222 ();
 sg13g2_decap_8 FILLER_152_1229 ();
 sg13g2_decap_8 FILLER_152_1236 ();
 sg13g2_decap_8 FILLER_152_1243 ();
 sg13g2_decap_8 FILLER_152_1250 ();
 sg13g2_decap_4 FILLER_152_1257 ();
 sg13g2_decap_8 FILLER_152_1265 ();
 sg13g2_decap_8 FILLER_152_1272 ();
 sg13g2_fill_2 FILLER_152_1279 ();
 sg13g2_fill_1 FILLER_152_1281 ();
 sg13g2_decap_8 FILLER_152_1287 ();
 sg13g2_decap_8 FILLER_152_1294 ();
 sg13g2_decap_8 FILLER_152_1301 ();
 sg13g2_decap_8 FILLER_152_1308 ();
 sg13g2_decap_8 FILLER_152_1315 ();
 sg13g2_decap_8 FILLER_152_1322 ();
 sg13g2_decap_8 FILLER_152_1329 ();
 sg13g2_decap_8 FILLER_152_1336 ();
 sg13g2_decap_8 FILLER_152_1343 ();
 sg13g2_decap_8 FILLER_152_1350 ();
 sg13g2_decap_8 FILLER_152_1357 ();
 sg13g2_decap_8 FILLER_152_1364 ();
 sg13g2_decap_8 FILLER_152_1371 ();
 sg13g2_decap_8 FILLER_152_1378 ();
 sg13g2_fill_1 FILLER_152_1385 ();
 sg13g2_decap_8 FILLER_152_1391 ();
 sg13g2_decap_8 FILLER_152_1398 ();
 sg13g2_decap_8 FILLER_152_1405 ();
 sg13g2_decap_8 FILLER_152_1412 ();
 sg13g2_fill_2 FILLER_152_1419 ();
 sg13g2_fill_2 FILLER_152_1426 ();
 sg13g2_decap_8 FILLER_152_1437 ();
 sg13g2_decap_8 FILLER_152_1444 ();
 sg13g2_decap_8 FILLER_152_1451 ();
 sg13g2_decap_8 FILLER_152_1458 ();
 sg13g2_decap_8 FILLER_152_1465 ();
 sg13g2_decap_8 FILLER_152_1472 ();
 sg13g2_decap_8 FILLER_152_1479 ();
 sg13g2_decap_8 FILLER_152_1486 ();
 sg13g2_decap_8 FILLER_152_1493 ();
 sg13g2_decap_8 FILLER_152_1500 ();
 sg13g2_decap_4 FILLER_152_1507 ();
 sg13g2_fill_2 FILLER_152_1511 ();
 sg13g2_decap_4 FILLER_152_1521 ();
 sg13g2_fill_1 FILLER_152_1525 ();
 sg13g2_decap_8 FILLER_152_1534 ();
 sg13g2_decap_8 FILLER_152_1541 ();
 sg13g2_decap_8 FILLER_152_1548 ();
 sg13g2_decap_8 FILLER_152_1555 ();
 sg13g2_decap_8 FILLER_152_1562 ();
 sg13g2_decap_8 FILLER_152_1569 ();
 sg13g2_decap_8 FILLER_152_1576 ();
 sg13g2_fill_2 FILLER_152_1583 ();
 sg13g2_fill_1 FILLER_152_1585 ();
 sg13g2_decap_8 FILLER_152_1598 ();
 sg13g2_decap_8 FILLER_152_1605 ();
 sg13g2_decap_8 FILLER_152_1612 ();
 sg13g2_decap_8 FILLER_152_1619 ();
 sg13g2_decap_8 FILLER_152_1626 ();
 sg13g2_decap_8 FILLER_152_1633 ();
 sg13g2_decap_8 FILLER_152_1640 ();
 sg13g2_decap_8 FILLER_152_1647 ();
 sg13g2_decap_8 FILLER_152_1654 ();
 sg13g2_decap_8 FILLER_152_1661 ();
 sg13g2_decap_8 FILLER_152_1668 ();
 sg13g2_decap_8 FILLER_152_1675 ();
 sg13g2_decap_8 FILLER_152_1682 ();
 sg13g2_decap_8 FILLER_152_1689 ();
 sg13g2_decap_8 FILLER_152_1696 ();
 sg13g2_decap_8 FILLER_152_1703 ();
 sg13g2_decap_8 FILLER_152_1710 ();
 sg13g2_decap_8 FILLER_152_1717 ();
 sg13g2_decap_8 FILLER_152_1724 ();
 sg13g2_decap_8 FILLER_152_1731 ();
 sg13g2_decap_8 FILLER_152_1738 ();
 sg13g2_decap_8 FILLER_152_1745 ();
 sg13g2_decap_8 FILLER_152_1752 ();
 sg13g2_decap_8 FILLER_152_1759 ();
 sg13g2_fill_2 FILLER_152_1766 ();
 sg13g2_decap_8 FILLER_153_0 ();
 sg13g2_decap_8 FILLER_153_7 ();
 sg13g2_decap_8 FILLER_153_14 ();
 sg13g2_fill_1 FILLER_153_34 ();
 sg13g2_decap_8 FILLER_153_56 ();
 sg13g2_decap_8 FILLER_153_63 ();
 sg13g2_decap_8 FILLER_153_70 ();
 sg13g2_decap_4 FILLER_153_77 ();
 sg13g2_fill_1 FILLER_153_81 ();
 sg13g2_decap_8 FILLER_153_94 ();
 sg13g2_decap_8 FILLER_153_101 ();
 sg13g2_decap_8 FILLER_153_108 ();
 sg13g2_fill_2 FILLER_153_115 ();
 sg13g2_fill_1 FILLER_153_117 ();
 sg13g2_decap_4 FILLER_153_135 ();
 sg13g2_decap_8 FILLER_153_143 ();
 sg13g2_decap_8 FILLER_153_150 ();
 sg13g2_decap_8 FILLER_153_157 ();
 sg13g2_fill_2 FILLER_153_164 ();
 sg13g2_fill_1 FILLER_153_166 ();
 sg13g2_decap_8 FILLER_153_201 ();
 sg13g2_decap_8 FILLER_153_208 ();
 sg13g2_decap_8 FILLER_153_215 ();
 sg13g2_decap_8 FILLER_153_222 ();
 sg13g2_decap_4 FILLER_153_229 ();
 sg13g2_decap_8 FILLER_153_237 ();
 sg13g2_fill_2 FILLER_153_244 ();
 sg13g2_fill_1 FILLER_153_246 ();
 sg13g2_fill_2 FILLER_153_273 ();
 sg13g2_fill_1 FILLER_153_275 ();
 sg13g2_decap_8 FILLER_153_289 ();
 sg13g2_decap_8 FILLER_153_296 ();
 sg13g2_decap_8 FILLER_153_303 ();
 sg13g2_decap_4 FILLER_153_310 ();
 sg13g2_fill_1 FILLER_153_314 ();
 sg13g2_decap_8 FILLER_153_320 ();
 sg13g2_decap_8 FILLER_153_365 ();
 sg13g2_decap_8 FILLER_153_372 ();
 sg13g2_decap_8 FILLER_153_379 ();
 sg13g2_decap_8 FILLER_153_386 ();
 sg13g2_decap_4 FILLER_153_393 ();
 sg13g2_fill_2 FILLER_153_397 ();
 sg13g2_decap_8 FILLER_153_424 ();
 sg13g2_decap_8 FILLER_153_431 ();
 sg13g2_decap_8 FILLER_153_438 ();
 sg13g2_decap_8 FILLER_153_445 ();
 sg13g2_fill_1 FILLER_153_452 ();
 sg13g2_decap_8 FILLER_153_471 ();
 sg13g2_decap_8 FILLER_153_478 ();
 sg13g2_decap_8 FILLER_153_485 ();
 sg13g2_decap_8 FILLER_153_492 ();
 sg13g2_decap_4 FILLER_153_499 ();
 sg13g2_fill_2 FILLER_153_503 ();
 sg13g2_decap_4 FILLER_153_514 ();
 sg13g2_fill_1 FILLER_153_518 ();
 sg13g2_decap_8 FILLER_153_543 ();
 sg13g2_decap_8 FILLER_153_550 ();
 sg13g2_fill_2 FILLER_153_560 ();
 sg13g2_decap_8 FILLER_153_566 ();
 sg13g2_decap_8 FILLER_153_573 ();
 sg13g2_decap_8 FILLER_153_580 ();
 sg13g2_decap_8 FILLER_153_587 ();
 sg13g2_decap_4 FILLER_153_594 ();
 sg13g2_fill_1 FILLER_153_598 ();
 sg13g2_decap_8 FILLER_153_618 ();
 sg13g2_decap_4 FILLER_153_625 ();
 sg13g2_decap_8 FILLER_153_642 ();
 sg13g2_fill_1 FILLER_153_649 ();
 sg13g2_fill_1 FILLER_153_658 ();
 sg13g2_fill_1 FILLER_153_679 ();
 sg13g2_decap_8 FILLER_153_688 ();
 sg13g2_decap_4 FILLER_153_695 ();
 sg13g2_decap_8 FILLER_153_716 ();
 sg13g2_decap_8 FILLER_153_723 ();
 sg13g2_decap_8 FILLER_153_730 ();
 sg13g2_decap_8 FILLER_153_737 ();
 sg13g2_decap_8 FILLER_153_744 ();
 sg13g2_decap_8 FILLER_153_751 ();
 sg13g2_decap_8 FILLER_153_758 ();
 sg13g2_decap_8 FILLER_153_765 ();
 sg13g2_fill_2 FILLER_153_772 ();
 sg13g2_fill_1 FILLER_153_782 ();
 sg13g2_decap_8 FILLER_153_796 ();
 sg13g2_fill_2 FILLER_153_803 ();
 sg13g2_decap_8 FILLER_153_811 ();
 sg13g2_decap_8 FILLER_153_835 ();
 sg13g2_fill_2 FILLER_153_842 ();
 sg13g2_decap_8 FILLER_153_847 ();
 sg13g2_decap_8 FILLER_153_854 ();
 sg13g2_decap_8 FILLER_153_861 ();
 sg13g2_decap_8 FILLER_153_868 ();
 sg13g2_decap_8 FILLER_153_875 ();
 sg13g2_fill_2 FILLER_153_882 ();
 sg13g2_fill_1 FILLER_153_884 ();
 sg13g2_decap_8 FILLER_153_947 ();
 sg13g2_decap_4 FILLER_153_954 ();
 sg13g2_decap_8 FILLER_153_968 ();
 sg13g2_decap_8 FILLER_153_975 ();
 sg13g2_decap_8 FILLER_153_982 ();
 sg13g2_decap_8 FILLER_153_989 ();
 sg13g2_decap_4 FILLER_153_996 ();
 sg13g2_decap_8 FILLER_153_1011 ();
 sg13g2_decap_8 FILLER_153_1018 ();
 sg13g2_decap_8 FILLER_153_1025 ();
 sg13g2_decap_8 FILLER_153_1032 ();
 sg13g2_decap_8 FILLER_153_1039 ();
 sg13g2_fill_1 FILLER_153_1046 ();
 sg13g2_fill_1 FILLER_153_1055 ();
 sg13g2_decap_8 FILLER_153_1061 ();
 sg13g2_fill_2 FILLER_153_1068 ();
 sg13g2_decap_8 FILLER_153_1075 ();
 sg13g2_decap_8 FILLER_153_1082 ();
 sg13g2_decap_8 FILLER_153_1089 ();
 sg13g2_decap_8 FILLER_153_1096 ();
 sg13g2_decap_8 FILLER_153_1103 ();
 sg13g2_decap_8 FILLER_153_1110 ();
 sg13g2_decap_8 FILLER_153_1117 ();
 sg13g2_decap_8 FILLER_153_1124 ();
 sg13g2_decap_4 FILLER_153_1131 ();
 sg13g2_decap_8 FILLER_153_1140 ();
 sg13g2_fill_1 FILLER_153_1147 ();
 sg13g2_decap_8 FILLER_153_1156 ();
 sg13g2_decap_8 FILLER_153_1163 ();
 sg13g2_decap_8 FILLER_153_1170 ();
 sg13g2_decap_8 FILLER_153_1177 ();
 sg13g2_decap_8 FILLER_153_1184 ();
 sg13g2_decap_8 FILLER_153_1191 ();
 sg13g2_decap_4 FILLER_153_1198 ();
 sg13g2_decap_8 FILLER_153_1223 ();
 sg13g2_decap_8 FILLER_153_1230 ();
 sg13g2_decap_8 FILLER_153_1237 ();
 sg13g2_decap_8 FILLER_153_1244 ();
 sg13g2_decap_4 FILLER_153_1251 ();
 sg13g2_decap_8 FILLER_153_1272 ();
 sg13g2_decap_8 FILLER_153_1279 ();
 sg13g2_decap_8 FILLER_153_1286 ();
 sg13g2_decap_8 FILLER_153_1293 ();
 sg13g2_decap_8 FILLER_153_1300 ();
 sg13g2_fill_2 FILLER_153_1307 ();
 sg13g2_decap_8 FILLER_153_1325 ();
 sg13g2_decap_8 FILLER_153_1332 ();
 sg13g2_decap_4 FILLER_153_1339 ();
 sg13g2_fill_2 FILLER_153_1343 ();
 sg13g2_decap_8 FILLER_153_1355 ();
 sg13g2_decap_8 FILLER_153_1362 ();
 sg13g2_decap_8 FILLER_153_1369 ();
 sg13g2_decap_4 FILLER_153_1376 ();
 sg13g2_fill_2 FILLER_153_1380 ();
 sg13g2_decap_8 FILLER_153_1402 ();
 sg13g2_decap_8 FILLER_153_1409 ();
 sg13g2_decap_4 FILLER_153_1416 ();
 sg13g2_fill_1 FILLER_153_1420 ();
 sg13g2_decap_8 FILLER_153_1437 ();
 sg13g2_decap_8 FILLER_153_1444 ();
 sg13g2_decap_8 FILLER_153_1451 ();
 sg13g2_fill_2 FILLER_153_1458 ();
 sg13g2_fill_1 FILLER_153_1460 ();
 sg13g2_fill_1 FILLER_153_1469 ();
 sg13g2_decap_8 FILLER_153_1478 ();
 sg13g2_decap_8 FILLER_153_1485 ();
 sg13g2_decap_8 FILLER_153_1492 ();
 sg13g2_decap_8 FILLER_153_1499 ();
 sg13g2_decap_4 FILLER_153_1506 ();
 sg13g2_decap_8 FILLER_153_1532 ();
 sg13g2_decap_8 FILLER_153_1539 ();
 sg13g2_decap_8 FILLER_153_1546 ();
 sg13g2_decap_4 FILLER_153_1553 ();
 sg13g2_decap_8 FILLER_153_1570 ();
 sg13g2_decap_8 FILLER_153_1577 ();
 sg13g2_fill_1 FILLER_153_1584 ();
 sg13g2_decap_8 FILLER_153_1598 ();
 sg13g2_decap_8 FILLER_153_1605 ();
 sg13g2_decap_8 FILLER_153_1612 ();
 sg13g2_decap_8 FILLER_153_1619 ();
 sg13g2_decap_8 FILLER_153_1626 ();
 sg13g2_decap_8 FILLER_153_1633 ();
 sg13g2_decap_8 FILLER_153_1640 ();
 sg13g2_decap_8 FILLER_153_1647 ();
 sg13g2_decap_8 FILLER_153_1654 ();
 sg13g2_decap_8 FILLER_153_1661 ();
 sg13g2_decap_8 FILLER_153_1668 ();
 sg13g2_decap_8 FILLER_153_1675 ();
 sg13g2_decap_8 FILLER_153_1682 ();
 sg13g2_decap_8 FILLER_153_1689 ();
 sg13g2_decap_8 FILLER_153_1696 ();
 sg13g2_decap_8 FILLER_153_1703 ();
 sg13g2_decap_8 FILLER_153_1710 ();
 sg13g2_decap_8 FILLER_153_1717 ();
 sg13g2_decap_8 FILLER_153_1724 ();
 sg13g2_decap_8 FILLER_153_1731 ();
 sg13g2_decap_8 FILLER_153_1738 ();
 sg13g2_decap_8 FILLER_153_1745 ();
 sg13g2_decap_8 FILLER_153_1752 ();
 sg13g2_decap_8 FILLER_153_1759 ();
 sg13g2_fill_2 FILLER_153_1766 ();
 sg13g2_decap_8 FILLER_154_0 ();
 sg13g2_decap_8 FILLER_154_7 ();
 sg13g2_decap_8 FILLER_154_14 ();
 sg13g2_decap_4 FILLER_154_21 ();
 sg13g2_fill_1 FILLER_154_25 ();
 sg13g2_decap_8 FILLER_154_46 ();
 sg13g2_decap_8 FILLER_154_53 ();
 sg13g2_decap_8 FILLER_154_60 ();
 sg13g2_decap_4 FILLER_154_67 ();
 sg13g2_fill_2 FILLER_154_71 ();
 sg13g2_decap_8 FILLER_154_86 ();
 sg13g2_decap_8 FILLER_154_93 ();
 sg13g2_decap_8 FILLER_154_100 ();
 sg13g2_decap_4 FILLER_154_107 ();
 sg13g2_fill_2 FILLER_154_111 ();
 sg13g2_decap_8 FILLER_154_117 ();
 sg13g2_decap_8 FILLER_154_124 ();
 sg13g2_decap_8 FILLER_154_131 ();
 sg13g2_decap_8 FILLER_154_138 ();
 sg13g2_decap_8 FILLER_154_145 ();
 sg13g2_decap_8 FILLER_154_152 ();
 sg13g2_decap_8 FILLER_154_159 ();
 sg13g2_decap_8 FILLER_154_166 ();
 sg13g2_decap_4 FILLER_154_173 ();
 sg13g2_fill_1 FILLER_154_177 ();
 sg13g2_decap_8 FILLER_154_182 ();
 sg13g2_decap_8 FILLER_154_189 ();
 sg13g2_decap_8 FILLER_154_196 ();
 sg13g2_decap_8 FILLER_154_203 ();
 sg13g2_decap_8 FILLER_154_210 ();
 sg13g2_decap_8 FILLER_154_217 ();
 sg13g2_decap_8 FILLER_154_224 ();
 sg13g2_decap_4 FILLER_154_231 ();
 sg13g2_decap_8 FILLER_154_245 ();
 sg13g2_decap_4 FILLER_154_252 ();
 sg13g2_fill_2 FILLER_154_256 ();
 sg13g2_decap_8 FILLER_154_262 ();
 sg13g2_decap_8 FILLER_154_269 ();
 sg13g2_decap_8 FILLER_154_276 ();
 sg13g2_decap_8 FILLER_154_283 ();
 sg13g2_decap_4 FILLER_154_290 ();
 sg13g2_fill_2 FILLER_154_294 ();
 sg13g2_fill_1 FILLER_154_348 ();
 sg13g2_decap_8 FILLER_154_375 ();
 sg13g2_decap_8 FILLER_154_382 ();
 sg13g2_decap_8 FILLER_154_389 ();
 sg13g2_decap_8 FILLER_154_396 ();
 sg13g2_decap_8 FILLER_154_403 ();
 sg13g2_decap_8 FILLER_154_410 ();
 sg13g2_decap_8 FILLER_154_417 ();
 sg13g2_decap_8 FILLER_154_424 ();
 sg13g2_decap_8 FILLER_154_431 ();
 sg13g2_decap_8 FILLER_154_438 ();
 sg13g2_decap_8 FILLER_154_465 ();
 sg13g2_decap_8 FILLER_154_472 ();
 sg13g2_decap_8 FILLER_154_479 ();
 sg13g2_decap_8 FILLER_154_486 ();
 sg13g2_decap_8 FILLER_154_493 ();
 sg13g2_decap_8 FILLER_154_508 ();
 sg13g2_decap_4 FILLER_154_515 ();
 sg13g2_fill_1 FILLER_154_531 ();
 sg13g2_decap_8 FILLER_154_545 ();
 sg13g2_fill_2 FILLER_154_552 ();
 sg13g2_fill_2 FILLER_154_562 ();
 sg13g2_decap_8 FILLER_154_573 ();
 sg13g2_decap_4 FILLER_154_580 ();
 sg13g2_decap_8 FILLER_154_610 ();
 sg13g2_decap_8 FILLER_154_617 ();
 sg13g2_decap_8 FILLER_154_624 ();
 sg13g2_decap_8 FILLER_154_631 ();
 sg13g2_decap_8 FILLER_154_638 ();
 sg13g2_decap_8 FILLER_154_645 ();
 sg13g2_fill_1 FILLER_154_652 ();
 sg13g2_decap_8 FILLER_154_663 ();
 sg13g2_fill_2 FILLER_154_670 ();
 sg13g2_decap_8 FILLER_154_689 ();
 sg13g2_decap_8 FILLER_154_696 ();
 sg13g2_decap_8 FILLER_154_703 ();
 sg13g2_fill_2 FILLER_154_710 ();
 sg13g2_decap_8 FILLER_154_724 ();
 sg13g2_decap_8 FILLER_154_731 ();
 sg13g2_decap_8 FILLER_154_738 ();
 sg13g2_fill_1 FILLER_154_745 ();
 sg13g2_fill_2 FILLER_154_755 ();
 sg13g2_decap_8 FILLER_154_761 ();
 sg13g2_decap_8 FILLER_154_768 ();
 sg13g2_decap_8 FILLER_154_775 ();
 sg13g2_decap_8 FILLER_154_782 ();
 sg13g2_fill_2 FILLER_154_789 ();
 sg13g2_fill_1 FILLER_154_791 ();
 sg13g2_decap_8 FILLER_154_806 ();
 sg13g2_decap_4 FILLER_154_813 ();
 sg13g2_fill_1 FILLER_154_817 ();
 sg13g2_decap_8 FILLER_154_839 ();
 sg13g2_fill_2 FILLER_154_846 ();
 sg13g2_decap_8 FILLER_154_863 ();
 sg13g2_decap_8 FILLER_154_870 ();
 sg13g2_decap_8 FILLER_154_877 ();
 sg13g2_decap_8 FILLER_154_884 ();
 sg13g2_decap_8 FILLER_154_891 ();
 sg13g2_decap_8 FILLER_154_898 ();
 sg13g2_decap_8 FILLER_154_905 ();
 sg13g2_decap_4 FILLER_154_912 ();
 sg13g2_fill_1 FILLER_154_916 ();
 sg13g2_decap_8 FILLER_154_931 ();
 sg13g2_decap_8 FILLER_154_938 ();
 sg13g2_decap_8 FILLER_154_945 ();
 sg13g2_decap_8 FILLER_154_952 ();
 sg13g2_decap_8 FILLER_154_959 ();
 sg13g2_fill_1 FILLER_154_966 ();
 sg13g2_fill_1 FILLER_154_993 ();
 sg13g2_decap_4 FILLER_154_997 ();
 sg13g2_fill_2 FILLER_154_1001 ();
 sg13g2_fill_2 FILLER_154_1007 ();
 sg13g2_decap_8 FILLER_154_1017 ();
 sg13g2_decap_8 FILLER_154_1024 ();
 sg13g2_decap_8 FILLER_154_1031 ();
 sg13g2_decap_8 FILLER_154_1050 ();
 sg13g2_decap_8 FILLER_154_1057 ();
 sg13g2_decap_8 FILLER_154_1064 ();
 sg13g2_decap_8 FILLER_154_1071 ();
 sg13g2_decap_8 FILLER_154_1078 ();
 sg13g2_decap_8 FILLER_154_1085 ();
 sg13g2_decap_8 FILLER_154_1092 ();
 sg13g2_decap_4 FILLER_154_1099 ();
 sg13g2_fill_2 FILLER_154_1103 ();
 sg13g2_decap_4 FILLER_154_1114 ();
 sg13g2_fill_1 FILLER_154_1118 ();
 sg13g2_fill_2 FILLER_154_1123 ();
 sg13g2_fill_1 FILLER_154_1125 ();
 sg13g2_decap_8 FILLER_154_1143 ();
 sg13g2_decap_4 FILLER_154_1150 ();
 sg13g2_fill_2 FILLER_154_1154 ();
 sg13g2_decap_8 FILLER_154_1172 ();
 sg13g2_decap_8 FILLER_154_1179 ();
 sg13g2_decap_4 FILLER_154_1186 ();
 sg13g2_fill_2 FILLER_154_1190 ();
 sg13g2_fill_2 FILLER_154_1208 ();
 sg13g2_decap_8 FILLER_154_1217 ();
 sg13g2_decap_8 FILLER_154_1224 ();
 sg13g2_decap_8 FILLER_154_1231 ();
 sg13g2_decap_8 FILLER_154_1238 ();
 sg13g2_decap_8 FILLER_154_1245 ();
 sg13g2_decap_4 FILLER_154_1252 ();
 sg13g2_fill_2 FILLER_154_1256 ();
 sg13g2_decap_8 FILLER_154_1271 ();
 sg13g2_decap_8 FILLER_154_1278 ();
 sg13g2_decap_4 FILLER_154_1285 ();
 sg13g2_fill_2 FILLER_154_1289 ();
 sg13g2_decap_8 FILLER_154_1299 ();
 sg13g2_decap_8 FILLER_154_1306 ();
 sg13g2_decap_8 FILLER_154_1313 ();
 sg13g2_fill_1 FILLER_154_1320 ();
 sg13g2_decap_8 FILLER_154_1325 ();
 sg13g2_decap_8 FILLER_154_1332 ();
 sg13g2_fill_1 FILLER_154_1339 ();
 sg13g2_decap_8 FILLER_154_1359 ();
 sg13g2_decap_8 FILLER_154_1366 ();
 sg13g2_decap_8 FILLER_154_1373 ();
 sg13g2_decap_8 FILLER_154_1380 ();
 sg13g2_fill_1 FILLER_154_1387 ();
 sg13g2_decap_8 FILLER_154_1401 ();
 sg13g2_fill_1 FILLER_154_1408 ();
 sg13g2_decap_8 FILLER_154_1424 ();
 sg13g2_decap_8 FILLER_154_1431 ();
 sg13g2_decap_8 FILLER_154_1438 ();
 sg13g2_decap_8 FILLER_154_1445 ();
 sg13g2_decap_8 FILLER_154_1452 ();
 sg13g2_fill_2 FILLER_154_1459 ();
 sg13g2_fill_1 FILLER_154_1461 ();
 sg13g2_decap_8 FILLER_154_1486 ();
 sg13g2_decap_8 FILLER_154_1493 ();
 sg13g2_decap_8 FILLER_154_1500 ();
 sg13g2_decap_8 FILLER_154_1507 ();
 sg13g2_fill_2 FILLER_154_1514 ();
 sg13g2_decap_8 FILLER_154_1524 ();
 sg13g2_decap_8 FILLER_154_1531 ();
 sg13g2_decap_8 FILLER_154_1538 ();
 sg13g2_decap_8 FILLER_154_1545 ();
 sg13g2_fill_1 FILLER_154_1552 ();
 sg13g2_decap_8 FILLER_154_1569 ();
 sg13g2_fill_2 FILLER_154_1576 ();
 sg13g2_decap_8 FILLER_154_1586 ();
 sg13g2_decap_8 FILLER_154_1593 ();
 sg13g2_decap_8 FILLER_154_1600 ();
 sg13g2_decap_8 FILLER_154_1607 ();
 sg13g2_decap_8 FILLER_154_1614 ();
 sg13g2_decap_8 FILLER_154_1621 ();
 sg13g2_decap_8 FILLER_154_1628 ();
 sg13g2_decap_8 FILLER_154_1635 ();
 sg13g2_decap_8 FILLER_154_1642 ();
 sg13g2_decap_8 FILLER_154_1649 ();
 sg13g2_decap_8 FILLER_154_1656 ();
 sg13g2_decap_8 FILLER_154_1663 ();
 sg13g2_decap_8 FILLER_154_1670 ();
 sg13g2_decap_8 FILLER_154_1677 ();
 sg13g2_decap_8 FILLER_154_1684 ();
 sg13g2_decap_8 FILLER_154_1691 ();
 sg13g2_decap_8 FILLER_154_1698 ();
 sg13g2_decap_8 FILLER_154_1705 ();
 sg13g2_decap_8 FILLER_154_1712 ();
 sg13g2_decap_8 FILLER_154_1719 ();
 sg13g2_decap_8 FILLER_154_1726 ();
 sg13g2_decap_8 FILLER_154_1733 ();
 sg13g2_decap_8 FILLER_154_1740 ();
 sg13g2_decap_8 FILLER_154_1747 ();
 sg13g2_decap_8 FILLER_154_1754 ();
 sg13g2_decap_8 FILLER_154_1761 ();
 sg13g2_decap_8 FILLER_155_0 ();
 sg13g2_decap_8 FILLER_155_7 ();
 sg13g2_decap_4 FILLER_155_14 ();
 sg13g2_fill_2 FILLER_155_18 ();
 sg13g2_decap_8 FILLER_155_40 ();
 sg13g2_decap_8 FILLER_155_47 ();
 sg13g2_decap_8 FILLER_155_54 ();
 sg13g2_decap_8 FILLER_155_61 ();
 sg13g2_decap_4 FILLER_155_68 ();
 sg13g2_fill_2 FILLER_155_72 ();
 sg13g2_decap_8 FILLER_155_95 ();
 sg13g2_decap_8 FILLER_155_102 ();
 sg13g2_decap_8 FILLER_155_109 ();
 sg13g2_decap_8 FILLER_155_126 ();
 sg13g2_decap_8 FILLER_155_133 ();
 sg13g2_decap_4 FILLER_155_140 ();
 sg13g2_decap_8 FILLER_155_152 ();
 sg13g2_decap_8 FILLER_155_159 ();
 sg13g2_decap_8 FILLER_155_166 ();
 sg13g2_decap_8 FILLER_155_173 ();
 sg13g2_decap_8 FILLER_155_180 ();
 sg13g2_fill_2 FILLER_155_187 ();
 sg13g2_fill_1 FILLER_155_189 ();
 sg13g2_decap_4 FILLER_155_201 ();
 sg13g2_decap_8 FILLER_155_249 ();
 sg13g2_decap_8 FILLER_155_256 ();
 sg13g2_decap_8 FILLER_155_263 ();
 sg13g2_decap_8 FILLER_155_270 ();
 sg13g2_decap_8 FILLER_155_277 ();
 sg13g2_decap_8 FILLER_155_284 ();
 sg13g2_fill_2 FILLER_155_291 ();
 sg13g2_fill_1 FILLER_155_293 ();
 sg13g2_fill_2 FILLER_155_308 ();
 sg13g2_fill_1 FILLER_155_310 ();
 sg13g2_decap_8 FILLER_155_320 ();
 sg13g2_decap_4 FILLER_155_327 ();
 sg13g2_fill_2 FILLER_155_331 ();
 sg13g2_decap_8 FILLER_155_337 ();
 sg13g2_decap_8 FILLER_155_344 ();
 sg13g2_decap_8 FILLER_155_351 ();
 sg13g2_fill_2 FILLER_155_358 ();
 sg13g2_decap_8 FILLER_155_364 ();
 sg13g2_decap_8 FILLER_155_371 ();
 sg13g2_decap_8 FILLER_155_378 ();
 sg13g2_decap_8 FILLER_155_385 ();
 sg13g2_decap_8 FILLER_155_392 ();
 sg13g2_decap_8 FILLER_155_399 ();
 sg13g2_decap_4 FILLER_155_406 ();
 sg13g2_fill_2 FILLER_155_410 ();
 sg13g2_decap_8 FILLER_155_431 ();
 sg13g2_decap_8 FILLER_155_438 ();
 sg13g2_decap_8 FILLER_155_445 ();
 sg13g2_decap_4 FILLER_155_452 ();
 sg13g2_fill_1 FILLER_155_456 ();
 sg13g2_decap_8 FILLER_155_465 ();
 sg13g2_decap_8 FILLER_155_472 ();
 sg13g2_decap_8 FILLER_155_479 ();
 sg13g2_decap_8 FILLER_155_486 ();
 sg13g2_decap_8 FILLER_155_493 ();
 sg13g2_decap_8 FILLER_155_500 ();
 sg13g2_decap_4 FILLER_155_527 ();
 sg13g2_fill_1 FILLER_155_531 ();
 sg13g2_fill_2 FILLER_155_540 ();
 sg13g2_fill_2 FILLER_155_550 ();
 sg13g2_decap_8 FILLER_155_560 ();
 sg13g2_decap_8 FILLER_155_567 ();
 sg13g2_decap_8 FILLER_155_574 ();
 sg13g2_decap_4 FILLER_155_581 ();
 sg13g2_fill_1 FILLER_155_585 ();
 sg13g2_decap_8 FILLER_155_590 ();
 sg13g2_decap_8 FILLER_155_597 ();
 sg13g2_decap_8 FILLER_155_604 ();
 sg13g2_decap_8 FILLER_155_629 ();
 sg13g2_decap_8 FILLER_155_636 ();
 sg13g2_decap_8 FILLER_155_643 ();
 sg13g2_decap_8 FILLER_155_650 ();
 sg13g2_decap_8 FILLER_155_657 ();
 sg13g2_decap_8 FILLER_155_664 ();
 sg13g2_fill_1 FILLER_155_671 ();
 sg13g2_decap_8 FILLER_155_685 ();
 sg13g2_decap_8 FILLER_155_692 ();
 sg13g2_decap_8 FILLER_155_699 ();
 sg13g2_decap_8 FILLER_155_706 ();
 sg13g2_decap_8 FILLER_155_713 ();
 sg13g2_fill_1 FILLER_155_720 ();
 sg13g2_fill_2 FILLER_155_729 ();
 sg13g2_fill_1 FILLER_155_731 ();
 sg13g2_decap_8 FILLER_155_740 ();
 sg13g2_fill_2 FILLER_155_747 ();
 sg13g2_fill_1 FILLER_155_749 ();
 sg13g2_decap_8 FILLER_155_772 ();
 sg13g2_fill_2 FILLER_155_779 ();
 sg13g2_fill_1 FILLER_155_781 ();
 sg13g2_decap_8 FILLER_155_803 ();
 sg13g2_decap_8 FILLER_155_810 ();
 sg13g2_decap_8 FILLER_155_817 ();
 sg13g2_decap_8 FILLER_155_824 ();
 sg13g2_decap_8 FILLER_155_831 ();
 sg13g2_decap_8 FILLER_155_838 ();
 sg13g2_decap_4 FILLER_155_845 ();
 sg13g2_fill_2 FILLER_155_849 ();
 sg13g2_decap_8 FILLER_155_856 ();
 sg13g2_decap_8 FILLER_155_863 ();
 sg13g2_decap_8 FILLER_155_870 ();
 sg13g2_decap_8 FILLER_155_877 ();
 sg13g2_decap_8 FILLER_155_884 ();
 sg13g2_decap_8 FILLER_155_891 ();
 sg13g2_decap_8 FILLER_155_898 ();
 sg13g2_decap_8 FILLER_155_905 ();
 sg13g2_decap_8 FILLER_155_912 ();
 sg13g2_decap_8 FILLER_155_919 ();
 sg13g2_fill_2 FILLER_155_926 ();
 sg13g2_decap_4 FILLER_155_932 ();
 sg13g2_fill_1 FILLER_155_936 ();
 sg13g2_decap_8 FILLER_155_942 ();
 sg13g2_decap_8 FILLER_155_949 ();
 sg13g2_decap_8 FILLER_155_956 ();
 sg13g2_decap_8 FILLER_155_963 ();
 sg13g2_decap_4 FILLER_155_970 ();
 sg13g2_decap_8 FILLER_155_986 ();
 sg13g2_decap_8 FILLER_155_1005 ();
 sg13g2_decap_8 FILLER_155_1012 ();
 sg13g2_decap_4 FILLER_155_1019 ();
 sg13g2_fill_2 FILLER_155_1023 ();
 sg13g2_decap_8 FILLER_155_1057 ();
 sg13g2_decap_8 FILLER_155_1064 ();
 sg13g2_decap_8 FILLER_155_1071 ();
 sg13g2_decap_8 FILLER_155_1078 ();
 sg13g2_decap_8 FILLER_155_1085 ();
 sg13g2_fill_2 FILLER_155_1092 ();
 sg13g2_decap_8 FILLER_155_1104 ();
 sg13g2_decap_8 FILLER_155_1111 ();
 sg13g2_decap_8 FILLER_155_1118 ();
 sg13g2_decap_8 FILLER_155_1125 ();
 sg13g2_decap_8 FILLER_155_1132 ();
 sg13g2_decap_8 FILLER_155_1139 ();
 sg13g2_decap_8 FILLER_155_1146 ();
 sg13g2_decap_4 FILLER_155_1153 ();
 sg13g2_fill_2 FILLER_155_1157 ();
 sg13g2_fill_1 FILLER_155_1167 ();
 sg13g2_decap_8 FILLER_155_1173 ();
 sg13g2_decap_8 FILLER_155_1180 ();
 sg13g2_decap_8 FILLER_155_1187 ();
 sg13g2_fill_2 FILLER_155_1194 ();
 sg13g2_fill_1 FILLER_155_1196 ();
 sg13g2_decap_4 FILLER_155_1213 ();
 sg13g2_fill_1 FILLER_155_1217 ();
 sg13g2_fill_2 FILLER_155_1226 ();
 sg13g2_fill_1 FILLER_155_1228 ();
 sg13g2_fill_2 FILLER_155_1258 ();
 sg13g2_fill_1 FILLER_155_1260 ();
 sg13g2_decap_8 FILLER_155_1265 ();
 sg13g2_decap_8 FILLER_155_1272 ();
 sg13g2_decap_8 FILLER_155_1279 ();
 sg13g2_decap_8 FILLER_155_1286 ();
 sg13g2_decap_8 FILLER_155_1299 ();
 sg13g2_decap_4 FILLER_155_1306 ();
 sg13g2_fill_2 FILLER_155_1310 ();
 sg13g2_decap_8 FILLER_155_1336 ();
 sg13g2_decap_8 FILLER_155_1343 ();
 sg13g2_decap_8 FILLER_155_1350 ();
 sg13g2_decap_8 FILLER_155_1357 ();
 sg13g2_decap_8 FILLER_155_1364 ();
 sg13g2_decap_8 FILLER_155_1371 ();
 sg13g2_decap_8 FILLER_155_1378 ();
 sg13g2_decap_8 FILLER_155_1385 ();
 sg13g2_decap_4 FILLER_155_1392 ();
 sg13g2_decap_4 FILLER_155_1404 ();
 sg13g2_fill_1 FILLER_155_1408 ();
 sg13g2_fill_2 FILLER_155_1422 ();
 sg13g2_decap_8 FILLER_155_1432 ();
 sg13g2_decap_8 FILLER_155_1439 ();
 sg13g2_decap_8 FILLER_155_1446 ();
 sg13g2_decap_8 FILLER_155_1453 ();
 sg13g2_decap_4 FILLER_155_1460 ();
 sg13g2_fill_2 FILLER_155_1464 ();
 sg13g2_decap_8 FILLER_155_1483 ();
 sg13g2_decap_8 FILLER_155_1490 ();
 sg13g2_decap_8 FILLER_155_1497 ();
 sg13g2_decap_8 FILLER_155_1504 ();
 sg13g2_decap_4 FILLER_155_1511 ();
 sg13g2_fill_2 FILLER_155_1515 ();
 sg13g2_decap_8 FILLER_155_1522 ();
 sg13g2_decap_8 FILLER_155_1529 ();
 sg13g2_decap_8 FILLER_155_1536 ();
 sg13g2_decap_8 FILLER_155_1543 ();
 sg13g2_decap_8 FILLER_155_1550 ();
 sg13g2_decap_8 FILLER_155_1557 ();
 sg13g2_decap_8 FILLER_155_1564 ();
 sg13g2_fill_1 FILLER_155_1571 ();
 sg13g2_decap_8 FILLER_155_1596 ();
 sg13g2_decap_8 FILLER_155_1603 ();
 sg13g2_decap_8 FILLER_155_1610 ();
 sg13g2_decap_8 FILLER_155_1617 ();
 sg13g2_decap_8 FILLER_155_1624 ();
 sg13g2_decap_8 FILLER_155_1631 ();
 sg13g2_decap_8 FILLER_155_1638 ();
 sg13g2_decap_8 FILLER_155_1645 ();
 sg13g2_decap_8 FILLER_155_1652 ();
 sg13g2_decap_8 FILLER_155_1659 ();
 sg13g2_decap_8 FILLER_155_1666 ();
 sg13g2_decap_8 FILLER_155_1673 ();
 sg13g2_decap_8 FILLER_155_1680 ();
 sg13g2_decap_8 FILLER_155_1687 ();
 sg13g2_decap_8 FILLER_155_1694 ();
 sg13g2_decap_8 FILLER_155_1701 ();
 sg13g2_decap_8 FILLER_155_1708 ();
 sg13g2_decap_8 FILLER_155_1715 ();
 sg13g2_decap_8 FILLER_155_1722 ();
 sg13g2_decap_8 FILLER_155_1729 ();
 sg13g2_decap_8 FILLER_155_1736 ();
 sg13g2_decap_8 FILLER_155_1743 ();
 sg13g2_decap_8 FILLER_155_1750 ();
 sg13g2_decap_8 FILLER_155_1757 ();
 sg13g2_decap_4 FILLER_155_1764 ();
 sg13g2_decap_8 FILLER_156_0 ();
 sg13g2_decap_8 FILLER_156_7 ();
 sg13g2_decap_4 FILLER_156_14 ();
 sg13g2_fill_1 FILLER_156_18 ();
 sg13g2_decap_8 FILLER_156_50 ();
 sg13g2_decap_8 FILLER_156_57 ();
 sg13g2_decap_8 FILLER_156_64 ();
 sg13g2_decap_8 FILLER_156_71 ();
 sg13g2_decap_4 FILLER_156_78 ();
 sg13g2_fill_2 FILLER_156_82 ();
 sg13g2_decap_8 FILLER_156_92 ();
 sg13g2_decap_4 FILLER_156_99 ();
 sg13g2_fill_1 FILLER_156_103 ();
 sg13g2_decap_8 FILLER_156_127 ();
 sg13g2_decap_8 FILLER_156_134 ();
 sg13g2_decap_8 FILLER_156_141 ();
 sg13g2_decap_8 FILLER_156_148 ();
 sg13g2_decap_8 FILLER_156_155 ();
 sg13g2_decap_8 FILLER_156_162 ();
 sg13g2_decap_8 FILLER_156_169 ();
 sg13g2_decap_8 FILLER_156_176 ();
 sg13g2_decap_8 FILLER_156_183 ();
 sg13g2_decap_8 FILLER_156_190 ();
 sg13g2_decap_8 FILLER_156_197 ();
 sg13g2_decap_8 FILLER_156_204 ();
 sg13g2_decap_4 FILLER_156_211 ();
 sg13g2_fill_1 FILLER_156_215 ();
 sg13g2_fill_2 FILLER_156_220 ();
 sg13g2_fill_1 FILLER_156_222 ();
 sg13g2_decap_8 FILLER_156_237 ();
 sg13g2_decap_8 FILLER_156_244 ();
 sg13g2_decap_8 FILLER_156_251 ();
 sg13g2_decap_8 FILLER_156_258 ();
 sg13g2_decap_8 FILLER_156_265 ();
 sg13g2_decap_8 FILLER_156_272 ();
 sg13g2_decap_8 FILLER_156_279 ();
 sg13g2_decap_8 FILLER_156_286 ();
 sg13g2_decap_8 FILLER_156_293 ();
 sg13g2_decap_8 FILLER_156_300 ();
 sg13g2_decap_8 FILLER_156_307 ();
 sg13g2_decap_8 FILLER_156_314 ();
 sg13g2_decap_8 FILLER_156_321 ();
 sg13g2_decap_8 FILLER_156_328 ();
 sg13g2_decap_8 FILLER_156_335 ();
 sg13g2_decap_8 FILLER_156_342 ();
 sg13g2_decap_8 FILLER_156_349 ();
 sg13g2_decap_8 FILLER_156_356 ();
 sg13g2_decap_8 FILLER_156_363 ();
 sg13g2_decap_4 FILLER_156_370 ();
 sg13g2_fill_1 FILLER_156_374 ();
 sg13g2_decap_8 FILLER_156_388 ();
 sg13g2_decap_8 FILLER_156_412 ();
 sg13g2_decap_8 FILLER_156_419 ();
 sg13g2_decap_8 FILLER_156_426 ();
 sg13g2_decap_8 FILLER_156_433 ();
 sg13g2_decap_8 FILLER_156_440 ();
 sg13g2_decap_8 FILLER_156_447 ();
 sg13g2_decap_8 FILLER_156_454 ();
 sg13g2_fill_2 FILLER_156_461 ();
 sg13g2_decap_8 FILLER_156_471 ();
 sg13g2_decap_8 FILLER_156_478 ();
 sg13g2_decap_8 FILLER_156_485 ();
 sg13g2_decap_8 FILLER_156_492 ();
 sg13g2_decap_8 FILLER_156_499 ();
 sg13g2_decap_8 FILLER_156_506 ();
 sg13g2_decap_8 FILLER_156_513 ();
 sg13g2_decap_8 FILLER_156_520 ();
 sg13g2_decap_8 FILLER_156_527 ();
 sg13g2_decap_8 FILLER_156_534 ();
 sg13g2_decap_8 FILLER_156_541 ();
 sg13g2_decap_8 FILLER_156_548 ();
 sg13g2_decap_8 FILLER_156_555 ();
 sg13g2_decap_8 FILLER_156_562 ();
 sg13g2_decap_8 FILLER_156_569 ();
 sg13g2_fill_2 FILLER_156_576 ();
 sg13g2_fill_1 FILLER_156_578 ();
 sg13g2_decap_4 FILLER_156_600 ();
 sg13g2_fill_2 FILLER_156_604 ();
 sg13g2_decap_8 FILLER_156_622 ();
 sg13g2_decap_8 FILLER_156_629 ();
 sg13g2_decap_8 FILLER_156_636 ();
 sg13g2_decap_8 FILLER_156_643 ();
 sg13g2_decap_8 FILLER_156_650 ();
 sg13g2_decap_8 FILLER_156_657 ();
 sg13g2_decap_8 FILLER_156_664 ();
 sg13g2_decap_8 FILLER_156_671 ();
 sg13g2_decap_8 FILLER_156_678 ();
 sg13g2_decap_8 FILLER_156_685 ();
 sg13g2_decap_4 FILLER_156_692 ();
 sg13g2_fill_1 FILLER_156_696 ();
 sg13g2_decap_8 FILLER_156_709 ();
 sg13g2_decap_4 FILLER_156_720 ();
 sg13g2_fill_1 FILLER_156_724 ();
 sg13g2_decap_8 FILLER_156_737 ();
 sg13g2_decap_8 FILLER_156_744 ();
 sg13g2_decap_4 FILLER_156_751 ();
 sg13g2_fill_1 FILLER_156_755 ();
 sg13g2_decap_8 FILLER_156_760 ();
 sg13g2_decap_4 FILLER_156_767 ();
 sg13g2_fill_2 FILLER_156_771 ();
 sg13g2_decap_8 FILLER_156_777 ();
 sg13g2_fill_1 FILLER_156_784 ();
 sg13g2_decap_8 FILLER_156_809 ();
 sg13g2_decap_8 FILLER_156_816 ();
 sg13g2_decap_8 FILLER_156_823 ();
 sg13g2_decap_8 FILLER_156_830 ();
 sg13g2_decap_8 FILLER_156_837 ();
 sg13g2_decap_8 FILLER_156_844 ();
 sg13g2_decap_8 FILLER_156_851 ();
 sg13g2_decap_8 FILLER_156_858 ();
 sg13g2_decap_8 FILLER_156_865 ();
 sg13g2_decap_4 FILLER_156_872 ();
 sg13g2_fill_2 FILLER_156_876 ();
 sg13g2_decap_8 FILLER_156_895 ();
 sg13g2_decap_8 FILLER_156_902 ();
 sg13g2_decap_8 FILLER_156_909 ();
 sg13g2_decap_4 FILLER_156_916 ();
 sg13g2_fill_2 FILLER_156_920 ();
 sg13g2_decap_8 FILLER_156_939 ();
 sg13g2_decap_4 FILLER_156_946 ();
 sg13g2_decap_8 FILLER_156_958 ();
 sg13g2_decap_8 FILLER_156_965 ();
 sg13g2_decap_8 FILLER_156_972 ();
 sg13g2_decap_8 FILLER_156_979 ();
 sg13g2_decap_8 FILLER_156_986 ();
 sg13g2_decap_8 FILLER_156_993 ();
 sg13g2_decap_8 FILLER_156_1000 ();
 sg13g2_decap_8 FILLER_156_1007 ();
 sg13g2_decap_8 FILLER_156_1014 ();
 sg13g2_decap_8 FILLER_156_1021 ();
 sg13g2_fill_2 FILLER_156_1028 ();
 sg13g2_decap_8 FILLER_156_1059 ();
 sg13g2_decap_8 FILLER_156_1066 ();
 sg13g2_decap_8 FILLER_156_1073 ();
 sg13g2_decap_8 FILLER_156_1080 ();
 sg13g2_fill_2 FILLER_156_1087 ();
 sg13g2_fill_1 FILLER_156_1089 ();
 sg13g2_decap_4 FILLER_156_1103 ();
 sg13g2_fill_1 FILLER_156_1107 ();
 sg13g2_decap_8 FILLER_156_1116 ();
 sg13g2_decap_8 FILLER_156_1123 ();
 sg13g2_decap_8 FILLER_156_1130 ();
 sg13g2_decap_8 FILLER_156_1137 ();
 sg13g2_decap_8 FILLER_156_1144 ();
 sg13g2_decap_8 FILLER_156_1151 ();
 sg13g2_decap_4 FILLER_156_1158 ();
 sg13g2_fill_2 FILLER_156_1162 ();
 sg13g2_decap_8 FILLER_156_1180 ();
 sg13g2_fill_2 FILLER_156_1187 ();
 sg13g2_decap_8 FILLER_156_1194 ();
 sg13g2_decap_8 FILLER_156_1201 ();
 sg13g2_decap_8 FILLER_156_1208 ();
 sg13g2_decap_8 FILLER_156_1219 ();
 sg13g2_decap_8 FILLER_156_1226 ();
 sg13g2_decap_8 FILLER_156_1233 ();
 sg13g2_decap_8 FILLER_156_1240 ();
 sg13g2_decap_8 FILLER_156_1247 ();
 sg13g2_fill_2 FILLER_156_1254 ();
 sg13g2_fill_1 FILLER_156_1256 ();
 sg13g2_decap_8 FILLER_156_1286 ();
 sg13g2_decap_8 FILLER_156_1293 ();
 sg13g2_decap_8 FILLER_156_1300 ();
 sg13g2_decap_8 FILLER_156_1307 ();
 sg13g2_decap_8 FILLER_156_1314 ();
 sg13g2_fill_2 FILLER_156_1321 ();
 sg13g2_decap_8 FILLER_156_1331 ();
 sg13g2_decap_4 FILLER_156_1338 ();
 sg13g2_decap_8 FILLER_156_1346 ();
 sg13g2_decap_8 FILLER_156_1353 ();
 sg13g2_decap_8 FILLER_156_1360 ();
 sg13g2_decap_8 FILLER_156_1367 ();
 sg13g2_decap_8 FILLER_156_1374 ();
 sg13g2_decap_8 FILLER_156_1381 ();
 sg13g2_decap_8 FILLER_156_1388 ();
 sg13g2_fill_2 FILLER_156_1395 ();
 sg13g2_fill_2 FILLER_156_1405 ();
 sg13g2_fill_1 FILLER_156_1414 ();
 sg13g2_decap_8 FILLER_156_1420 ();
 sg13g2_fill_2 FILLER_156_1427 ();
 sg13g2_decap_8 FILLER_156_1433 ();
 sg13g2_decap_8 FILLER_156_1440 ();
 sg13g2_decap_8 FILLER_156_1447 ();
 sg13g2_decap_8 FILLER_156_1454 ();
 sg13g2_decap_8 FILLER_156_1461 ();
 sg13g2_fill_1 FILLER_156_1468 ();
 sg13g2_decap_8 FILLER_156_1490 ();
 sg13g2_decap_8 FILLER_156_1497 ();
 sg13g2_decap_8 FILLER_156_1504 ();
 sg13g2_fill_2 FILLER_156_1511 ();
 sg13g2_fill_1 FILLER_156_1513 ();
 sg13g2_decap_8 FILLER_156_1527 ();
 sg13g2_decap_8 FILLER_156_1534 ();
 sg13g2_decap_8 FILLER_156_1549 ();
 sg13g2_decap_8 FILLER_156_1556 ();
 sg13g2_decap_4 FILLER_156_1563 ();
 sg13g2_fill_2 FILLER_156_1576 ();
 sg13g2_decap_8 FILLER_156_1583 ();
 sg13g2_decap_8 FILLER_156_1590 ();
 sg13g2_decap_8 FILLER_156_1597 ();
 sg13g2_decap_8 FILLER_156_1604 ();
 sg13g2_decap_8 FILLER_156_1611 ();
 sg13g2_decap_8 FILLER_156_1618 ();
 sg13g2_decap_8 FILLER_156_1625 ();
 sg13g2_decap_8 FILLER_156_1632 ();
 sg13g2_decap_8 FILLER_156_1639 ();
 sg13g2_decap_8 FILLER_156_1646 ();
 sg13g2_decap_8 FILLER_156_1653 ();
 sg13g2_decap_8 FILLER_156_1660 ();
 sg13g2_decap_8 FILLER_156_1667 ();
 sg13g2_decap_8 FILLER_156_1674 ();
 sg13g2_decap_8 FILLER_156_1681 ();
 sg13g2_decap_8 FILLER_156_1688 ();
 sg13g2_decap_8 FILLER_156_1695 ();
 sg13g2_decap_8 FILLER_156_1702 ();
 sg13g2_decap_8 FILLER_156_1709 ();
 sg13g2_decap_8 FILLER_156_1716 ();
 sg13g2_decap_8 FILLER_156_1723 ();
 sg13g2_decap_8 FILLER_156_1730 ();
 sg13g2_decap_8 FILLER_156_1737 ();
 sg13g2_decap_8 FILLER_156_1744 ();
 sg13g2_decap_8 FILLER_156_1751 ();
 sg13g2_decap_8 FILLER_156_1758 ();
 sg13g2_fill_2 FILLER_156_1765 ();
 sg13g2_fill_1 FILLER_156_1767 ();
 sg13g2_decap_8 FILLER_157_0 ();
 sg13g2_decap_8 FILLER_157_7 ();
 sg13g2_decap_8 FILLER_157_14 ();
 sg13g2_decap_8 FILLER_157_21 ();
 sg13g2_fill_2 FILLER_157_28 ();
 sg13g2_fill_1 FILLER_157_30 ();
 sg13g2_decap_8 FILLER_157_53 ();
 sg13g2_decap_8 FILLER_157_60 ();
 sg13g2_decap_8 FILLER_157_67 ();
 sg13g2_decap_8 FILLER_157_74 ();
 sg13g2_decap_8 FILLER_157_81 ();
 sg13g2_decap_8 FILLER_157_88 ();
 sg13g2_decap_8 FILLER_157_95 ();
 sg13g2_decap_8 FILLER_157_102 ();
 sg13g2_decap_8 FILLER_157_109 ();
 sg13g2_decap_8 FILLER_157_116 ();
 sg13g2_decap_8 FILLER_157_123 ();
 sg13g2_decap_8 FILLER_157_130 ();
 sg13g2_decap_8 FILLER_157_137 ();
 sg13g2_decap_8 FILLER_157_144 ();
 sg13g2_decap_8 FILLER_157_151 ();
 sg13g2_decap_8 FILLER_157_158 ();
 sg13g2_decap_8 FILLER_157_165 ();
 sg13g2_decap_4 FILLER_157_172 ();
 sg13g2_fill_1 FILLER_157_176 ();
 sg13g2_decap_4 FILLER_157_202 ();
 sg13g2_fill_1 FILLER_157_206 ();
 sg13g2_fill_1 FILLER_157_232 ();
 sg13g2_decap_8 FILLER_157_238 ();
 sg13g2_decap_4 FILLER_157_245 ();
 sg13g2_decap_8 FILLER_157_254 ();
 sg13g2_fill_1 FILLER_157_261 ();
 sg13g2_decap_8 FILLER_157_272 ();
 sg13g2_fill_2 FILLER_157_279 ();
 sg13g2_decap_4 FILLER_157_307 ();
 sg13g2_fill_2 FILLER_157_311 ();
 sg13g2_fill_2 FILLER_157_318 ();
 sg13g2_decap_8 FILLER_157_330 ();
 sg13g2_decap_4 FILLER_157_337 ();
 sg13g2_decap_8 FILLER_157_345 ();
 sg13g2_decap_8 FILLER_157_352 ();
 sg13g2_decap_4 FILLER_157_359 ();
 sg13g2_fill_1 FILLER_157_363 ();
 sg13g2_decap_8 FILLER_157_377 ();
 sg13g2_decap_8 FILLER_157_384 ();
 sg13g2_fill_2 FILLER_157_391 ();
 sg13g2_decap_8 FILLER_157_423 ();
 sg13g2_decap_8 FILLER_157_430 ();
 sg13g2_decap_8 FILLER_157_437 ();
 sg13g2_decap_8 FILLER_157_444 ();
 sg13g2_decap_8 FILLER_157_451 ();
 sg13g2_fill_2 FILLER_157_458 ();
 sg13g2_fill_2 FILLER_157_467 ();
 sg13g2_decap_8 FILLER_157_485 ();
 sg13g2_decap_8 FILLER_157_492 ();
 sg13g2_decap_8 FILLER_157_499 ();
 sg13g2_decap_8 FILLER_157_506 ();
 sg13g2_fill_2 FILLER_157_513 ();
 sg13g2_decap_8 FILLER_157_519 ();
 sg13g2_decap_8 FILLER_157_526 ();
 sg13g2_decap_8 FILLER_157_533 ();
 sg13g2_decap_8 FILLER_157_540 ();
 sg13g2_decap_4 FILLER_157_547 ();
 sg13g2_fill_1 FILLER_157_551 ();
 sg13g2_decap_8 FILLER_157_556 ();
 sg13g2_decap_8 FILLER_157_563 ();
 sg13g2_decap_4 FILLER_157_570 ();
 sg13g2_fill_2 FILLER_157_574 ();
 sg13g2_decap_8 FILLER_157_592 ();
 sg13g2_decap_8 FILLER_157_599 ();
 sg13g2_decap_8 FILLER_157_606 ();
 sg13g2_decap_8 FILLER_157_613 ();
 sg13g2_decap_8 FILLER_157_620 ();
 sg13g2_decap_8 FILLER_157_627 ();
 sg13g2_decap_4 FILLER_157_634 ();
 sg13g2_fill_2 FILLER_157_638 ();
 sg13g2_decap_8 FILLER_157_657 ();
 sg13g2_decap_8 FILLER_157_664 ();
 sg13g2_decap_8 FILLER_157_671 ();
 sg13g2_decap_8 FILLER_157_678 ();
 sg13g2_decap_8 FILLER_157_685 ();
 sg13g2_decap_8 FILLER_157_692 ();
 sg13g2_decap_8 FILLER_157_699 ();
 sg13g2_decap_8 FILLER_157_706 ();
 sg13g2_fill_2 FILLER_157_713 ();
 sg13g2_decap_8 FILLER_157_733 ();
 sg13g2_decap_8 FILLER_157_740 ();
 sg13g2_decap_8 FILLER_157_747 ();
 sg13g2_decap_8 FILLER_157_754 ();
 sg13g2_decap_4 FILLER_157_761 ();
 sg13g2_decap_8 FILLER_157_774 ();
 sg13g2_fill_2 FILLER_157_781 ();
 sg13g2_decap_8 FILLER_157_799 ();
 sg13g2_decap_8 FILLER_157_806 ();
 sg13g2_decap_8 FILLER_157_813 ();
 sg13g2_decap_8 FILLER_157_820 ();
 sg13g2_decap_8 FILLER_157_827 ();
 sg13g2_decap_8 FILLER_157_834 ();
 sg13g2_decap_8 FILLER_157_850 ();
 sg13g2_decap_8 FILLER_157_857 ();
 sg13g2_decap_4 FILLER_157_864 ();
 sg13g2_fill_1 FILLER_157_868 ();
 sg13g2_fill_2 FILLER_157_878 ();
 sg13g2_decap_8 FILLER_157_892 ();
 sg13g2_decap_8 FILLER_157_899 ();
 sg13g2_decap_4 FILLER_157_906 ();
 sg13g2_fill_1 FILLER_157_910 ();
 sg13g2_decap_8 FILLER_157_919 ();
 sg13g2_decap_8 FILLER_157_934 ();
 sg13g2_decap_8 FILLER_157_941 ();
 sg13g2_fill_2 FILLER_157_948 ();
 sg13g2_fill_1 FILLER_157_950 ();
 sg13g2_decap_8 FILLER_157_955 ();
 sg13g2_decap_8 FILLER_157_962 ();
 sg13g2_decap_8 FILLER_157_969 ();
 sg13g2_decap_8 FILLER_157_976 ();
 sg13g2_decap_4 FILLER_157_983 ();
 sg13g2_fill_2 FILLER_157_987 ();
 sg13g2_decap_8 FILLER_157_997 ();
 sg13g2_decap_8 FILLER_157_1004 ();
 sg13g2_decap_8 FILLER_157_1011 ();
 sg13g2_decap_8 FILLER_157_1018 ();
 sg13g2_decap_8 FILLER_157_1025 ();
 sg13g2_fill_2 FILLER_157_1032 ();
 sg13g2_fill_1 FILLER_157_1034 ();
 sg13g2_fill_2 FILLER_157_1040 ();
 sg13g2_decap_8 FILLER_157_1050 ();
 sg13g2_decap_8 FILLER_157_1057 ();
 sg13g2_decap_8 FILLER_157_1064 ();
 sg13g2_decap_8 FILLER_157_1071 ();
 sg13g2_fill_2 FILLER_157_1078 ();
 sg13g2_fill_1 FILLER_157_1080 ();
 sg13g2_decap_8 FILLER_157_1094 ();
 sg13g2_decap_8 FILLER_157_1101 ();
 sg13g2_fill_2 FILLER_157_1108 ();
 sg13g2_decap_8 FILLER_157_1128 ();
 sg13g2_decap_8 FILLER_157_1135 ();
 sg13g2_decap_8 FILLER_157_1142 ();
 sg13g2_decap_8 FILLER_157_1149 ();
 sg13g2_decap_4 FILLER_157_1156 ();
 sg13g2_fill_2 FILLER_157_1160 ();
 sg13g2_decap_8 FILLER_157_1178 ();
 sg13g2_decap_4 FILLER_157_1185 ();
 sg13g2_decap_8 FILLER_157_1193 ();
 sg13g2_decap_8 FILLER_157_1204 ();
 sg13g2_fill_2 FILLER_157_1211 ();
 sg13g2_fill_1 FILLER_157_1213 ();
 sg13g2_decap_8 FILLER_157_1222 ();
 sg13g2_decap_8 FILLER_157_1229 ();
 sg13g2_decap_8 FILLER_157_1236 ();
 sg13g2_decap_8 FILLER_157_1243 ();
 sg13g2_decap_4 FILLER_157_1250 ();
 sg13g2_fill_2 FILLER_157_1254 ();
 sg13g2_decap_4 FILLER_157_1272 ();
 sg13g2_decap_8 FILLER_157_1284 ();
 sg13g2_decap_8 FILLER_157_1291 ();
 sg13g2_decap_8 FILLER_157_1298 ();
 sg13g2_decap_8 FILLER_157_1305 ();
 sg13g2_decap_8 FILLER_157_1312 ();
 sg13g2_decap_8 FILLER_157_1319 ();
 sg13g2_decap_4 FILLER_157_1326 ();
 sg13g2_fill_2 FILLER_157_1330 ();
 sg13g2_decap_8 FILLER_157_1357 ();
 sg13g2_decap_8 FILLER_157_1364 ();
 sg13g2_decap_8 FILLER_157_1371 ();
 sg13g2_decap_8 FILLER_157_1378 ();
 sg13g2_decap_8 FILLER_157_1385 ();
 sg13g2_decap_8 FILLER_157_1392 ();
 sg13g2_decap_8 FILLER_157_1399 ();
 sg13g2_decap_8 FILLER_157_1406 ();
 sg13g2_fill_2 FILLER_157_1413 ();
 sg13g2_fill_1 FILLER_157_1415 ();
 sg13g2_decap_8 FILLER_157_1435 ();
 sg13g2_decap_8 FILLER_157_1442 ();
 sg13g2_decap_8 FILLER_157_1449 ();
 sg13g2_decap_8 FILLER_157_1456 ();
 sg13g2_decap_4 FILLER_157_1463 ();
 sg13g2_fill_1 FILLER_157_1467 ();
 sg13g2_decap_8 FILLER_157_1488 ();
 sg13g2_decap_8 FILLER_157_1495 ();
 sg13g2_decap_4 FILLER_157_1502 ();
 sg13g2_decap_8 FILLER_157_1519 ();
 sg13g2_decap_4 FILLER_157_1526 ();
 sg13g2_fill_1 FILLER_157_1530 ();
 sg13g2_fill_2 FILLER_157_1543 ();
 sg13g2_fill_1 FILLER_157_1545 ();
 sg13g2_decap_8 FILLER_157_1554 ();
 sg13g2_decap_8 FILLER_157_1561 ();
 sg13g2_decap_8 FILLER_157_1568 ();
 sg13g2_decap_8 FILLER_157_1575 ();
 sg13g2_decap_8 FILLER_157_1582 ();
 sg13g2_decap_8 FILLER_157_1589 ();
 sg13g2_decap_8 FILLER_157_1596 ();
 sg13g2_decap_8 FILLER_157_1603 ();
 sg13g2_decap_8 FILLER_157_1610 ();
 sg13g2_decap_8 FILLER_157_1617 ();
 sg13g2_decap_8 FILLER_157_1624 ();
 sg13g2_decap_8 FILLER_157_1631 ();
 sg13g2_decap_8 FILLER_157_1638 ();
 sg13g2_decap_8 FILLER_157_1645 ();
 sg13g2_decap_8 FILLER_157_1652 ();
 sg13g2_decap_8 FILLER_157_1659 ();
 sg13g2_decap_8 FILLER_157_1666 ();
 sg13g2_decap_8 FILLER_157_1673 ();
 sg13g2_decap_8 FILLER_157_1680 ();
 sg13g2_decap_8 FILLER_157_1687 ();
 sg13g2_decap_8 FILLER_157_1694 ();
 sg13g2_decap_8 FILLER_157_1701 ();
 sg13g2_decap_8 FILLER_157_1708 ();
 sg13g2_decap_8 FILLER_157_1715 ();
 sg13g2_decap_8 FILLER_157_1722 ();
 sg13g2_decap_8 FILLER_157_1729 ();
 sg13g2_decap_8 FILLER_157_1736 ();
 sg13g2_decap_8 FILLER_157_1743 ();
 sg13g2_decap_8 FILLER_157_1750 ();
 sg13g2_decap_8 FILLER_157_1757 ();
 sg13g2_decap_4 FILLER_157_1764 ();
 sg13g2_decap_8 FILLER_158_0 ();
 sg13g2_decap_8 FILLER_158_7 ();
 sg13g2_decap_8 FILLER_158_14 ();
 sg13g2_decap_8 FILLER_158_21 ();
 sg13g2_decap_8 FILLER_158_28 ();
 sg13g2_fill_1 FILLER_158_35 ();
 sg13g2_decap_8 FILLER_158_56 ();
 sg13g2_decap_8 FILLER_158_63 ();
 sg13g2_decap_8 FILLER_158_70 ();
 sg13g2_decap_8 FILLER_158_77 ();
 sg13g2_decap_8 FILLER_158_84 ();
 sg13g2_decap_8 FILLER_158_91 ();
 sg13g2_fill_1 FILLER_158_103 ();
 sg13g2_decap_8 FILLER_158_115 ();
 sg13g2_decap_8 FILLER_158_122 ();
 sg13g2_decap_8 FILLER_158_129 ();
 sg13g2_decap_8 FILLER_158_136 ();
 sg13g2_decap_8 FILLER_158_143 ();
 sg13g2_decap_8 FILLER_158_150 ();
 sg13g2_fill_2 FILLER_158_157 ();
 sg13g2_fill_1 FILLER_158_159 ();
 sg13g2_decap_8 FILLER_158_196 ();
 sg13g2_decap_8 FILLER_158_203 ();
 sg13g2_decap_8 FILLER_158_210 ();
 sg13g2_decap_8 FILLER_158_217 ();
 sg13g2_fill_2 FILLER_158_224 ();
 sg13g2_fill_2 FILLER_158_234 ();
 sg13g2_fill_1 FILLER_158_236 ();
 sg13g2_fill_1 FILLER_158_289 ();
 sg13g2_decap_8 FILLER_158_299 ();
 sg13g2_decap_8 FILLER_158_306 ();
 sg13g2_decap_8 FILLER_158_313 ();
 sg13g2_decap_8 FILLER_158_320 ();
 sg13g2_fill_2 FILLER_158_327 ();
 sg13g2_fill_1 FILLER_158_329 ();
 sg13g2_decap_8 FILLER_158_356 ();
 sg13g2_decap_8 FILLER_158_363 ();
 sg13g2_decap_8 FILLER_158_370 ();
 sg13g2_decap_8 FILLER_158_377 ();
 sg13g2_decap_8 FILLER_158_384 ();
 sg13g2_decap_8 FILLER_158_391 ();
 sg13g2_fill_1 FILLER_158_398 ();
 sg13g2_decap_8 FILLER_158_415 ();
 sg13g2_fill_2 FILLER_158_422 ();
 sg13g2_decap_8 FILLER_158_432 ();
 sg13g2_decap_8 FILLER_158_439 ();
 sg13g2_decap_4 FILLER_158_446 ();
 sg13g2_decap_8 FILLER_158_460 ();
 sg13g2_decap_8 FILLER_158_467 ();
 sg13g2_decap_8 FILLER_158_474 ();
 sg13g2_decap_4 FILLER_158_481 ();
 sg13g2_fill_2 FILLER_158_485 ();
 sg13g2_decap_8 FILLER_158_491 ();
 sg13g2_fill_2 FILLER_158_498 ();
 sg13g2_fill_1 FILLER_158_500 ();
 sg13g2_fill_1 FILLER_158_509 ();
 sg13g2_decap_4 FILLER_158_527 ();
 sg13g2_fill_2 FILLER_158_539 ();
 sg13g2_decap_8 FILLER_158_558 ();
 sg13g2_decap_8 FILLER_158_565 ();
 sg13g2_decap_8 FILLER_158_572 ();
 sg13g2_decap_4 FILLER_158_579 ();
 sg13g2_fill_2 FILLER_158_583 ();
 sg13g2_decap_8 FILLER_158_588 ();
 sg13g2_decap_8 FILLER_158_595 ();
 sg13g2_decap_8 FILLER_158_602 ();
 sg13g2_decap_4 FILLER_158_609 ();
 sg13g2_fill_1 FILLER_158_613 ();
 sg13g2_decap_8 FILLER_158_622 ();
 sg13g2_decap_8 FILLER_158_629 ();
 sg13g2_fill_1 FILLER_158_636 ();
 sg13g2_decap_4 FILLER_158_641 ();
 sg13g2_decap_8 FILLER_158_653 ();
 sg13g2_decap_8 FILLER_158_660 ();
 sg13g2_decap_8 FILLER_158_667 ();
 sg13g2_decap_8 FILLER_158_674 ();
 sg13g2_decap_8 FILLER_158_681 ();
 sg13g2_decap_8 FILLER_158_688 ();
 sg13g2_decap_8 FILLER_158_695 ();
 sg13g2_decap_4 FILLER_158_702 ();
 sg13g2_fill_2 FILLER_158_706 ();
 sg13g2_fill_1 FILLER_158_716 ();
 sg13g2_fill_1 FILLER_158_725 ();
 sg13g2_decap_8 FILLER_158_734 ();
 sg13g2_decap_8 FILLER_158_741 ();
 sg13g2_decap_8 FILLER_158_748 ();
 sg13g2_decap_4 FILLER_158_755 ();
 sg13g2_fill_2 FILLER_158_759 ();
 sg13g2_decap_8 FILLER_158_764 ();
 sg13g2_decap_8 FILLER_158_771 ();
 sg13g2_fill_2 FILLER_158_778 ();
 sg13g2_fill_2 FILLER_158_792 ();
 sg13g2_fill_1 FILLER_158_794 ();
 sg13g2_decap_8 FILLER_158_803 ();
 sg13g2_decap_8 FILLER_158_810 ();
 sg13g2_decap_8 FILLER_158_817 ();
 sg13g2_decap_8 FILLER_158_824 ();
 sg13g2_decap_8 FILLER_158_831 ();
 sg13g2_decap_8 FILLER_158_838 ();
 sg13g2_decap_8 FILLER_158_845 ();
 sg13g2_decap_4 FILLER_158_852 ();
 sg13g2_fill_1 FILLER_158_856 ();
 sg13g2_fill_2 FILLER_158_881 ();
 sg13g2_fill_1 FILLER_158_883 ();
 sg13g2_decap_8 FILLER_158_896 ();
 sg13g2_fill_1 FILLER_158_903 ();
 sg13g2_decap_8 FILLER_158_912 ();
 sg13g2_decap_8 FILLER_158_919 ();
 sg13g2_decap_8 FILLER_158_926 ();
 sg13g2_decap_8 FILLER_158_933 ();
 sg13g2_decap_8 FILLER_158_940 ();
 sg13g2_decap_4 FILLER_158_947 ();
 sg13g2_fill_2 FILLER_158_951 ();
 sg13g2_fill_1 FILLER_158_961 ();
 sg13g2_decap_8 FILLER_158_970 ();
 sg13g2_fill_2 FILLER_158_977 ();
 sg13g2_fill_1 FILLER_158_979 ();
 sg13g2_decap_8 FILLER_158_986 ();
 sg13g2_decap_8 FILLER_158_1001 ();
 sg13g2_decap_8 FILLER_158_1008 ();
 sg13g2_decap_8 FILLER_158_1015 ();
 sg13g2_decap_8 FILLER_158_1022 ();
 sg13g2_fill_1 FILLER_158_1029 ();
 sg13g2_decap_8 FILLER_158_1046 ();
 sg13g2_decap_8 FILLER_158_1053 ();
 sg13g2_decap_8 FILLER_158_1060 ();
 sg13g2_decap_8 FILLER_158_1088 ();
 sg13g2_decap_8 FILLER_158_1095 ();
 sg13g2_decap_8 FILLER_158_1102 ();
 sg13g2_fill_2 FILLER_158_1109 ();
 sg13g2_decap_8 FILLER_158_1124 ();
 sg13g2_decap_8 FILLER_158_1131 ();
 sg13g2_decap_8 FILLER_158_1138 ();
 sg13g2_decap_8 FILLER_158_1145 ();
 sg13g2_decap_8 FILLER_158_1152 ();
 sg13g2_decap_4 FILLER_158_1159 ();
 sg13g2_fill_1 FILLER_158_1163 ();
 sg13g2_decap_8 FILLER_158_1176 ();
 sg13g2_decap_8 FILLER_158_1183 ();
 sg13g2_decap_4 FILLER_158_1190 ();
 sg13g2_fill_1 FILLER_158_1194 ();
 sg13g2_decap_8 FILLER_158_1219 ();
 sg13g2_decap_8 FILLER_158_1226 ();
 sg13g2_decap_8 FILLER_158_1233 ();
 sg13g2_decap_8 FILLER_158_1240 ();
 sg13g2_decap_8 FILLER_158_1247 ();
 sg13g2_fill_2 FILLER_158_1254 ();
 sg13g2_decap_8 FILLER_158_1264 ();
 sg13g2_decap_8 FILLER_158_1271 ();
 sg13g2_decap_8 FILLER_158_1278 ();
 sg13g2_decap_8 FILLER_158_1285 ();
 sg13g2_decap_8 FILLER_158_1292 ();
 sg13g2_decap_8 FILLER_158_1299 ();
 sg13g2_decap_8 FILLER_158_1306 ();
 sg13g2_decap_8 FILLER_158_1313 ();
 sg13g2_decap_8 FILLER_158_1320 ();
 sg13g2_decap_8 FILLER_158_1327 ();
 sg13g2_decap_8 FILLER_158_1334 ();
 sg13g2_decap_8 FILLER_158_1341 ();
 sg13g2_decap_8 FILLER_158_1348 ();
 sg13g2_fill_2 FILLER_158_1355 ();
 sg13g2_fill_1 FILLER_158_1357 ();
 sg13g2_decap_8 FILLER_158_1375 ();
 sg13g2_decap_8 FILLER_158_1382 ();
 sg13g2_decap_8 FILLER_158_1389 ();
 sg13g2_decap_8 FILLER_158_1396 ();
 sg13g2_decap_8 FILLER_158_1403 ();
 sg13g2_decap_8 FILLER_158_1410 ();
 sg13g2_decap_8 FILLER_158_1417 ();
 sg13g2_decap_8 FILLER_158_1432 ();
 sg13g2_decap_8 FILLER_158_1439 ();
 sg13g2_decap_8 FILLER_158_1446 ();
 sg13g2_decap_8 FILLER_158_1453 ();
 sg13g2_decap_8 FILLER_158_1460 ();
 sg13g2_fill_1 FILLER_158_1467 ();
 sg13g2_decap_8 FILLER_158_1486 ();
 sg13g2_decap_8 FILLER_158_1493 ();
 sg13g2_decap_8 FILLER_158_1500 ();
 sg13g2_decap_8 FILLER_158_1507 ();
 sg13g2_decap_4 FILLER_158_1514 ();
 sg13g2_fill_2 FILLER_158_1538 ();
 sg13g2_decap_8 FILLER_158_1557 ();
 sg13g2_decap_8 FILLER_158_1564 ();
 sg13g2_decap_8 FILLER_158_1571 ();
 sg13g2_decap_8 FILLER_158_1578 ();
 sg13g2_decap_8 FILLER_158_1585 ();
 sg13g2_decap_8 FILLER_158_1592 ();
 sg13g2_decap_8 FILLER_158_1599 ();
 sg13g2_decap_8 FILLER_158_1606 ();
 sg13g2_decap_8 FILLER_158_1613 ();
 sg13g2_decap_8 FILLER_158_1620 ();
 sg13g2_decap_8 FILLER_158_1627 ();
 sg13g2_decap_8 FILLER_158_1634 ();
 sg13g2_decap_8 FILLER_158_1641 ();
 sg13g2_decap_8 FILLER_158_1648 ();
 sg13g2_decap_8 FILLER_158_1655 ();
 sg13g2_decap_8 FILLER_158_1662 ();
 sg13g2_decap_8 FILLER_158_1669 ();
 sg13g2_decap_8 FILLER_158_1676 ();
 sg13g2_decap_8 FILLER_158_1683 ();
 sg13g2_decap_8 FILLER_158_1690 ();
 sg13g2_decap_8 FILLER_158_1697 ();
 sg13g2_decap_8 FILLER_158_1704 ();
 sg13g2_decap_8 FILLER_158_1711 ();
 sg13g2_decap_8 FILLER_158_1718 ();
 sg13g2_decap_8 FILLER_158_1725 ();
 sg13g2_decap_8 FILLER_158_1732 ();
 sg13g2_decap_8 FILLER_158_1739 ();
 sg13g2_decap_8 FILLER_158_1746 ();
 sg13g2_decap_8 FILLER_158_1753 ();
 sg13g2_decap_8 FILLER_158_1760 ();
 sg13g2_fill_1 FILLER_158_1767 ();
 sg13g2_decap_8 FILLER_159_0 ();
 sg13g2_decap_8 FILLER_159_7 ();
 sg13g2_decap_8 FILLER_159_14 ();
 sg13g2_decap_8 FILLER_159_21 ();
 sg13g2_decap_8 FILLER_159_28 ();
 sg13g2_decap_8 FILLER_159_35 ();
 sg13g2_fill_2 FILLER_159_42 ();
 sg13g2_fill_2 FILLER_159_49 ();
 sg13g2_decap_8 FILLER_159_64 ();
 sg13g2_decap_8 FILLER_159_71 ();
 sg13g2_decap_8 FILLER_159_78 ();
 sg13g2_decap_4 FILLER_159_85 ();
 sg13g2_fill_2 FILLER_159_89 ();
 sg13g2_fill_1 FILLER_159_103 ();
 sg13g2_decap_8 FILLER_159_123 ();
 sg13g2_decap_8 FILLER_159_130 ();
 sg13g2_decap_8 FILLER_159_137 ();
 sg13g2_decap_8 FILLER_159_144 ();
 sg13g2_fill_1 FILLER_159_151 ();
 sg13g2_fill_2 FILLER_159_178 ();
 sg13g2_decap_8 FILLER_159_184 ();
 sg13g2_decap_8 FILLER_159_191 ();
 sg13g2_decap_8 FILLER_159_198 ();
 sg13g2_decap_8 FILLER_159_205 ();
 sg13g2_fill_1 FILLER_159_247 ();
 sg13g2_fill_1 FILLER_159_252 ();
 sg13g2_decap_8 FILLER_159_261 ();
 sg13g2_decap_4 FILLER_159_268 ();
 sg13g2_fill_2 FILLER_159_272 ();
 sg13g2_decap_8 FILLER_159_278 ();
 sg13g2_decap_8 FILLER_159_285 ();
 sg13g2_decap_4 FILLER_159_292 ();
 sg13g2_fill_1 FILLER_159_296 ();
 sg13g2_decap_8 FILLER_159_301 ();
 sg13g2_decap_8 FILLER_159_308 ();
 sg13g2_decap_8 FILLER_159_315 ();
 sg13g2_decap_8 FILLER_159_322 ();
 sg13g2_decap_4 FILLER_159_329 ();
 sg13g2_decap_8 FILLER_159_338 ();
 sg13g2_decap_8 FILLER_159_345 ();
 sg13g2_decap_8 FILLER_159_352 ();
 sg13g2_decap_8 FILLER_159_359 ();
 sg13g2_decap_4 FILLER_159_366 ();
 sg13g2_fill_2 FILLER_159_370 ();
 sg13g2_decap_8 FILLER_159_376 ();
 sg13g2_decap_8 FILLER_159_383 ();
 sg13g2_decap_8 FILLER_159_390 ();
 sg13g2_decap_8 FILLER_159_397 ();
 sg13g2_decap_8 FILLER_159_404 ();
 sg13g2_decap_8 FILLER_159_411 ();
 sg13g2_decap_4 FILLER_159_418 ();
 sg13g2_fill_1 FILLER_159_430 ();
 sg13g2_decap_4 FILLER_159_444 ();
 sg13g2_fill_1 FILLER_159_448 ();
 sg13g2_decap_8 FILLER_159_454 ();
 sg13g2_decap_8 FILLER_159_461 ();
 sg13g2_decap_8 FILLER_159_468 ();
 sg13g2_fill_2 FILLER_159_475 ();
 sg13g2_decap_8 FILLER_159_498 ();
 sg13g2_decap_8 FILLER_159_505 ();
 sg13g2_decap_8 FILLER_159_512 ();
 sg13g2_decap_8 FILLER_159_519 ();
 sg13g2_decap_8 FILLER_159_526 ();
 sg13g2_decap_4 FILLER_159_533 ();
 sg13g2_fill_2 FILLER_159_537 ();
 sg13g2_decap_4 FILLER_159_544 ();
 sg13g2_fill_1 FILLER_159_548 ();
 sg13g2_decap_8 FILLER_159_557 ();
 sg13g2_decap_8 FILLER_159_564 ();
 sg13g2_fill_2 FILLER_159_571 ();
 sg13g2_decap_8 FILLER_159_590 ();
 sg13g2_decap_8 FILLER_159_597 ();
 sg13g2_decap_8 FILLER_159_604 ();
 sg13g2_decap_8 FILLER_159_611 ();
 sg13g2_decap_8 FILLER_159_618 ();
 sg13g2_decap_8 FILLER_159_625 ();
 sg13g2_decap_4 FILLER_159_632 ();
 sg13g2_fill_1 FILLER_159_648 ();
 sg13g2_decap_8 FILLER_159_658 ();
 sg13g2_decap_8 FILLER_159_665 ();
 sg13g2_decap_8 FILLER_159_672 ();
 sg13g2_decap_8 FILLER_159_679 ();
 sg13g2_decap_4 FILLER_159_686 ();
 sg13g2_decap_8 FILLER_159_706 ();
 sg13g2_fill_2 FILLER_159_721 ();
 sg13g2_decap_8 FILLER_159_728 ();
 sg13g2_decap_8 FILLER_159_735 ();
 sg13g2_decap_8 FILLER_159_742 ();
 sg13g2_decap_8 FILLER_159_749 ();
 sg13g2_decap_4 FILLER_159_756 ();
 sg13g2_fill_1 FILLER_159_760 ();
 sg13g2_decap_8 FILLER_159_769 ();
 sg13g2_decap_4 FILLER_159_776 ();
 sg13g2_fill_2 FILLER_159_780 ();
 sg13g2_decap_8 FILLER_159_790 ();
 sg13g2_decap_8 FILLER_159_797 ();
 sg13g2_decap_8 FILLER_159_804 ();
 sg13g2_decap_8 FILLER_159_811 ();
 sg13g2_decap_8 FILLER_159_818 ();
 sg13g2_fill_2 FILLER_159_825 ();
 sg13g2_fill_1 FILLER_159_827 ();
 sg13g2_decap_8 FILLER_159_838 ();
 sg13g2_fill_1 FILLER_159_845 ();
 sg13g2_fill_2 FILLER_159_854 ();
 sg13g2_fill_1 FILLER_159_864 ();
 sg13g2_decap_8 FILLER_159_870 ();
 sg13g2_decap_8 FILLER_159_877 ();
 sg13g2_decap_8 FILLER_159_884 ();
 sg13g2_decap_8 FILLER_159_891 ();
 sg13g2_decap_8 FILLER_159_898 ();
 sg13g2_decap_8 FILLER_159_905 ();
 sg13g2_fill_2 FILLER_159_912 ();
 sg13g2_decap_8 FILLER_159_924 ();
 sg13g2_decap_8 FILLER_159_931 ();
 sg13g2_decap_8 FILLER_159_938 ();
 sg13g2_decap_8 FILLER_159_945 ();
 sg13g2_decap_8 FILLER_159_952 ();
 sg13g2_decap_8 FILLER_159_959 ();
 sg13g2_decap_8 FILLER_159_966 ();
 sg13g2_decap_8 FILLER_159_973 ();
 sg13g2_decap_8 FILLER_159_980 ();
 sg13g2_decap_8 FILLER_159_987 ();
 sg13g2_decap_8 FILLER_159_994 ();
 sg13g2_decap_8 FILLER_159_1001 ();
 sg13g2_decap_8 FILLER_159_1008 ();
 sg13g2_decap_8 FILLER_159_1015 ();
 sg13g2_decap_4 FILLER_159_1032 ();
 sg13g2_decap_8 FILLER_159_1049 ();
 sg13g2_decap_8 FILLER_159_1056 ();
 sg13g2_decap_8 FILLER_159_1063 ();
 sg13g2_decap_8 FILLER_159_1070 ();
 sg13g2_fill_1 FILLER_159_1077 ();
 sg13g2_decap_8 FILLER_159_1086 ();
 sg13g2_decap_8 FILLER_159_1093 ();
 sg13g2_decap_4 FILLER_159_1100 ();
 sg13g2_fill_1 FILLER_159_1104 ();
 sg13g2_fill_2 FILLER_159_1114 ();
 sg13g2_fill_1 FILLER_159_1116 ();
 sg13g2_decap_8 FILLER_159_1125 ();
 sg13g2_decap_8 FILLER_159_1132 ();
 sg13g2_decap_8 FILLER_159_1139 ();
 sg13g2_decap_8 FILLER_159_1146 ();
 sg13g2_decap_4 FILLER_159_1153 ();
 sg13g2_decap_8 FILLER_159_1185 ();
 sg13g2_decap_4 FILLER_159_1192 ();
 sg13g2_fill_2 FILLER_159_1196 ();
 sg13g2_decap_8 FILLER_159_1206 ();
 sg13g2_decap_8 FILLER_159_1213 ();
 sg13g2_decap_8 FILLER_159_1220 ();
 sg13g2_decap_8 FILLER_159_1227 ();
 sg13g2_decap_8 FILLER_159_1234 ();
 sg13g2_decap_8 FILLER_159_1241 ();
 sg13g2_decap_8 FILLER_159_1248 ();
 sg13g2_decap_8 FILLER_159_1255 ();
 sg13g2_fill_1 FILLER_159_1262 ();
 sg13g2_decap_4 FILLER_159_1266 ();
 sg13g2_fill_1 FILLER_159_1270 ();
 sg13g2_decap_4 FILLER_159_1280 ();
 sg13g2_fill_2 FILLER_159_1284 ();
 sg13g2_decap_8 FILLER_159_1294 ();
 sg13g2_decap_8 FILLER_159_1301 ();
 sg13g2_decap_8 FILLER_159_1308 ();
 sg13g2_decap_8 FILLER_159_1315 ();
 sg13g2_decap_8 FILLER_159_1322 ();
 sg13g2_decap_8 FILLER_159_1329 ();
 sg13g2_decap_8 FILLER_159_1336 ();
 sg13g2_decap_8 FILLER_159_1343 ();
 sg13g2_decap_4 FILLER_159_1350 ();
 sg13g2_fill_2 FILLER_159_1354 ();
 sg13g2_fill_1 FILLER_159_1365 ();
 sg13g2_decap_8 FILLER_159_1390 ();
 sg13g2_decap_8 FILLER_159_1397 ();
 sg13g2_decap_4 FILLER_159_1404 ();
 sg13g2_fill_2 FILLER_159_1408 ();
 sg13g2_decap_8 FILLER_159_1415 ();
 sg13g2_decap_4 FILLER_159_1422 ();
 sg13g2_fill_2 FILLER_159_1426 ();
 sg13g2_decap_8 FILLER_159_1437 ();
 sg13g2_decap_8 FILLER_159_1444 ();
 sg13g2_decap_8 FILLER_159_1451 ();
 sg13g2_decap_8 FILLER_159_1458 ();
 sg13g2_decap_8 FILLER_159_1465 ();
 sg13g2_decap_8 FILLER_159_1472 ();
 sg13g2_fill_1 FILLER_159_1479 ();
 sg13g2_decap_8 FILLER_159_1493 ();
 sg13g2_decap_8 FILLER_159_1500 ();
 sg13g2_decap_8 FILLER_159_1507 ();
 sg13g2_decap_8 FILLER_159_1514 ();
 sg13g2_decap_8 FILLER_159_1521 ();
 sg13g2_decap_8 FILLER_159_1528 ();
 sg13g2_decap_8 FILLER_159_1539 ();
 sg13g2_decap_8 FILLER_159_1550 ();
 sg13g2_decap_8 FILLER_159_1557 ();
 sg13g2_decap_8 FILLER_159_1564 ();
 sg13g2_decap_8 FILLER_159_1571 ();
 sg13g2_decap_8 FILLER_159_1578 ();
 sg13g2_decap_8 FILLER_159_1585 ();
 sg13g2_decap_8 FILLER_159_1592 ();
 sg13g2_decap_8 FILLER_159_1599 ();
 sg13g2_decap_8 FILLER_159_1606 ();
 sg13g2_decap_8 FILLER_159_1613 ();
 sg13g2_decap_8 FILLER_159_1620 ();
 sg13g2_decap_8 FILLER_159_1627 ();
 sg13g2_decap_8 FILLER_159_1634 ();
 sg13g2_decap_8 FILLER_159_1641 ();
 sg13g2_decap_8 FILLER_159_1648 ();
 sg13g2_decap_8 FILLER_159_1655 ();
 sg13g2_decap_8 FILLER_159_1662 ();
 sg13g2_decap_8 FILLER_159_1669 ();
 sg13g2_decap_8 FILLER_159_1676 ();
 sg13g2_decap_8 FILLER_159_1683 ();
 sg13g2_decap_8 FILLER_159_1690 ();
 sg13g2_decap_8 FILLER_159_1697 ();
 sg13g2_decap_8 FILLER_159_1704 ();
 sg13g2_decap_8 FILLER_159_1711 ();
 sg13g2_decap_8 FILLER_159_1718 ();
 sg13g2_decap_8 FILLER_159_1725 ();
 sg13g2_decap_8 FILLER_159_1732 ();
 sg13g2_decap_8 FILLER_159_1739 ();
 sg13g2_decap_8 FILLER_159_1746 ();
 sg13g2_decap_8 FILLER_159_1753 ();
 sg13g2_decap_8 FILLER_159_1760 ();
 sg13g2_fill_1 FILLER_159_1767 ();
 sg13g2_decap_8 FILLER_160_0 ();
 sg13g2_decap_8 FILLER_160_7 ();
 sg13g2_decap_8 FILLER_160_14 ();
 sg13g2_decap_8 FILLER_160_21 ();
 sg13g2_decap_8 FILLER_160_28 ();
 sg13g2_decap_8 FILLER_160_35 ();
 sg13g2_fill_1 FILLER_160_42 ();
 sg13g2_decap_8 FILLER_160_71 ();
 sg13g2_decap_8 FILLER_160_78 ();
 sg13g2_decap_8 FILLER_160_85 ();
 sg13g2_decap_8 FILLER_160_92 ();
 sg13g2_fill_2 FILLER_160_99 ();
 sg13g2_fill_2 FILLER_160_105 ();
 sg13g2_decap_8 FILLER_160_127 ();
 sg13g2_decap_8 FILLER_160_134 ();
 sg13g2_decap_8 FILLER_160_141 ();
 sg13g2_decap_8 FILLER_160_148 ();
 sg13g2_decap_4 FILLER_160_155 ();
 sg13g2_decap_8 FILLER_160_173 ();
 sg13g2_decap_8 FILLER_160_180 ();
 sg13g2_decap_8 FILLER_160_187 ();
 sg13g2_decap_8 FILLER_160_194 ();
 sg13g2_decap_8 FILLER_160_201 ();
 sg13g2_decap_8 FILLER_160_208 ();
 sg13g2_decap_8 FILLER_160_215 ();
 sg13g2_fill_1 FILLER_160_222 ();
 sg13g2_decap_8 FILLER_160_227 ();
 sg13g2_decap_8 FILLER_160_234 ();
 sg13g2_decap_8 FILLER_160_241 ();
 sg13g2_decap_8 FILLER_160_248 ();
 sg13g2_decap_8 FILLER_160_255 ();
 sg13g2_decap_8 FILLER_160_262 ();
 sg13g2_decap_8 FILLER_160_269 ();
 sg13g2_decap_8 FILLER_160_276 ();
 sg13g2_decap_8 FILLER_160_283 ();
 sg13g2_fill_1 FILLER_160_290 ();
 sg13g2_decap_8 FILLER_160_301 ();
 sg13g2_decap_8 FILLER_160_308 ();
 sg13g2_decap_8 FILLER_160_315 ();
 sg13g2_fill_1 FILLER_160_322 ();
 sg13g2_decap_4 FILLER_160_333 ();
 sg13g2_decap_8 FILLER_160_346 ();
 sg13g2_decap_8 FILLER_160_353 ();
 sg13g2_fill_1 FILLER_160_360 ();
 sg13g2_decap_8 FILLER_160_387 ();
 sg13g2_decap_8 FILLER_160_394 ();
 sg13g2_decap_8 FILLER_160_401 ();
 sg13g2_decap_8 FILLER_160_408 ();
 sg13g2_decap_8 FILLER_160_415 ();
 sg13g2_decap_8 FILLER_160_422 ();
 sg13g2_decap_8 FILLER_160_429 ();
 sg13g2_decap_4 FILLER_160_436 ();
 sg13g2_fill_2 FILLER_160_440 ();
 sg13g2_decap_8 FILLER_160_458 ();
 sg13g2_decap_8 FILLER_160_465 ();
 sg13g2_decap_8 FILLER_160_472 ();
 sg13g2_decap_8 FILLER_160_479 ();
 sg13g2_fill_1 FILLER_160_486 ();
 sg13g2_decap_8 FILLER_160_491 ();
 sg13g2_decap_8 FILLER_160_498 ();
 sg13g2_decap_8 FILLER_160_505 ();
 sg13g2_decap_8 FILLER_160_512 ();
 sg13g2_fill_2 FILLER_160_519 ();
 sg13g2_fill_1 FILLER_160_521 ();
 sg13g2_fill_2 FILLER_160_532 ();
 sg13g2_fill_1 FILLER_160_534 ();
 sg13g2_decap_8 FILLER_160_540 ();
 sg13g2_decap_8 FILLER_160_547 ();
 sg13g2_decap_8 FILLER_160_554 ();
 sg13g2_decap_8 FILLER_160_561 ();
 sg13g2_decap_8 FILLER_160_568 ();
 sg13g2_decap_8 FILLER_160_575 ();
 sg13g2_decap_4 FILLER_160_582 ();
 sg13g2_decap_8 FILLER_160_590 ();
 sg13g2_decap_8 FILLER_160_597 ();
 sg13g2_decap_8 FILLER_160_604 ();
 sg13g2_fill_2 FILLER_160_611 ();
 sg13g2_decap_8 FILLER_160_623 ();
 sg13g2_decap_4 FILLER_160_630 ();
 sg13g2_fill_2 FILLER_160_634 ();
 sg13g2_decap_8 FILLER_160_656 ();
 sg13g2_decap_8 FILLER_160_663 ();
 sg13g2_decap_8 FILLER_160_670 ();
 sg13g2_decap_8 FILLER_160_677 ();
 sg13g2_decap_8 FILLER_160_684 ();
 sg13g2_decap_4 FILLER_160_691 ();
 sg13g2_fill_1 FILLER_160_695 ();
 sg13g2_fill_2 FILLER_160_705 ();
 sg13g2_fill_1 FILLER_160_707 ();
 sg13g2_decap_4 FILLER_160_713 ();
 sg13g2_fill_2 FILLER_160_717 ();
 sg13g2_decap_4 FILLER_160_723 ();
 sg13g2_fill_1 FILLER_160_727 ();
 sg13g2_decap_8 FILLER_160_740 ();
 sg13g2_decap_8 FILLER_160_747 ();
 sg13g2_decap_8 FILLER_160_754 ();
 sg13g2_decap_8 FILLER_160_761 ();
 sg13g2_decap_8 FILLER_160_768 ();
 sg13g2_decap_8 FILLER_160_775 ();
 sg13g2_fill_2 FILLER_160_782 ();
 sg13g2_decap_8 FILLER_160_789 ();
 sg13g2_decap_8 FILLER_160_796 ();
 sg13g2_decap_8 FILLER_160_803 ();
 sg13g2_decap_8 FILLER_160_810 ();
 sg13g2_decap_4 FILLER_160_817 ();
 sg13g2_fill_1 FILLER_160_821 ();
 sg13g2_fill_2 FILLER_160_827 ();
 sg13g2_fill_1 FILLER_160_829 ();
 sg13g2_fill_2 FILLER_160_835 ();
 sg13g2_decap_8 FILLER_160_855 ();
 sg13g2_decap_8 FILLER_160_862 ();
 sg13g2_decap_8 FILLER_160_869 ();
 sg13g2_fill_1 FILLER_160_876 ();
 sg13g2_decap_4 FILLER_160_881 ();
 sg13g2_fill_1 FILLER_160_885 ();
 sg13g2_fill_2 FILLER_160_891 ();
 sg13g2_fill_1 FILLER_160_893 ();
 sg13g2_decap_8 FILLER_160_902 ();
 sg13g2_decap_4 FILLER_160_909 ();
 sg13g2_decap_8 FILLER_160_926 ();
 sg13g2_decap_8 FILLER_160_933 ();
 sg13g2_decap_8 FILLER_160_940 ();
 sg13g2_decap_8 FILLER_160_947 ();
 sg13g2_decap_8 FILLER_160_954 ();
 sg13g2_fill_2 FILLER_160_961 ();
 sg13g2_decap_4 FILLER_160_978 ();
 sg13g2_fill_2 FILLER_160_982 ();
 sg13g2_decap_8 FILLER_160_987 ();
 sg13g2_decap_8 FILLER_160_994 ();
 sg13g2_decap_8 FILLER_160_1001 ();
 sg13g2_decap_8 FILLER_160_1008 ();
 sg13g2_decap_8 FILLER_160_1015 ();
 sg13g2_fill_1 FILLER_160_1022 ();
 sg13g2_decap_4 FILLER_160_1028 ();
 sg13g2_fill_2 FILLER_160_1032 ();
 sg13g2_decap_8 FILLER_160_1052 ();
 sg13g2_decap_8 FILLER_160_1059 ();
 sg13g2_decap_8 FILLER_160_1066 ();
 sg13g2_decap_8 FILLER_160_1073 ();
 sg13g2_decap_8 FILLER_160_1080 ();
 sg13g2_decap_8 FILLER_160_1087 ();
 sg13g2_decap_8 FILLER_160_1099 ();
 sg13g2_decap_8 FILLER_160_1106 ();
 sg13g2_decap_4 FILLER_160_1113 ();
 sg13g2_fill_2 FILLER_160_1117 ();
 sg13g2_decap_8 FILLER_160_1131 ();
 sg13g2_decap_8 FILLER_160_1138 ();
 sg13g2_decap_8 FILLER_160_1145 ();
 sg13g2_decap_8 FILLER_160_1152 ();
 sg13g2_decap_4 FILLER_160_1159 ();
 sg13g2_fill_1 FILLER_160_1163 ();
 sg13g2_decap_4 FILLER_160_1172 ();
 sg13g2_decap_8 FILLER_160_1184 ();
 sg13g2_decap_8 FILLER_160_1191 ();
 sg13g2_decap_8 FILLER_160_1198 ();
 sg13g2_decap_8 FILLER_160_1205 ();
 sg13g2_decap_4 FILLER_160_1212 ();
 sg13g2_fill_2 FILLER_160_1224 ();
 sg13g2_fill_1 FILLER_160_1226 ();
 sg13g2_decap_8 FILLER_160_1248 ();
 sg13g2_decap_4 FILLER_160_1255 ();
 sg13g2_decap_8 FILLER_160_1267 ();
 sg13g2_decap_8 FILLER_160_1274 ();
 sg13g2_decap_4 FILLER_160_1281 ();
 sg13g2_fill_1 FILLER_160_1285 ();
 sg13g2_decap_4 FILLER_160_1295 ();
 sg13g2_fill_2 FILLER_160_1299 ();
 sg13g2_decap_8 FILLER_160_1319 ();
 sg13g2_decap_8 FILLER_160_1326 ();
 sg13g2_decap_4 FILLER_160_1333 ();
 sg13g2_decap_8 FILLER_160_1340 ();
 sg13g2_decap_8 FILLER_160_1347 ();
 sg13g2_decap_8 FILLER_160_1354 ();
 sg13g2_fill_2 FILLER_160_1361 ();
 sg13g2_fill_1 FILLER_160_1363 ();
 sg13g2_decap_4 FILLER_160_1369 ();
 sg13g2_fill_1 FILLER_160_1373 ();
 sg13g2_decap_8 FILLER_160_1387 ();
 sg13g2_fill_2 FILLER_160_1394 ();
 sg13g2_fill_1 FILLER_160_1396 ();
 sg13g2_fill_2 FILLER_160_1413 ();
 sg13g2_fill_1 FILLER_160_1415 ();
 sg13g2_decap_4 FILLER_160_1424 ();
 sg13g2_fill_1 FILLER_160_1428 ();
 sg13g2_decap_8 FILLER_160_1442 ();
 sg13g2_decap_8 FILLER_160_1449 ();
 sg13g2_decap_8 FILLER_160_1456 ();
 sg13g2_decap_8 FILLER_160_1463 ();
 sg13g2_decap_8 FILLER_160_1494 ();
 sg13g2_decap_8 FILLER_160_1501 ();
 sg13g2_decap_8 FILLER_160_1508 ();
 sg13g2_decap_8 FILLER_160_1515 ();
 sg13g2_decap_8 FILLER_160_1546 ();
 sg13g2_decap_8 FILLER_160_1553 ();
 sg13g2_decap_8 FILLER_160_1560 ();
 sg13g2_decap_8 FILLER_160_1567 ();
 sg13g2_decap_8 FILLER_160_1574 ();
 sg13g2_decap_8 FILLER_160_1581 ();
 sg13g2_decap_8 FILLER_160_1588 ();
 sg13g2_decap_8 FILLER_160_1595 ();
 sg13g2_decap_8 FILLER_160_1602 ();
 sg13g2_decap_8 FILLER_160_1609 ();
 sg13g2_decap_8 FILLER_160_1616 ();
 sg13g2_decap_8 FILLER_160_1623 ();
 sg13g2_decap_8 FILLER_160_1630 ();
 sg13g2_decap_8 FILLER_160_1637 ();
 sg13g2_decap_8 FILLER_160_1644 ();
 sg13g2_decap_8 FILLER_160_1651 ();
 sg13g2_decap_8 FILLER_160_1658 ();
 sg13g2_decap_8 FILLER_160_1665 ();
 sg13g2_decap_8 FILLER_160_1672 ();
 sg13g2_decap_8 FILLER_160_1679 ();
 sg13g2_decap_8 FILLER_160_1686 ();
 sg13g2_decap_8 FILLER_160_1693 ();
 sg13g2_decap_8 FILLER_160_1700 ();
 sg13g2_decap_8 FILLER_160_1707 ();
 sg13g2_decap_8 FILLER_160_1714 ();
 sg13g2_decap_8 FILLER_160_1721 ();
 sg13g2_decap_8 FILLER_160_1728 ();
 sg13g2_decap_8 FILLER_160_1735 ();
 sg13g2_decap_8 FILLER_160_1742 ();
 sg13g2_decap_8 FILLER_160_1749 ();
 sg13g2_decap_8 FILLER_160_1756 ();
 sg13g2_decap_4 FILLER_160_1763 ();
 sg13g2_fill_1 FILLER_160_1767 ();
 sg13g2_decap_8 FILLER_161_0 ();
 sg13g2_decap_8 FILLER_161_7 ();
 sg13g2_decap_8 FILLER_161_14 ();
 sg13g2_decap_8 FILLER_161_21 ();
 sg13g2_decap_8 FILLER_161_28 ();
 sg13g2_decap_8 FILLER_161_35 ();
 sg13g2_decap_4 FILLER_161_42 ();
 sg13g2_fill_2 FILLER_161_46 ();
 sg13g2_decap_8 FILLER_161_74 ();
 sg13g2_decap_8 FILLER_161_81 ();
 sg13g2_decap_8 FILLER_161_88 ();
 sg13g2_decap_8 FILLER_161_95 ();
 sg13g2_fill_2 FILLER_161_102 ();
 sg13g2_fill_1 FILLER_161_104 ();
 sg13g2_decap_8 FILLER_161_133 ();
 sg13g2_decap_8 FILLER_161_140 ();
 sg13g2_decap_8 FILLER_161_147 ();
 sg13g2_decap_4 FILLER_161_154 ();
 sg13g2_fill_1 FILLER_161_158 ();
 sg13g2_decap_8 FILLER_161_168 ();
 sg13g2_decap_8 FILLER_161_175 ();
 sg13g2_decap_8 FILLER_161_182 ();
 sg13g2_decap_8 FILLER_161_189 ();
 sg13g2_decap_8 FILLER_161_196 ();
 sg13g2_decap_8 FILLER_161_203 ();
 sg13g2_decap_8 FILLER_161_210 ();
 sg13g2_decap_8 FILLER_161_217 ();
 sg13g2_decap_8 FILLER_161_224 ();
 sg13g2_decap_8 FILLER_161_231 ();
 sg13g2_decap_8 FILLER_161_238 ();
 sg13g2_decap_8 FILLER_161_245 ();
 sg13g2_decap_8 FILLER_161_252 ();
 sg13g2_decap_8 FILLER_161_259 ();
 sg13g2_decap_8 FILLER_161_266 ();
 sg13g2_fill_2 FILLER_161_273 ();
 sg13g2_fill_1 FILLER_161_275 ();
 sg13g2_decap_8 FILLER_161_311 ();
 sg13g2_decap_4 FILLER_161_318 ();
 sg13g2_fill_2 FILLER_161_322 ();
 sg13g2_decap_4 FILLER_161_350 ();
 sg13g2_fill_2 FILLER_161_354 ();
 sg13g2_decap_8 FILLER_161_361 ();
 sg13g2_decap_8 FILLER_161_368 ();
 sg13g2_decap_4 FILLER_161_375 ();
 sg13g2_decap_8 FILLER_161_388 ();
 sg13g2_decap_8 FILLER_161_395 ();
 sg13g2_decap_8 FILLER_161_402 ();
 sg13g2_fill_2 FILLER_161_409 ();
 sg13g2_decap_8 FILLER_161_427 ();
 sg13g2_decap_8 FILLER_161_434 ();
 sg13g2_decap_8 FILLER_161_441 ();
 sg13g2_fill_1 FILLER_161_448 ();
 sg13g2_fill_2 FILLER_161_461 ();
 sg13g2_fill_1 FILLER_161_463 ();
 sg13g2_decap_8 FILLER_161_472 ();
 sg13g2_decap_8 FILLER_161_479 ();
 sg13g2_decap_8 FILLER_161_486 ();
 sg13g2_fill_2 FILLER_161_493 ();
 sg13g2_fill_2 FILLER_161_499 ();
 sg13g2_fill_1 FILLER_161_501 ();
 sg13g2_decap_8 FILLER_161_507 ();
 sg13g2_fill_2 FILLER_161_514 ();
 sg13g2_decap_8 FILLER_161_526 ();
 sg13g2_decap_8 FILLER_161_533 ();
 sg13g2_fill_1 FILLER_161_540 ();
 sg13g2_decap_8 FILLER_161_552 ();
 sg13g2_decap_8 FILLER_161_559 ();
 sg13g2_decap_8 FILLER_161_566 ();
 sg13g2_decap_4 FILLER_161_573 ();
 sg13g2_fill_1 FILLER_161_577 ();
 sg13g2_decap_8 FILLER_161_598 ();
 sg13g2_decap_8 FILLER_161_605 ();
 sg13g2_fill_1 FILLER_161_612 ();
 sg13g2_decap_8 FILLER_161_621 ();
 sg13g2_fill_2 FILLER_161_628 ();
 sg13g2_fill_1 FILLER_161_630 ();
 sg13g2_decap_8 FILLER_161_652 ();
 sg13g2_decap_8 FILLER_161_659 ();
 sg13g2_decap_8 FILLER_161_666 ();
 sg13g2_decap_8 FILLER_161_673 ();
 sg13g2_decap_8 FILLER_161_680 ();
 sg13g2_decap_8 FILLER_161_687 ();
 sg13g2_fill_2 FILLER_161_694 ();
 sg13g2_fill_1 FILLER_161_696 ();
 sg13g2_decap_8 FILLER_161_718 ();
 sg13g2_decap_8 FILLER_161_725 ();
 sg13g2_decap_8 FILLER_161_732 ();
 sg13g2_decap_8 FILLER_161_739 ();
 sg13g2_decap_8 FILLER_161_746 ();
 sg13g2_decap_8 FILLER_161_753 ();
 sg13g2_decap_8 FILLER_161_760 ();
 sg13g2_decap_8 FILLER_161_767 ();
 sg13g2_decap_8 FILLER_161_774 ();
 sg13g2_decap_8 FILLER_161_809 ();
 sg13g2_fill_2 FILLER_161_816 ();
 sg13g2_decap_8 FILLER_161_826 ();
 sg13g2_decap_8 FILLER_161_833 ();
 sg13g2_decap_8 FILLER_161_840 ();
 sg13g2_decap_8 FILLER_161_847 ();
 sg13g2_decap_8 FILLER_161_854 ();
 sg13g2_decap_8 FILLER_161_861 ();
 sg13g2_decap_8 FILLER_161_868 ();
 sg13g2_decap_8 FILLER_161_875 ();
 sg13g2_decap_8 FILLER_161_882 ();
 sg13g2_decap_4 FILLER_161_889 ();
 sg13g2_fill_2 FILLER_161_893 ();
 sg13g2_decap_8 FILLER_161_915 ();
 sg13g2_decap_8 FILLER_161_922 ();
 sg13g2_decap_8 FILLER_161_929 ();
 sg13g2_decap_8 FILLER_161_936 ();
 sg13g2_decap_8 FILLER_161_943 ();
 sg13g2_decap_8 FILLER_161_950 ();
 sg13g2_decap_8 FILLER_161_957 ();
 sg13g2_decap_4 FILLER_161_964 ();
 sg13g2_fill_1 FILLER_161_981 ();
 sg13g2_decap_8 FILLER_161_998 ();
 sg13g2_decap_8 FILLER_161_1005 ();
 sg13g2_fill_2 FILLER_161_1012 ();
 sg13g2_fill_1 FILLER_161_1014 ();
 sg13g2_fill_2 FILLER_161_1030 ();
 sg13g2_decap_8 FILLER_161_1048 ();
 sg13g2_decap_8 FILLER_161_1055 ();
 sg13g2_decap_8 FILLER_161_1062 ();
 sg13g2_decap_8 FILLER_161_1069 ();
 sg13g2_decap_8 FILLER_161_1076 ();
 sg13g2_fill_2 FILLER_161_1083 ();
 sg13g2_fill_1 FILLER_161_1085 ();
 sg13g2_decap_8 FILLER_161_1104 ();
 sg13g2_decap_8 FILLER_161_1111 ();
 sg13g2_decap_4 FILLER_161_1118 ();
 sg13g2_fill_1 FILLER_161_1122 ();
 sg13g2_decap_8 FILLER_161_1131 ();
 sg13g2_decap_8 FILLER_161_1138 ();
 sg13g2_decap_8 FILLER_161_1145 ();
 sg13g2_decap_8 FILLER_161_1152 ();
 sg13g2_decap_8 FILLER_161_1159 ();
 sg13g2_decap_8 FILLER_161_1175 ();
 sg13g2_decap_8 FILLER_161_1182 ();
 sg13g2_decap_8 FILLER_161_1189 ();
 sg13g2_fill_2 FILLER_161_1196 ();
 sg13g2_fill_1 FILLER_161_1198 ();
 sg13g2_decap_8 FILLER_161_1207 ();
 sg13g2_decap_8 FILLER_161_1214 ();
 sg13g2_fill_2 FILLER_161_1221 ();
 sg13g2_fill_1 FILLER_161_1223 ();
 sg13g2_decap_8 FILLER_161_1243 ();
 sg13g2_decap_8 FILLER_161_1250 ();
 sg13g2_decap_8 FILLER_161_1257 ();
 sg13g2_decap_8 FILLER_161_1264 ();
 sg13g2_fill_1 FILLER_161_1271 ();
 sg13g2_fill_2 FILLER_161_1284 ();
 sg13g2_decap_8 FILLER_161_1310 ();
 sg13g2_decap_8 FILLER_161_1317 ();
 sg13g2_decap_8 FILLER_161_1332 ();
 sg13g2_decap_8 FILLER_161_1339 ();
 sg13g2_decap_8 FILLER_161_1346 ();
 sg13g2_decap_8 FILLER_161_1353 ();
 sg13g2_fill_1 FILLER_161_1360 ();
 sg13g2_fill_2 FILLER_161_1374 ();
 sg13g2_decap_8 FILLER_161_1381 ();
 sg13g2_decap_8 FILLER_161_1388 ();
 sg13g2_decap_8 FILLER_161_1395 ();
 sg13g2_decap_8 FILLER_161_1402 ();
 sg13g2_decap_8 FILLER_161_1409 ();
 sg13g2_decap_8 FILLER_161_1416 ();
 sg13g2_fill_1 FILLER_161_1423 ();
 sg13g2_decap_8 FILLER_161_1439 ();
 sg13g2_decap_8 FILLER_161_1446 ();
 sg13g2_decap_8 FILLER_161_1453 ();
 sg13g2_decap_8 FILLER_161_1460 ();
 sg13g2_decap_8 FILLER_161_1467 ();
 sg13g2_decap_4 FILLER_161_1474 ();
 sg13g2_decap_8 FILLER_161_1483 ();
 sg13g2_decap_4 FILLER_161_1490 ();
 sg13g2_fill_1 FILLER_161_1494 ();
 sg13g2_decap_8 FILLER_161_1500 ();
 sg13g2_decap_8 FILLER_161_1507 ();
 sg13g2_decap_8 FILLER_161_1514 ();
 sg13g2_decap_4 FILLER_161_1521 ();
 sg13g2_fill_2 FILLER_161_1525 ();
 sg13g2_decap_8 FILLER_161_1539 ();
 sg13g2_decap_8 FILLER_161_1546 ();
 sg13g2_decap_8 FILLER_161_1553 ();
 sg13g2_decap_8 FILLER_161_1560 ();
 sg13g2_decap_8 FILLER_161_1567 ();
 sg13g2_decap_8 FILLER_161_1574 ();
 sg13g2_decap_8 FILLER_161_1581 ();
 sg13g2_decap_8 FILLER_161_1588 ();
 sg13g2_decap_8 FILLER_161_1595 ();
 sg13g2_decap_8 FILLER_161_1602 ();
 sg13g2_decap_8 FILLER_161_1609 ();
 sg13g2_decap_8 FILLER_161_1616 ();
 sg13g2_decap_8 FILLER_161_1623 ();
 sg13g2_decap_8 FILLER_161_1630 ();
 sg13g2_decap_8 FILLER_161_1637 ();
 sg13g2_decap_8 FILLER_161_1644 ();
 sg13g2_decap_8 FILLER_161_1651 ();
 sg13g2_decap_8 FILLER_161_1658 ();
 sg13g2_decap_8 FILLER_161_1665 ();
 sg13g2_decap_8 FILLER_161_1672 ();
 sg13g2_decap_8 FILLER_161_1679 ();
 sg13g2_decap_8 FILLER_161_1686 ();
 sg13g2_decap_8 FILLER_161_1693 ();
 sg13g2_decap_8 FILLER_161_1700 ();
 sg13g2_decap_8 FILLER_161_1707 ();
 sg13g2_decap_8 FILLER_161_1714 ();
 sg13g2_decap_8 FILLER_161_1721 ();
 sg13g2_decap_8 FILLER_161_1728 ();
 sg13g2_decap_8 FILLER_161_1735 ();
 sg13g2_decap_8 FILLER_161_1742 ();
 sg13g2_decap_8 FILLER_161_1749 ();
 sg13g2_decap_8 FILLER_161_1756 ();
 sg13g2_decap_4 FILLER_161_1763 ();
 sg13g2_fill_1 FILLER_161_1767 ();
 sg13g2_decap_8 FILLER_162_0 ();
 sg13g2_decap_8 FILLER_162_7 ();
 sg13g2_decap_8 FILLER_162_14 ();
 sg13g2_decap_8 FILLER_162_21 ();
 sg13g2_decap_8 FILLER_162_28 ();
 sg13g2_decap_8 FILLER_162_35 ();
 sg13g2_decap_8 FILLER_162_42 ();
 sg13g2_fill_2 FILLER_162_49 ();
 sg13g2_fill_1 FILLER_162_51 ();
 sg13g2_decap_8 FILLER_162_82 ();
 sg13g2_decap_8 FILLER_162_89 ();
 sg13g2_decap_8 FILLER_162_96 ();
 sg13g2_fill_2 FILLER_162_103 ();
 sg13g2_fill_1 FILLER_162_105 ();
 sg13g2_fill_2 FILLER_162_116 ();
 sg13g2_decap_8 FILLER_162_136 ();
 sg13g2_decap_8 FILLER_162_143 ();
 sg13g2_decap_8 FILLER_162_150 ();
 sg13g2_decap_8 FILLER_162_157 ();
 sg13g2_decap_8 FILLER_162_164 ();
 sg13g2_decap_8 FILLER_162_171 ();
 sg13g2_decap_8 FILLER_162_178 ();
 sg13g2_decap_8 FILLER_162_185 ();
 sg13g2_decap_8 FILLER_162_192 ();
 sg13g2_decap_8 FILLER_162_199 ();
 sg13g2_decap_8 FILLER_162_206 ();
 sg13g2_decap_8 FILLER_162_213 ();
 sg13g2_decap_8 FILLER_162_220 ();
 sg13g2_decap_4 FILLER_162_227 ();
 sg13g2_fill_1 FILLER_162_231 ();
 sg13g2_fill_2 FILLER_162_237 ();
 sg13g2_decap_8 FILLER_162_249 ();
 sg13g2_decap_8 FILLER_162_256 ();
 sg13g2_decap_8 FILLER_162_263 ();
 sg13g2_decap_8 FILLER_162_270 ();
 sg13g2_decap_8 FILLER_162_277 ();
 sg13g2_fill_2 FILLER_162_284 ();
 sg13g2_decap_8 FILLER_162_290 ();
 sg13g2_decap_8 FILLER_162_297 ();
 sg13g2_decap_8 FILLER_162_304 ();
 sg13g2_decap_8 FILLER_162_311 ();
 sg13g2_decap_8 FILLER_162_318 ();
 sg13g2_fill_1 FILLER_162_325 ();
 sg13g2_fill_1 FILLER_162_334 ();
 sg13g2_decap_8 FILLER_162_339 ();
 sg13g2_decap_8 FILLER_162_346 ();
 sg13g2_decap_8 FILLER_162_353 ();
 sg13g2_decap_8 FILLER_162_360 ();
 sg13g2_decap_8 FILLER_162_367 ();
 sg13g2_decap_4 FILLER_162_374 ();
 sg13g2_fill_1 FILLER_162_378 ();
 sg13g2_decap_4 FILLER_162_384 ();
 sg13g2_fill_1 FILLER_162_388 ();
 sg13g2_decap_8 FILLER_162_399 ();
 sg13g2_decap_4 FILLER_162_406 ();
 sg13g2_fill_2 FILLER_162_418 ();
 sg13g2_decap_4 FILLER_162_428 ();
 sg13g2_fill_1 FILLER_162_432 ();
 sg13g2_decap_4 FILLER_162_449 ();
 sg13g2_fill_2 FILLER_162_453 ();
 sg13g2_fill_2 FILLER_162_459 ();
 sg13g2_fill_1 FILLER_162_461 ();
 sg13g2_decap_8 FILLER_162_467 ();
 sg13g2_decap_8 FILLER_162_474 ();
 sg13g2_fill_2 FILLER_162_481 ();
 sg13g2_fill_2 FILLER_162_493 ();
 sg13g2_fill_1 FILLER_162_495 ();
 sg13g2_fill_2 FILLER_162_504 ();
 sg13g2_fill_1 FILLER_162_506 ();
 sg13g2_decap_8 FILLER_162_515 ();
 sg13g2_decap_8 FILLER_162_522 ();
 sg13g2_decap_8 FILLER_162_529 ();
 sg13g2_decap_8 FILLER_162_536 ();
 sg13g2_decap_8 FILLER_162_543 ();
 sg13g2_fill_2 FILLER_162_550 ();
 sg13g2_fill_1 FILLER_162_552 ();
 sg13g2_decap_8 FILLER_162_561 ();
 sg13g2_decap_8 FILLER_162_568 ();
 sg13g2_decap_8 FILLER_162_575 ();
 sg13g2_decap_8 FILLER_162_582 ();
 sg13g2_decap_8 FILLER_162_589 ();
 sg13g2_fill_1 FILLER_162_596 ();
 sg13g2_decap_8 FILLER_162_605 ();
 sg13g2_decap_8 FILLER_162_612 ();
 sg13g2_decap_8 FILLER_162_619 ();
 sg13g2_decap_8 FILLER_162_626 ();
 sg13g2_decap_8 FILLER_162_640 ();
 sg13g2_decap_8 FILLER_162_647 ();
 sg13g2_decap_8 FILLER_162_654 ();
 sg13g2_decap_8 FILLER_162_661 ();
 sg13g2_decap_8 FILLER_162_668 ();
 sg13g2_decap_8 FILLER_162_675 ();
 sg13g2_decap_8 FILLER_162_682 ();
 sg13g2_decap_8 FILLER_162_689 ();
 sg13g2_decap_8 FILLER_162_696 ();
 sg13g2_decap_4 FILLER_162_703 ();
 sg13g2_fill_1 FILLER_162_707 ();
 sg13g2_decap_8 FILLER_162_716 ();
 sg13g2_decap_4 FILLER_162_723 ();
 sg13g2_decap_8 FILLER_162_743 ();
 sg13g2_decap_4 FILLER_162_750 ();
 sg13g2_fill_2 FILLER_162_754 ();
 sg13g2_decap_8 FILLER_162_760 ();
 sg13g2_fill_2 FILLER_162_767 ();
 sg13g2_fill_1 FILLER_162_769 ();
 sg13g2_decap_4 FILLER_162_775 ();
 sg13g2_fill_1 FILLER_162_792 ();
 sg13g2_decap_8 FILLER_162_815 ();
 sg13g2_decap_8 FILLER_162_822 ();
 sg13g2_decap_4 FILLER_162_829 ();
 sg13g2_fill_2 FILLER_162_833 ();
 sg13g2_fill_1 FILLER_162_844 ();
 sg13g2_decap_8 FILLER_162_857 ();
 sg13g2_decap_8 FILLER_162_864 ();
 sg13g2_decap_8 FILLER_162_871 ();
 sg13g2_decap_8 FILLER_162_890 ();
 sg13g2_decap_8 FILLER_162_897 ();
 sg13g2_decap_8 FILLER_162_904 ();
 sg13g2_decap_8 FILLER_162_911 ();
 sg13g2_decap_8 FILLER_162_918 ();
 sg13g2_decap_8 FILLER_162_925 ();
 sg13g2_decap_8 FILLER_162_932 ();
 sg13g2_decap_8 FILLER_162_939 ();
 sg13g2_decap_8 FILLER_162_946 ();
 sg13g2_decap_8 FILLER_162_953 ();
 sg13g2_decap_8 FILLER_162_960 ();
 sg13g2_decap_8 FILLER_162_967 ();
 sg13g2_decap_8 FILLER_162_974 ();
 sg13g2_fill_2 FILLER_162_981 ();
 sg13g2_fill_1 FILLER_162_983 ();
 sg13g2_decap_8 FILLER_162_1005 ();
 sg13g2_decap_8 FILLER_162_1012 ();
 sg13g2_fill_2 FILLER_162_1019 ();
 sg13g2_decap_8 FILLER_162_1030 ();
 sg13g2_decap_8 FILLER_162_1037 ();
 sg13g2_decap_8 FILLER_162_1044 ();
 sg13g2_decap_8 FILLER_162_1051 ();
 sg13g2_decap_8 FILLER_162_1058 ();
 sg13g2_decap_8 FILLER_162_1065 ();
 sg13g2_decap_8 FILLER_162_1072 ();
 sg13g2_fill_1 FILLER_162_1079 ();
 sg13g2_decap_8 FILLER_162_1088 ();
 sg13g2_decap_8 FILLER_162_1095 ();
 sg13g2_decap_4 FILLER_162_1102 ();
 sg13g2_decap_8 FILLER_162_1119 ();
 sg13g2_decap_8 FILLER_162_1126 ();
 sg13g2_decap_8 FILLER_162_1133 ();
 sg13g2_decap_8 FILLER_162_1140 ();
 sg13g2_decap_8 FILLER_162_1147 ();
 sg13g2_decap_4 FILLER_162_1154 ();
 sg13g2_decap_8 FILLER_162_1179 ();
 sg13g2_decap_8 FILLER_162_1186 ();
 sg13g2_decap_4 FILLER_162_1193 ();
 sg13g2_fill_2 FILLER_162_1197 ();
 sg13g2_decap_8 FILLER_162_1212 ();
 sg13g2_decap_4 FILLER_162_1219 ();
 sg13g2_decap_4 FILLER_162_1228 ();
 sg13g2_fill_2 FILLER_162_1232 ();
 sg13g2_decap_8 FILLER_162_1242 ();
 sg13g2_decap_8 FILLER_162_1249 ();
 sg13g2_decap_8 FILLER_162_1256 ();
 sg13g2_decap_4 FILLER_162_1263 ();
 sg13g2_fill_2 FILLER_162_1267 ();
 sg13g2_decap_4 FILLER_162_1274 ();
 sg13g2_fill_2 FILLER_162_1282 ();
 sg13g2_fill_1 FILLER_162_1284 ();
 sg13g2_decap_8 FILLER_162_1297 ();
 sg13g2_decap_8 FILLER_162_1304 ();
 sg13g2_decap_8 FILLER_162_1311 ();
 sg13g2_decap_8 FILLER_162_1318 ();
 sg13g2_decap_8 FILLER_162_1325 ();
 sg13g2_decap_8 FILLER_162_1332 ();
 sg13g2_decap_8 FILLER_162_1339 ();
 sg13g2_decap_4 FILLER_162_1346 ();
 sg13g2_decap_8 FILLER_162_1353 ();
 sg13g2_decap_8 FILLER_162_1360 ();
 sg13g2_decap_4 FILLER_162_1367 ();
 sg13g2_fill_1 FILLER_162_1371 ();
 sg13g2_decap_8 FILLER_162_1375 ();
 sg13g2_decap_8 FILLER_162_1382 ();
 sg13g2_decap_8 FILLER_162_1389 ();
 sg13g2_decap_8 FILLER_162_1396 ();
 sg13g2_decap_4 FILLER_162_1403 ();
 sg13g2_fill_2 FILLER_162_1415 ();
 sg13g2_fill_1 FILLER_162_1417 ();
 sg13g2_decap_8 FILLER_162_1426 ();
 sg13g2_decap_8 FILLER_162_1433 ();
 sg13g2_decap_8 FILLER_162_1440 ();
 sg13g2_decap_8 FILLER_162_1447 ();
 sg13g2_decap_8 FILLER_162_1454 ();
 sg13g2_decap_8 FILLER_162_1461 ();
 sg13g2_decap_8 FILLER_162_1468 ();
 sg13g2_fill_2 FILLER_162_1475 ();
 sg13g2_decap_4 FILLER_162_1480 ();
 sg13g2_fill_2 FILLER_162_1484 ();
 sg13g2_decap_8 FILLER_162_1508 ();
 sg13g2_fill_2 FILLER_162_1515 ();
 sg13g2_decap_8 FILLER_162_1520 ();
 sg13g2_decap_8 FILLER_162_1527 ();
 sg13g2_decap_8 FILLER_162_1534 ();
 sg13g2_decap_8 FILLER_162_1541 ();
 sg13g2_decap_8 FILLER_162_1548 ();
 sg13g2_decap_8 FILLER_162_1555 ();
 sg13g2_decap_8 FILLER_162_1562 ();
 sg13g2_decap_8 FILLER_162_1569 ();
 sg13g2_decap_8 FILLER_162_1576 ();
 sg13g2_decap_8 FILLER_162_1583 ();
 sg13g2_decap_8 FILLER_162_1590 ();
 sg13g2_decap_8 FILLER_162_1597 ();
 sg13g2_decap_8 FILLER_162_1604 ();
 sg13g2_decap_8 FILLER_162_1611 ();
 sg13g2_decap_8 FILLER_162_1618 ();
 sg13g2_decap_8 FILLER_162_1625 ();
 sg13g2_decap_8 FILLER_162_1632 ();
 sg13g2_decap_8 FILLER_162_1639 ();
 sg13g2_decap_8 FILLER_162_1646 ();
 sg13g2_decap_8 FILLER_162_1653 ();
 sg13g2_decap_8 FILLER_162_1660 ();
 sg13g2_decap_8 FILLER_162_1667 ();
 sg13g2_decap_8 FILLER_162_1674 ();
 sg13g2_decap_8 FILLER_162_1681 ();
 sg13g2_decap_8 FILLER_162_1688 ();
 sg13g2_decap_8 FILLER_162_1695 ();
 sg13g2_decap_8 FILLER_162_1702 ();
 sg13g2_decap_8 FILLER_162_1709 ();
 sg13g2_decap_8 FILLER_162_1716 ();
 sg13g2_decap_8 FILLER_162_1723 ();
 sg13g2_decap_8 FILLER_162_1730 ();
 sg13g2_decap_8 FILLER_162_1737 ();
 sg13g2_decap_8 FILLER_162_1744 ();
 sg13g2_decap_8 FILLER_162_1751 ();
 sg13g2_decap_8 FILLER_162_1758 ();
 sg13g2_fill_2 FILLER_162_1765 ();
 sg13g2_fill_1 FILLER_162_1767 ();
 sg13g2_decap_8 FILLER_163_0 ();
 sg13g2_decap_8 FILLER_163_7 ();
 sg13g2_decap_8 FILLER_163_14 ();
 sg13g2_decap_8 FILLER_163_21 ();
 sg13g2_decap_8 FILLER_163_28 ();
 sg13g2_decap_8 FILLER_163_35 ();
 sg13g2_decap_8 FILLER_163_42 ();
 sg13g2_decap_8 FILLER_163_49 ();
 sg13g2_decap_4 FILLER_163_56 ();
 sg13g2_decap_8 FILLER_163_76 ();
 sg13g2_decap_8 FILLER_163_83 ();
 sg13g2_decap_8 FILLER_163_90 ();
 sg13g2_decap_8 FILLER_163_97 ();
 sg13g2_decap_8 FILLER_163_104 ();
 sg13g2_fill_1 FILLER_163_111 ();
 sg13g2_fill_2 FILLER_163_131 ();
 sg13g2_decap_8 FILLER_163_141 ();
 sg13g2_decap_8 FILLER_163_148 ();
 sg13g2_decap_8 FILLER_163_155 ();
 sg13g2_decap_8 FILLER_163_162 ();
 sg13g2_decap_8 FILLER_163_169 ();
 sg13g2_decap_8 FILLER_163_176 ();
 sg13g2_decap_8 FILLER_163_183 ();
 sg13g2_fill_2 FILLER_163_190 ();
 sg13g2_decap_8 FILLER_163_201 ();
 sg13g2_decap_8 FILLER_163_208 ();
 sg13g2_decap_8 FILLER_163_215 ();
 sg13g2_fill_1 FILLER_163_222 ();
 sg13g2_fill_2 FILLER_163_232 ();
 sg13g2_fill_1 FILLER_163_252 ();
 sg13g2_decap_8 FILLER_163_256 ();
 sg13g2_decap_8 FILLER_163_263 ();
 sg13g2_decap_8 FILLER_163_270 ();
 sg13g2_decap_8 FILLER_163_277 ();
 sg13g2_decap_8 FILLER_163_284 ();
 sg13g2_decap_8 FILLER_163_291 ();
 sg13g2_decap_8 FILLER_163_298 ();
 sg13g2_decap_8 FILLER_163_305 ();
 sg13g2_decap_8 FILLER_163_312 ();
 sg13g2_decap_8 FILLER_163_319 ();
 sg13g2_fill_2 FILLER_163_326 ();
 sg13g2_fill_1 FILLER_163_328 ();
 sg13g2_decap_8 FILLER_163_333 ();
 sg13g2_decap_8 FILLER_163_340 ();
 sg13g2_decap_8 FILLER_163_347 ();
 sg13g2_decap_8 FILLER_163_354 ();
 sg13g2_decap_4 FILLER_163_361 ();
 sg13g2_fill_2 FILLER_163_376 ();
 sg13g2_fill_1 FILLER_163_378 ();
 sg13g2_decap_8 FILLER_163_400 ();
 sg13g2_decap_8 FILLER_163_407 ();
 sg13g2_decap_8 FILLER_163_414 ();
 sg13g2_decap_8 FILLER_163_421 ();
 sg13g2_decap_8 FILLER_163_428 ();
 sg13g2_fill_2 FILLER_163_435 ();
 sg13g2_decap_8 FILLER_163_450 ();
 sg13g2_decap_8 FILLER_163_457 ();
 sg13g2_decap_8 FILLER_163_464 ();
 sg13g2_decap_8 FILLER_163_471 ();
 sg13g2_decap_8 FILLER_163_478 ();
 sg13g2_decap_4 FILLER_163_488 ();
 sg13g2_fill_2 FILLER_163_492 ();
 sg13g2_fill_2 FILLER_163_498 ();
 sg13g2_decap_8 FILLER_163_517 ();
 sg13g2_decap_8 FILLER_163_524 ();
 sg13g2_decap_8 FILLER_163_531 ();
 sg13g2_fill_2 FILLER_163_538 ();
 sg13g2_fill_1 FILLER_163_540 ();
 sg13g2_decap_8 FILLER_163_558 ();
 sg13g2_decap_8 FILLER_163_565 ();
 sg13g2_decap_8 FILLER_163_572 ();
 sg13g2_decap_4 FILLER_163_579 ();
 sg13g2_fill_1 FILLER_163_583 ();
 sg13g2_decap_8 FILLER_163_587 ();
 sg13g2_decap_8 FILLER_163_598 ();
 sg13g2_decap_8 FILLER_163_605 ();
 sg13g2_fill_1 FILLER_163_612 ();
 sg13g2_decap_8 FILLER_163_617 ();
 sg13g2_decap_8 FILLER_163_624 ();
 sg13g2_decap_4 FILLER_163_631 ();
 sg13g2_decap_8 FILLER_163_643 ();
 sg13g2_decap_4 FILLER_163_650 ();
 sg13g2_decap_8 FILLER_163_663 ();
 sg13g2_decap_8 FILLER_163_670 ();
 sg13g2_decap_8 FILLER_163_677 ();
 sg13g2_decap_8 FILLER_163_684 ();
 sg13g2_decap_8 FILLER_163_691 ();
 sg13g2_decap_8 FILLER_163_698 ();
 sg13g2_decap_8 FILLER_163_705 ();
 sg13g2_decap_8 FILLER_163_712 ();
 sg13g2_decap_8 FILLER_163_719 ();
 sg13g2_decap_4 FILLER_163_726 ();
 sg13g2_fill_1 FILLER_163_730 ();
 sg13g2_decap_8 FILLER_163_740 ();
 sg13g2_fill_2 FILLER_163_747 ();
 sg13g2_fill_1 FILLER_163_749 ();
 sg13g2_fill_2 FILLER_163_767 ();
 sg13g2_fill_1 FILLER_163_769 ();
 sg13g2_decap_8 FILLER_163_774 ();
 sg13g2_decap_4 FILLER_163_781 ();
 sg13g2_fill_2 FILLER_163_785 ();
 sg13g2_decap_8 FILLER_163_799 ();
 sg13g2_decap_8 FILLER_163_806 ();
 sg13g2_decap_4 FILLER_163_813 ();
 sg13g2_decap_8 FILLER_163_825 ();
 sg13g2_decap_8 FILLER_163_832 ();
 sg13g2_decap_8 FILLER_163_839 ();
 sg13g2_decap_8 FILLER_163_863 ();
 sg13g2_decap_4 FILLER_163_870 ();
 sg13g2_fill_2 FILLER_163_874 ();
 sg13g2_decap_8 FILLER_163_884 ();
 sg13g2_decap_8 FILLER_163_891 ();
 sg13g2_decap_4 FILLER_163_898 ();
 sg13g2_fill_1 FILLER_163_902 ();
 sg13g2_fill_1 FILLER_163_911 ();
 sg13g2_decap_8 FILLER_163_920 ();
 sg13g2_decap_8 FILLER_163_927 ();
 sg13g2_decap_8 FILLER_163_934 ();
 sg13g2_decap_8 FILLER_163_941 ();
 sg13g2_decap_8 FILLER_163_948 ();
 sg13g2_decap_8 FILLER_163_955 ();
 sg13g2_decap_8 FILLER_163_962 ();
 sg13g2_decap_8 FILLER_163_969 ();
 sg13g2_decap_8 FILLER_163_976 ();
 sg13g2_fill_2 FILLER_163_983 ();
 sg13g2_fill_2 FILLER_163_997 ();
 sg13g2_fill_1 FILLER_163_999 ();
 sg13g2_decap_8 FILLER_163_1008 ();
 sg13g2_decap_8 FILLER_163_1015 ();
 sg13g2_decap_8 FILLER_163_1022 ();
 sg13g2_fill_2 FILLER_163_1029 ();
 sg13g2_fill_1 FILLER_163_1031 ();
 sg13g2_fill_1 FILLER_163_1036 ();
 sg13g2_fill_1 FILLER_163_1041 ();
 sg13g2_decap_8 FILLER_163_1047 ();
 sg13g2_decap_8 FILLER_163_1054 ();
 sg13g2_decap_8 FILLER_163_1061 ();
 sg13g2_decap_8 FILLER_163_1068 ();
 sg13g2_decap_4 FILLER_163_1075 ();
 sg13g2_fill_2 FILLER_163_1079 ();
 sg13g2_decap_8 FILLER_163_1094 ();
 sg13g2_fill_2 FILLER_163_1101 ();
 sg13g2_decap_8 FILLER_163_1124 ();
 sg13g2_decap_8 FILLER_163_1131 ();
 sg13g2_decap_8 FILLER_163_1138 ();
 sg13g2_decap_8 FILLER_163_1145 ();
 sg13g2_decap_8 FILLER_163_1152 ();
 sg13g2_decap_4 FILLER_163_1159 ();
 sg13g2_fill_1 FILLER_163_1163 ();
 sg13g2_decap_8 FILLER_163_1174 ();
 sg13g2_decap_8 FILLER_163_1181 ();
 sg13g2_decap_8 FILLER_163_1188 ();
 sg13g2_decap_8 FILLER_163_1195 ();
 sg13g2_decap_8 FILLER_163_1202 ();
 sg13g2_decap_8 FILLER_163_1209 ();
 sg13g2_decap_8 FILLER_163_1216 ();
 sg13g2_fill_1 FILLER_163_1223 ();
 sg13g2_decap_8 FILLER_163_1232 ();
 sg13g2_decap_8 FILLER_163_1239 ();
 sg13g2_decap_8 FILLER_163_1246 ();
 sg13g2_decap_8 FILLER_163_1253 ();
 sg13g2_decap_8 FILLER_163_1260 ();
 sg13g2_fill_2 FILLER_163_1267 ();
 sg13g2_fill_1 FILLER_163_1277 ();
 sg13g2_decap_8 FILLER_163_1282 ();
 sg13g2_decap_8 FILLER_163_1293 ();
 sg13g2_decap_8 FILLER_163_1300 ();
 sg13g2_decap_8 FILLER_163_1307 ();
 sg13g2_decap_8 FILLER_163_1314 ();
 sg13g2_decap_8 FILLER_163_1321 ();
 sg13g2_decap_8 FILLER_163_1328 ();
 sg13g2_decap_8 FILLER_163_1335 ();
 sg13g2_decap_8 FILLER_163_1342 ();
 sg13g2_decap_8 FILLER_163_1349 ();
 sg13g2_decap_8 FILLER_163_1356 ();
 sg13g2_decap_8 FILLER_163_1363 ();
 sg13g2_decap_8 FILLER_163_1370 ();
 sg13g2_decap_8 FILLER_163_1377 ();
 sg13g2_decap_8 FILLER_163_1384 ();
 sg13g2_decap_8 FILLER_163_1391 ();
 sg13g2_decap_8 FILLER_163_1398 ();
 sg13g2_decap_8 FILLER_163_1405 ();
 sg13g2_fill_2 FILLER_163_1412 ();
 sg13g2_decap_8 FILLER_163_1418 ();
 sg13g2_decap_4 FILLER_163_1425 ();
 sg13g2_fill_2 FILLER_163_1429 ();
 sg13g2_fill_1 FILLER_163_1436 ();
 sg13g2_fill_2 FILLER_163_1441 ();
 sg13g2_decap_8 FILLER_163_1448 ();
 sg13g2_decap_8 FILLER_163_1455 ();
 sg13g2_decap_8 FILLER_163_1462 ();
 sg13g2_fill_2 FILLER_163_1469 ();
 sg13g2_fill_2 FILLER_163_1476 ();
 sg13g2_decap_8 FILLER_163_1504 ();
 sg13g2_decap_8 FILLER_163_1511 ();
 sg13g2_decap_8 FILLER_163_1518 ();
 sg13g2_decap_8 FILLER_163_1525 ();
 sg13g2_decap_8 FILLER_163_1532 ();
 sg13g2_decap_8 FILLER_163_1539 ();
 sg13g2_decap_8 FILLER_163_1546 ();
 sg13g2_decap_8 FILLER_163_1553 ();
 sg13g2_decap_8 FILLER_163_1560 ();
 sg13g2_decap_8 FILLER_163_1567 ();
 sg13g2_decap_8 FILLER_163_1574 ();
 sg13g2_decap_8 FILLER_163_1581 ();
 sg13g2_decap_8 FILLER_163_1588 ();
 sg13g2_decap_8 FILLER_163_1595 ();
 sg13g2_decap_8 FILLER_163_1602 ();
 sg13g2_decap_8 FILLER_163_1609 ();
 sg13g2_decap_8 FILLER_163_1616 ();
 sg13g2_decap_8 FILLER_163_1623 ();
 sg13g2_decap_8 FILLER_163_1630 ();
 sg13g2_decap_8 FILLER_163_1637 ();
 sg13g2_decap_8 FILLER_163_1644 ();
 sg13g2_decap_8 FILLER_163_1651 ();
 sg13g2_decap_8 FILLER_163_1658 ();
 sg13g2_decap_8 FILLER_163_1665 ();
 sg13g2_decap_8 FILLER_163_1672 ();
 sg13g2_decap_8 FILLER_163_1679 ();
 sg13g2_decap_8 FILLER_163_1686 ();
 sg13g2_decap_8 FILLER_163_1693 ();
 sg13g2_decap_8 FILLER_163_1700 ();
 sg13g2_decap_8 FILLER_163_1707 ();
 sg13g2_decap_8 FILLER_163_1714 ();
 sg13g2_decap_8 FILLER_163_1721 ();
 sg13g2_decap_8 FILLER_163_1728 ();
 sg13g2_decap_8 FILLER_163_1735 ();
 sg13g2_decap_8 FILLER_163_1742 ();
 sg13g2_decap_8 FILLER_163_1749 ();
 sg13g2_decap_8 FILLER_163_1756 ();
 sg13g2_decap_4 FILLER_163_1763 ();
 sg13g2_fill_1 FILLER_163_1767 ();
 sg13g2_decap_8 FILLER_164_0 ();
 sg13g2_decap_8 FILLER_164_7 ();
 sg13g2_decap_8 FILLER_164_14 ();
 sg13g2_decap_8 FILLER_164_21 ();
 sg13g2_decap_8 FILLER_164_28 ();
 sg13g2_decap_8 FILLER_164_35 ();
 sg13g2_decap_8 FILLER_164_42 ();
 sg13g2_decap_8 FILLER_164_49 ();
 sg13g2_decap_8 FILLER_164_56 ();
 sg13g2_decap_8 FILLER_164_63 ();
 sg13g2_decap_8 FILLER_164_70 ();
 sg13g2_decap_8 FILLER_164_77 ();
 sg13g2_decap_8 FILLER_164_84 ();
 sg13g2_decap_8 FILLER_164_91 ();
 sg13g2_decap_8 FILLER_164_98 ();
 sg13g2_decap_8 FILLER_164_105 ();
 sg13g2_decap_4 FILLER_164_112 ();
 sg13g2_fill_2 FILLER_164_126 ();
 sg13g2_decap_8 FILLER_164_149 ();
 sg13g2_decap_8 FILLER_164_156 ();
 sg13g2_decap_8 FILLER_164_163 ();
 sg13g2_decap_8 FILLER_164_170 ();
 sg13g2_decap_4 FILLER_164_177 ();
 sg13g2_fill_2 FILLER_164_181 ();
 sg13g2_fill_2 FILLER_164_192 ();
 sg13g2_fill_1 FILLER_164_199 ();
 sg13g2_decap_8 FILLER_164_210 ();
 sg13g2_decap_8 FILLER_164_217 ();
 sg13g2_fill_1 FILLER_164_224 ();
 sg13g2_fill_1 FILLER_164_239 ();
 sg13g2_fill_1 FILLER_164_250 ();
 sg13g2_fill_1 FILLER_164_255 ();
 sg13g2_decap_8 FILLER_164_271 ();
 sg13g2_decap_8 FILLER_164_278 ();
 sg13g2_decap_8 FILLER_164_285 ();
 sg13g2_decap_8 FILLER_164_292 ();
 sg13g2_decap_8 FILLER_164_299 ();
 sg13g2_decap_8 FILLER_164_306 ();
 sg13g2_decap_4 FILLER_164_313 ();
 sg13g2_fill_1 FILLER_164_317 ();
 sg13g2_fill_2 FILLER_164_321 ();
 sg13g2_fill_1 FILLER_164_323 ();
 sg13g2_decap_8 FILLER_164_344 ();
 sg13g2_decap_8 FILLER_164_351 ();
 sg13g2_decap_8 FILLER_164_358 ();
 sg13g2_decap_8 FILLER_164_365 ();
 sg13g2_decap_8 FILLER_164_372 ();
 sg13g2_fill_1 FILLER_164_379 ();
 sg13g2_decap_8 FILLER_164_390 ();
 sg13g2_decap_8 FILLER_164_397 ();
 sg13g2_fill_1 FILLER_164_404 ();
 sg13g2_decap_8 FILLER_164_409 ();
 sg13g2_decap_8 FILLER_164_416 ();
 sg13g2_decap_8 FILLER_164_423 ();
 sg13g2_decap_8 FILLER_164_430 ();
 sg13g2_decap_8 FILLER_164_437 ();
 sg13g2_decap_8 FILLER_164_444 ();
 sg13g2_decap_8 FILLER_164_463 ();
 sg13g2_decap_8 FILLER_164_470 ();
 sg13g2_decap_8 FILLER_164_477 ();
 sg13g2_fill_2 FILLER_164_484 ();
 sg13g2_fill_1 FILLER_164_486 ();
 sg13g2_decap_4 FILLER_164_495 ();
 sg13g2_fill_1 FILLER_164_499 ();
 sg13g2_decap_4 FILLER_164_505 ();
 sg13g2_fill_1 FILLER_164_509 ();
 sg13g2_decap_8 FILLER_164_515 ();
 sg13g2_decap_8 FILLER_164_522 ();
 sg13g2_decap_8 FILLER_164_529 ();
 sg13g2_decap_4 FILLER_164_536 ();
 sg13g2_fill_1 FILLER_164_540 ();
 sg13g2_decap_8 FILLER_164_565 ();
 sg13g2_decap_8 FILLER_164_572 ();
 sg13g2_fill_2 FILLER_164_579 ();
 sg13g2_fill_1 FILLER_164_581 ();
 sg13g2_fill_2 FILLER_164_599 ();
 sg13g2_fill_1 FILLER_164_611 ();
 sg13g2_decap_8 FILLER_164_624 ();
 sg13g2_decap_8 FILLER_164_631 ();
 sg13g2_decap_8 FILLER_164_638 ();
 sg13g2_decap_8 FILLER_164_645 ();
 sg13g2_fill_2 FILLER_164_652 ();
 sg13g2_decap_8 FILLER_164_684 ();
 sg13g2_fill_2 FILLER_164_691 ();
 sg13g2_decap_4 FILLER_164_698 ();
 sg13g2_fill_2 FILLER_164_702 ();
 sg13g2_decap_8 FILLER_164_717 ();
 sg13g2_decap_8 FILLER_164_724 ();
 sg13g2_fill_1 FILLER_164_744 ();
 sg13g2_decap_4 FILLER_164_753 ();
 sg13g2_fill_1 FILLER_164_757 ();
 sg13g2_decap_8 FILLER_164_766 ();
 sg13g2_decap_8 FILLER_164_773 ();
 sg13g2_decap_8 FILLER_164_780 ();
 sg13g2_decap_8 FILLER_164_787 ();
 sg13g2_decap_8 FILLER_164_794 ();
 sg13g2_decap_8 FILLER_164_809 ();
 sg13g2_fill_2 FILLER_164_816 ();
 sg13g2_fill_1 FILLER_164_818 ();
 sg13g2_decap_8 FILLER_164_829 ();
 sg13g2_decap_8 FILLER_164_836 ();
 sg13g2_decap_8 FILLER_164_843 ();
 sg13g2_decap_8 FILLER_164_850 ();
 sg13g2_decap_8 FILLER_164_857 ();
 sg13g2_fill_2 FILLER_164_864 ();
 sg13g2_fill_2 FILLER_164_870 ();
 sg13g2_decap_8 FILLER_164_886 ();
 sg13g2_decap_8 FILLER_164_893 ();
 sg13g2_decap_8 FILLER_164_900 ();
 sg13g2_decap_4 FILLER_164_913 ();
 sg13g2_decap_8 FILLER_164_933 ();
 sg13g2_decap_8 FILLER_164_940 ();
 sg13g2_decap_8 FILLER_164_947 ();
 sg13g2_decap_8 FILLER_164_954 ();
 sg13g2_decap_8 FILLER_164_961 ();
 sg13g2_decap_4 FILLER_164_968 ();
 sg13g2_decap_8 FILLER_164_981 ();
 sg13g2_decap_4 FILLER_164_988 ();
 sg13g2_fill_1 FILLER_164_992 ();
 sg13g2_decap_8 FILLER_164_997 ();
 sg13g2_decap_8 FILLER_164_1004 ();
 sg13g2_decap_8 FILLER_164_1011 ();
 sg13g2_fill_1 FILLER_164_1018 ();
 sg13g2_decap_8 FILLER_164_1053 ();
 sg13g2_decap_8 FILLER_164_1060 ();
 sg13g2_decap_8 FILLER_164_1067 ();
 sg13g2_decap_8 FILLER_164_1074 ();
 sg13g2_decap_4 FILLER_164_1081 ();
 sg13g2_decap_8 FILLER_164_1118 ();
 sg13g2_decap_8 FILLER_164_1125 ();
 sg13g2_decap_8 FILLER_164_1132 ();
 sg13g2_decap_8 FILLER_164_1139 ();
 sg13g2_decap_8 FILLER_164_1146 ();
 sg13g2_decap_4 FILLER_164_1153 ();
 sg13g2_decap_8 FILLER_164_1165 ();
 sg13g2_decap_8 FILLER_164_1172 ();
 sg13g2_decap_8 FILLER_164_1179 ();
 sg13g2_decap_8 FILLER_164_1186 ();
 sg13g2_decap_8 FILLER_164_1193 ();
 sg13g2_decap_8 FILLER_164_1200 ();
 sg13g2_decap_8 FILLER_164_1207 ();
 sg13g2_decap_4 FILLER_164_1214 ();
 sg13g2_fill_1 FILLER_164_1218 ();
 sg13g2_decap_8 FILLER_164_1224 ();
 sg13g2_decap_8 FILLER_164_1231 ();
 sg13g2_decap_4 FILLER_164_1238 ();
 sg13g2_fill_1 FILLER_164_1242 ();
 sg13g2_decap_8 FILLER_164_1261 ();
 sg13g2_decap_4 FILLER_164_1268 ();
 sg13g2_fill_2 FILLER_164_1272 ();
 sg13g2_decap_8 FILLER_164_1302 ();
 sg13g2_decap_8 FILLER_164_1309 ();
 sg13g2_decap_8 FILLER_164_1316 ();
 sg13g2_decap_8 FILLER_164_1323 ();
 sg13g2_decap_4 FILLER_164_1330 ();
 sg13g2_fill_2 FILLER_164_1334 ();
 sg13g2_fill_2 FILLER_164_1343 ();
 sg13g2_fill_1 FILLER_164_1345 ();
 sg13g2_decap_4 FILLER_164_1351 ();
 sg13g2_fill_1 FILLER_164_1355 ();
 sg13g2_fill_2 FILLER_164_1366 ();
 sg13g2_fill_1 FILLER_164_1376 ();
 sg13g2_fill_2 FILLER_164_1389 ();
 sg13g2_fill_1 FILLER_164_1391 ();
 sg13g2_decap_8 FILLER_164_1400 ();
 sg13g2_decap_8 FILLER_164_1407 ();
 sg13g2_decap_4 FILLER_164_1414 ();
 sg13g2_fill_2 FILLER_164_1418 ();
 sg13g2_fill_2 FILLER_164_1424 ();
 sg13g2_fill_1 FILLER_164_1426 ();
 sg13g2_decap_8 FILLER_164_1455 ();
 sg13g2_decap_4 FILLER_164_1462 ();
 sg13g2_fill_1 FILLER_164_1466 ();
 sg13g2_decap_8 FILLER_164_1494 ();
 sg13g2_decap_8 FILLER_164_1501 ();
 sg13g2_decap_8 FILLER_164_1508 ();
 sg13g2_decap_8 FILLER_164_1515 ();
 sg13g2_decap_8 FILLER_164_1522 ();
 sg13g2_decap_8 FILLER_164_1529 ();
 sg13g2_decap_8 FILLER_164_1536 ();
 sg13g2_decap_8 FILLER_164_1543 ();
 sg13g2_decap_8 FILLER_164_1550 ();
 sg13g2_decap_8 FILLER_164_1557 ();
 sg13g2_decap_8 FILLER_164_1564 ();
 sg13g2_decap_8 FILLER_164_1571 ();
 sg13g2_decap_8 FILLER_164_1578 ();
 sg13g2_decap_8 FILLER_164_1585 ();
 sg13g2_decap_8 FILLER_164_1592 ();
 sg13g2_decap_8 FILLER_164_1599 ();
 sg13g2_decap_8 FILLER_164_1606 ();
 sg13g2_decap_8 FILLER_164_1613 ();
 sg13g2_decap_8 FILLER_164_1620 ();
 sg13g2_decap_8 FILLER_164_1627 ();
 sg13g2_decap_8 FILLER_164_1634 ();
 sg13g2_decap_8 FILLER_164_1641 ();
 sg13g2_decap_8 FILLER_164_1648 ();
 sg13g2_decap_8 FILLER_164_1655 ();
 sg13g2_decap_8 FILLER_164_1662 ();
 sg13g2_decap_8 FILLER_164_1669 ();
 sg13g2_decap_8 FILLER_164_1676 ();
 sg13g2_decap_8 FILLER_164_1683 ();
 sg13g2_decap_8 FILLER_164_1690 ();
 sg13g2_decap_8 FILLER_164_1697 ();
 sg13g2_decap_8 FILLER_164_1704 ();
 sg13g2_decap_8 FILLER_164_1711 ();
 sg13g2_decap_8 FILLER_164_1718 ();
 sg13g2_decap_8 FILLER_164_1725 ();
 sg13g2_decap_8 FILLER_164_1732 ();
 sg13g2_decap_8 FILLER_164_1739 ();
 sg13g2_decap_8 FILLER_164_1746 ();
 sg13g2_decap_8 FILLER_164_1753 ();
 sg13g2_decap_8 FILLER_164_1760 ();
 sg13g2_fill_1 FILLER_164_1767 ();
 sg13g2_decap_8 FILLER_165_0 ();
 sg13g2_decap_8 FILLER_165_7 ();
 sg13g2_decap_8 FILLER_165_14 ();
 sg13g2_decap_8 FILLER_165_21 ();
 sg13g2_decap_8 FILLER_165_28 ();
 sg13g2_decap_8 FILLER_165_35 ();
 sg13g2_decap_8 FILLER_165_42 ();
 sg13g2_decap_8 FILLER_165_49 ();
 sg13g2_decap_8 FILLER_165_56 ();
 sg13g2_decap_8 FILLER_165_63 ();
 sg13g2_decap_8 FILLER_165_70 ();
 sg13g2_decap_8 FILLER_165_77 ();
 sg13g2_decap_8 FILLER_165_84 ();
 sg13g2_decap_8 FILLER_165_91 ();
 sg13g2_decap_8 FILLER_165_98 ();
 sg13g2_decap_8 FILLER_165_105 ();
 sg13g2_decap_8 FILLER_165_112 ();
 sg13g2_decap_8 FILLER_165_119 ();
 sg13g2_fill_2 FILLER_165_126 ();
 sg13g2_decap_4 FILLER_165_138 ();
 sg13g2_fill_2 FILLER_165_142 ();
 sg13g2_decap_8 FILLER_165_152 ();
 sg13g2_decap_8 FILLER_165_159 ();
 sg13g2_decap_8 FILLER_165_166 ();
 sg13g2_decap_8 FILLER_165_173 ();
 sg13g2_fill_1 FILLER_165_180 ();
 sg13g2_fill_2 FILLER_165_187 ();
 sg13g2_decap_8 FILLER_165_221 ();
 sg13g2_decap_8 FILLER_165_228 ();
 sg13g2_decap_4 FILLER_165_235 ();
 sg13g2_fill_2 FILLER_165_239 ();
 sg13g2_decap_8 FILLER_165_244 ();
 sg13g2_decap_8 FILLER_165_251 ();
 sg13g2_decap_8 FILLER_165_258 ();
 sg13g2_decap_8 FILLER_165_265 ();
 sg13g2_decap_8 FILLER_165_272 ();
 sg13g2_decap_8 FILLER_165_279 ();
 sg13g2_decap_4 FILLER_165_286 ();
 sg13g2_fill_1 FILLER_165_290 ();
 sg13g2_decap_8 FILLER_165_296 ();
 sg13g2_decap_8 FILLER_165_303 ();
 sg13g2_fill_2 FILLER_165_315 ();
 sg13g2_fill_1 FILLER_165_322 ();
 sg13g2_decap_8 FILLER_165_331 ();
 sg13g2_decap_8 FILLER_165_338 ();
 sg13g2_fill_2 FILLER_165_345 ();
 sg13g2_decap_8 FILLER_165_355 ();
 sg13g2_decap_8 FILLER_165_362 ();
 sg13g2_decap_8 FILLER_165_369 ();
 sg13g2_decap_8 FILLER_165_376 ();
 sg13g2_decap_8 FILLER_165_383 ();
 sg13g2_decap_4 FILLER_165_390 ();
 sg13g2_decap_8 FILLER_165_420 ();
 sg13g2_decap_8 FILLER_165_427 ();
 sg13g2_decap_8 FILLER_165_434 ();
 sg13g2_decap_8 FILLER_165_441 ();
 sg13g2_decap_8 FILLER_165_448 ();
 sg13g2_decap_8 FILLER_165_455 ();
 sg13g2_decap_8 FILLER_165_462 ();
 sg13g2_fill_2 FILLER_165_469 ();
 sg13g2_fill_1 FILLER_165_471 ();
 sg13g2_decap_8 FILLER_165_477 ();
 sg13g2_decap_8 FILLER_165_484 ();
 sg13g2_decap_8 FILLER_165_491 ();
 sg13g2_decap_8 FILLER_165_498 ();
 sg13g2_decap_8 FILLER_165_505 ();
 sg13g2_decap_4 FILLER_165_512 ();
 sg13g2_decap_8 FILLER_165_519 ();
 sg13g2_decap_8 FILLER_165_526 ();
 sg13g2_decap_8 FILLER_165_533 ();
 sg13g2_fill_1 FILLER_165_540 ();
 sg13g2_decap_8 FILLER_165_549 ();
 sg13g2_decap_8 FILLER_165_556 ();
 sg13g2_decap_8 FILLER_165_563 ();
 sg13g2_decap_8 FILLER_165_570 ();
 sg13g2_decap_8 FILLER_165_577 ();
 sg13g2_decap_8 FILLER_165_584 ();
 sg13g2_fill_2 FILLER_165_591 ();
 sg13g2_fill_1 FILLER_165_593 ();
 sg13g2_fill_2 FILLER_165_602 ();
 sg13g2_decap_8 FILLER_165_609 ();
 sg13g2_decap_8 FILLER_165_616 ();
 sg13g2_decap_8 FILLER_165_623 ();
 sg13g2_decap_8 FILLER_165_630 ();
 sg13g2_decap_8 FILLER_165_637 ();
 sg13g2_decap_8 FILLER_165_644 ();
 sg13g2_decap_8 FILLER_165_651 ();
 sg13g2_fill_1 FILLER_165_658 ();
 sg13g2_fill_1 FILLER_165_695 ();
 sg13g2_decap_8 FILLER_165_705 ();
 sg13g2_decap_8 FILLER_165_712 ();
 sg13g2_decap_8 FILLER_165_719 ();
 sg13g2_decap_8 FILLER_165_726 ();
 sg13g2_decap_4 FILLER_165_733 ();
 sg13g2_fill_2 FILLER_165_737 ();
 sg13g2_decap_8 FILLER_165_742 ();
 sg13g2_decap_8 FILLER_165_749 ();
 sg13g2_decap_8 FILLER_165_756 ();
 sg13g2_decap_8 FILLER_165_763 ();
 sg13g2_decap_8 FILLER_165_770 ();
 sg13g2_decap_8 FILLER_165_777 ();
 sg13g2_decap_4 FILLER_165_784 ();
 sg13g2_decap_8 FILLER_165_792 ();
 sg13g2_decap_8 FILLER_165_799 ();
 sg13g2_decap_8 FILLER_165_806 ();
 sg13g2_decap_4 FILLER_165_813 ();
 sg13g2_fill_2 FILLER_165_817 ();
 sg13g2_decap_8 FILLER_165_832 ();
 sg13g2_decap_8 FILLER_165_839 ();
 sg13g2_decap_8 FILLER_165_846 ();
 sg13g2_decap_8 FILLER_165_853 ();
 sg13g2_decap_8 FILLER_165_860 ();
 sg13g2_decap_8 FILLER_165_875 ();
 sg13g2_fill_1 FILLER_165_882 ();
 sg13g2_decap_8 FILLER_165_888 ();
 sg13g2_decap_8 FILLER_165_895 ();
 sg13g2_decap_8 FILLER_165_902 ();
 sg13g2_decap_8 FILLER_165_909 ();
 sg13g2_fill_2 FILLER_165_916 ();
 sg13g2_decap_8 FILLER_165_934 ();
 sg13g2_decap_8 FILLER_165_941 ();
 sg13g2_decap_8 FILLER_165_948 ();
 sg13g2_decap_8 FILLER_165_955 ();
 sg13g2_decap_4 FILLER_165_962 ();
 sg13g2_decap_8 FILLER_165_977 ();
 sg13g2_decap_8 FILLER_165_984 ();
 sg13g2_decap_8 FILLER_165_991 ();
 sg13g2_decap_8 FILLER_165_998 ();
 sg13g2_decap_8 FILLER_165_1005 ();
 sg13g2_decap_8 FILLER_165_1012 ();
 sg13g2_decap_8 FILLER_165_1019 ();
 sg13g2_decap_8 FILLER_165_1026 ();
 sg13g2_decap_4 FILLER_165_1033 ();
 sg13g2_fill_2 FILLER_165_1041 ();
 sg13g2_decap_8 FILLER_165_1051 ();
 sg13g2_decap_8 FILLER_165_1058 ();
 sg13g2_decap_8 FILLER_165_1065 ();
 sg13g2_fill_2 FILLER_165_1072 ();
 sg13g2_fill_1 FILLER_165_1074 ();
 sg13g2_decap_8 FILLER_165_1079 ();
 sg13g2_decap_8 FILLER_165_1086 ();
 sg13g2_decap_8 FILLER_165_1093 ();
 sg13g2_decap_8 FILLER_165_1100 ();
 sg13g2_decap_8 FILLER_165_1107 ();
 sg13g2_decap_8 FILLER_165_1114 ();
 sg13g2_decap_8 FILLER_165_1121 ();
 sg13g2_decap_8 FILLER_165_1128 ();
 sg13g2_decap_8 FILLER_165_1135 ();
 sg13g2_fill_2 FILLER_165_1142 ();
 sg13g2_decap_8 FILLER_165_1170 ();
 sg13g2_decap_8 FILLER_165_1177 ();
 sg13g2_decap_8 FILLER_165_1184 ();
 sg13g2_decap_8 FILLER_165_1191 ();
 sg13g2_decap_8 FILLER_165_1198 ();
 sg13g2_fill_2 FILLER_165_1205 ();
 sg13g2_fill_1 FILLER_165_1207 ();
 sg13g2_fill_2 FILLER_165_1233 ();
 sg13g2_decap_8 FILLER_165_1250 ();
 sg13g2_decap_8 FILLER_165_1257 ();
 sg13g2_decap_8 FILLER_165_1264 ();
 sg13g2_decap_8 FILLER_165_1271 ();
 sg13g2_decap_4 FILLER_165_1278 ();
 sg13g2_fill_1 FILLER_165_1282 ();
 sg13g2_decap_8 FILLER_165_1288 ();
 sg13g2_decap_8 FILLER_165_1295 ();
 sg13g2_decap_8 FILLER_165_1302 ();
 sg13g2_decap_8 FILLER_165_1309 ();
 sg13g2_decap_8 FILLER_165_1316 ();
 sg13g2_fill_2 FILLER_165_1323 ();
 sg13g2_fill_1 FILLER_165_1325 ();
 sg13g2_decap_8 FILLER_165_1398 ();
 sg13g2_decap_8 FILLER_165_1405 ();
 sg13g2_fill_2 FILLER_165_1412 ();
 sg13g2_fill_1 FILLER_165_1414 ();
 sg13g2_decap_4 FILLER_165_1439 ();
 sg13g2_fill_1 FILLER_165_1443 ();
 sg13g2_decap_8 FILLER_165_1448 ();
 sg13g2_decap_8 FILLER_165_1455 ();
 sg13g2_decap_8 FILLER_165_1462 ();
 sg13g2_decap_4 FILLER_165_1469 ();
 sg13g2_fill_1 FILLER_165_1473 ();
 sg13g2_decap_8 FILLER_165_1484 ();
 sg13g2_decap_8 FILLER_165_1491 ();
 sg13g2_decap_8 FILLER_165_1498 ();
 sg13g2_decap_8 FILLER_165_1505 ();
 sg13g2_decap_8 FILLER_165_1512 ();
 sg13g2_decap_8 FILLER_165_1519 ();
 sg13g2_decap_8 FILLER_165_1526 ();
 sg13g2_decap_8 FILLER_165_1533 ();
 sg13g2_decap_8 FILLER_165_1540 ();
 sg13g2_decap_8 FILLER_165_1547 ();
 sg13g2_decap_8 FILLER_165_1554 ();
 sg13g2_decap_8 FILLER_165_1561 ();
 sg13g2_decap_8 FILLER_165_1568 ();
 sg13g2_decap_8 FILLER_165_1575 ();
 sg13g2_decap_8 FILLER_165_1582 ();
 sg13g2_decap_8 FILLER_165_1589 ();
 sg13g2_decap_8 FILLER_165_1596 ();
 sg13g2_decap_8 FILLER_165_1603 ();
 sg13g2_decap_8 FILLER_165_1610 ();
 sg13g2_decap_8 FILLER_165_1617 ();
 sg13g2_decap_8 FILLER_165_1624 ();
 sg13g2_decap_8 FILLER_165_1631 ();
 sg13g2_decap_8 FILLER_165_1638 ();
 sg13g2_decap_8 FILLER_165_1645 ();
 sg13g2_decap_8 FILLER_165_1652 ();
 sg13g2_decap_8 FILLER_165_1659 ();
 sg13g2_decap_8 FILLER_165_1666 ();
 sg13g2_decap_8 FILLER_165_1673 ();
 sg13g2_decap_8 FILLER_165_1680 ();
 sg13g2_decap_8 FILLER_165_1687 ();
 sg13g2_decap_8 FILLER_165_1694 ();
 sg13g2_decap_8 FILLER_165_1701 ();
 sg13g2_decap_8 FILLER_165_1708 ();
 sg13g2_decap_8 FILLER_165_1715 ();
 sg13g2_decap_8 FILLER_165_1722 ();
 sg13g2_decap_8 FILLER_165_1729 ();
 sg13g2_decap_8 FILLER_165_1736 ();
 sg13g2_decap_8 FILLER_165_1743 ();
 sg13g2_decap_8 FILLER_165_1750 ();
 sg13g2_decap_8 FILLER_165_1757 ();
 sg13g2_decap_4 FILLER_165_1764 ();
 sg13g2_decap_8 FILLER_166_0 ();
 sg13g2_decap_8 FILLER_166_7 ();
 sg13g2_decap_8 FILLER_166_14 ();
 sg13g2_decap_8 FILLER_166_21 ();
 sg13g2_decap_8 FILLER_166_28 ();
 sg13g2_decap_8 FILLER_166_35 ();
 sg13g2_decap_8 FILLER_166_42 ();
 sg13g2_decap_8 FILLER_166_49 ();
 sg13g2_decap_8 FILLER_166_56 ();
 sg13g2_decap_8 FILLER_166_63 ();
 sg13g2_decap_8 FILLER_166_70 ();
 sg13g2_decap_8 FILLER_166_77 ();
 sg13g2_decap_8 FILLER_166_84 ();
 sg13g2_decap_8 FILLER_166_91 ();
 sg13g2_decap_8 FILLER_166_98 ();
 sg13g2_decap_8 FILLER_166_105 ();
 sg13g2_decap_8 FILLER_166_112 ();
 sg13g2_decap_8 FILLER_166_119 ();
 sg13g2_decap_8 FILLER_166_126 ();
 sg13g2_decap_8 FILLER_166_133 ();
 sg13g2_decap_8 FILLER_166_140 ();
 sg13g2_decap_8 FILLER_166_147 ();
 sg13g2_decap_8 FILLER_166_154 ();
 sg13g2_decap_8 FILLER_166_161 ();
 sg13g2_decap_4 FILLER_166_168 ();
 sg13g2_fill_1 FILLER_166_172 ();
 sg13g2_fill_1 FILLER_166_205 ();
 sg13g2_decap_8 FILLER_166_209 ();
 sg13g2_decap_8 FILLER_166_216 ();
 sg13g2_decap_8 FILLER_166_223 ();
 sg13g2_decap_8 FILLER_166_230 ();
 sg13g2_decap_8 FILLER_166_237 ();
 sg13g2_decap_8 FILLER_166_244 ();
 sg13g2_decap_8 FILLER_166_251 ();
 sg13g2_decap_8 FILLER_166_258 ();
 sg13g2_decap_8 FILLER_166_265 ();
 sg13g2_decap_8 FILLER_166_272 ();
 sg13g2_decap_4 FILLER_166_279 ();
 sg13g2_fill_2 FILLER_166_283 ();
 sg13g2_fill_2 FILLER_166_300 ();
 sg13g2_fill_1 FILLER_166_302 ();
 sg13g2_decap_8 FILLER_166_332 ();
 sg13g2_decap_8 FILLER_166_339 ();
 sg13g2_decap_8 FILLER_166_346 ();
 sg13g2_decap_4 FILLER_166_353 ();
 sg13g2_decap_8 FILLER_166_363 ();
 sg13g2_decap_8 FILLER_166_370 ();
 sg13g2_decap_8 FILLER_166_377 ();
 sg13g2_decap_8 FILLER_166_384 ();
 sg13g2_decap_8 FILLER_166_391 ();
 sg13g2_decap_8 FILLER_166_398 ();
 sg13g2_decap_8 FILLER_166_405 ();
 sg13g2_decap_8 FILLER_166_412 ();
 sg13g2_decap_8 FILLER_166_419 ();
 sg13g2_decap_8 FILLER_166_426 ();
 sg13g2_decap_8 FILLER_166_433 ();
 sg13g2_decap_4 FILLER_166_440 ();
 sg13g2_fill_1 FILLER_166_460 ();
 sg13g2_decap_8 FILLER_166_473 ();
 sg13g2_decap_8 FILLER_166_480 ();
 sg13g2_decap_4 FILLER_166_487 ();
 sg13g2_fill_2 FILLER_166_491 ();
 sg13g2_decap_8 FILLER_166_505 ();
 sg13g2_decap_8 FILLER_166_520 ();
 sg13g2_decap_8 FILLER_166_532 ();
 sg13g2_decap_8 FILLER_166_539 ();
 sg13g2_decap_8 FILLER_166_546 ();
 sg13g2_decap_8 FILLER_166_553 ();
 sg13g2_decap_8 FILLER_166_560 ();
 sg13g2_decap_8 FILLER_166_567 ();
 sg13g2_decap_8 FILLER_166_574 ();
 sg13g2_decap_4 FILLER_166_581 ();
 sg13g2_fill_2 FILLER_166_585 ();
 sg13g2_fill_2 FILLER_166_600 ();
 sg13g2_decap_8 FILLER_166_620 ();
 sg13g2_decap_8 FILLER_166_627 ();
 sg13g2_decap_8 FILLER_166_634 ();
 sg13g2_decap_8 FILLER_166_641 ();
 sg13g2_decap_8 FILLER_166_648 ();
 sg13g2_decap_8 FILLER_166_655 ();
 sg13g2_decap_8 FILLER_166_662 ();
 sg13g2_decap_8 FILLER_166_669 ();
 sg13g2_decap_4 FILLER_166_676 ();
 sg13g2_decap_8 FILLER_166_684 ();
 sg13g2_decap_8 FILLER_166_691 ();
 sg13g2_decap_8 FILLER_166_698 ();
 sg13g2_fill_1 FILLER_166_705 ();
 sg13g2_decap_8 FILLER_166_716 ();
 sg13g2_decap_8 FILLER_166_723 ();
 sg13g2_decap_4 FILLER_166_730 ();
 sg13g2_fill_1 FILLER_166_734 ();
 sg13g2_decap_4 FILLER_166_739 ();
 sg13g2_fill_2 FILLER_166_743 ();
 sg13g2_decap_8 FILLER_166_753 ();
 sg13g2_decap_8 FILLER_166_760 ();
 sg13g2_decap_8 FILLER_166_767 ();
 sg13g2_decap_8 FILLER_166_774 ();
 sg13g2_fill_1 FILLER_166_781 ();
 sg13g2_decap_8 FILLER_166_802 ();
 sg13g2_decap_8 FILLER_166_809 ();
 sg13g2_decap_4 FILLER_166_816 ();
 sg13g2_fill_2 FILLER_166_820 ();
 sg13g2_decap_8 FILLER_166_827 ();
 sg13g2_decap_8 FILLER_166_834 ();
 sg13g2_decap_8 FILLER_166_841 ();
 sg13g2_decap_4 FILLER_166_848 ();
 sg13g2_decap_8 FILLER_166_855 ();
 sg13g2_decap_8 FILLER_166_862 ();
 sg13g2_decap_8 FILLER_166_869 ();
 sg13g2_decap_4 FILLER_166_876 ();
 sg13g2_fill_1 FILLER_166_880 ();
 sg13g2_decap_8 FILLER_166_894 ();
 sg13g2_decap_8 FILLER_166_901 ();
 sg13g2_decap_8 FILLER_166_908 ();
 sg13g2_decap_8 FILLER_166_915 ();
 sg13g2_decap_8 FILLER_166_922 ();
 sg13g2_decap_8 FILLER_166_929 ();
 sg13g2_decap_8 FILLER_166_936 ();
 sg13g2_decap_8 FILLER_166_943 ();
 sg13g2_decap_8 FILLER_166_950 ();
 sg13g2_fill_2 FILLER_166_957 ();
 sg13g2_decap_8 FILLER_166_984 ();
 sg13g2_decap_8 FILLER_166_991 ();
 sg13g2_decap_4 FILLER_166_998 ();
 sg13g2_decap_8 FILLER_166_1006 ();
 sg13g2_decap_8 FILLER_166_1034 ();
 sg13g2_decap_8 FILLER_166_1041 ();
 sg13g2_decap_8 FILLER_166_1048 ();
 sg13g2_decap_8 FILLER_166_1055 ();
 sg13g2_decap_8 FILLER_166_1062 ();
 sg13g2_fill_1 FILLER_166_1069 ();
 sg13g2_decap_8 FILLER_166_1079 ();
 sg13g2_decap_8 FILLER_166_1086 ();
 sg13g2_decap_8 FILLER_166_1093 ();
 sg13g2_decap_8 FILLER_166_1100 ();
 sg13g2_decap_8 FILLER_166_1107 ();
 sg13g2_decap_8 FILLER_166_1114 ();
 sg13g2_decap_8 FILLER_166_1121 ();
 sg13g2_decap_4 FILLER_166_1128 ();
 sg13g2_fill_1 FILLER_166_1132 ();
 sg13g2_fill_1 FILLER_166_1141 ();
 sg13g2_decap_8 FILLER_166_1176 ();
 sg13g2_decap_8 FILLER_166_1183 ();
 sg13g2_decap_8 FILLER_166_1190 ();
 sg13g2_decap_8 FILLER_166_1197 ();
 sg13g2_decap_4 FILLER_166_1204 ();
 sg13g2_fill_1 FILLER_166_1208 ();
 sg13g2_decap_8 FILLER_166_1225 ();
 sg13g2_fill_1 FILLER_166_1232 ();
 sg13g2_decap_8 FILLER_166_1238 ();
 sg13g2_decap_8 FILLER_166_1245 ();
 sg13g2_decap_4 FILLER_166_1252 ();
 sg13g2_fill_2 FILLER_166_1256 ();
 sg13g2_decap_8 FILLER_166_1262 ();
 sg13g2_decap_8 FILLER_166_1269 ();
 sg13g2_decap_8 FILLER_166_1276 ();
 sg13g2_decap_8 FILLER_166_1283 ();
 sg13g2_decap_8 FILLER_166_1290 ();
 sg13g2_decap_8 FILLER_166_1297 ();
 sg13g2_decap_8 FILLER_166_1304 ();
 sg13g2_decap_8 FILLER_166_1311 ();
 sg13g2_decap_8 FILLER_166_1318 ();
 sg13g2_decap_8 FILLER_166_1325 ();
 sg13g2_fill_1 FILLER_166_1332 ();
 sg13g2_decap_8 FILLER_166_1338 ();
 sg13g2_decap_8 FILLER_166_1345 ();
 sg13g2_decap_8 FILLER_166_1352 ();
 sg13g2_fill_2 FILLER_166_1382 ();
 sg13g2_decap_8 FILLER_166_1389 ();
 sg13g2_decap_8 FILLER_166_1396 ();
 sg13g2_decap_4 FILLER_166_1403 ();
 sg13g2_fill_2 FILLER_166_1407 ();
 sg13g2_decap_4 FILLER_166_1423 ();
 sg13g2_decap_8 FILLER_166_1438 ();
 sg13g2_decap_8 FILLER_166_1445 ();
 sg13g2_decap_8 FILLER_166_1452 ();
 sg13g2_decap_8 FILLER_166_1459 ();
 sg13g2_decap_8 FILLER_166_1466 ();
 sg13g2_decap_8 FILLER_166_1473 ();
 sg13g2_decap_8 FILLER_166_1480 ();
 sg13g2_decap_8 FILLER_166_1487 ();
 sg13g2_decap_8 FILLER_166_1494 ();
 sg13g2_decap_8 FILLER_166_1501 ();
 sg13g2_decap_8 FILLER_166_1508 ();
 sg13g2_decap_8 FILLER_166_1515 ();
 sg13g2_decap_8 FILLER_166_1522 ();
 sg13g2_decap_8 FILLER_166_1529 ();
 sg13g2_decap_8 FILLER_166_1536 ();
 sg13g2_decap_8 FILLER_166_1543 ();
 sg13g2_decap_8 FILLER_166_1550 ();
 sg13g2_decap_8 FILLER_166_1557 ();
 sg13g2_decap_8 FILLER_166_1564 ();
 sg13g2_decap_8 FILLER_166_1571 ();
 sg13g2_decap_8 FILLER_166_1578 ();
 sg13g2_decap_8 FILLER_166_1585 ();
 sg13g2_decap_8 FILLER_166_1592 ();
 sg13g2_decap_8 FILLER_166_1599 ();
 sg13g2_decap_8 FILLER_166_1606 ();
 sg13g2_decap_8 FILLER_166_1613 ();
 sg13g2_decap_8 FILLER_166_1620 ();
 sg13g2_decap_8 FILLER_166_1627 ();
 sg13g2_decap_8 FILLER_166_1634 ();
 sg13g2_decap_8 FILLER_166_1641 ();
 sg13g2_decap_8 FILLER_166_1648 ();
 sg13g2_decap_8 FILLER_166_1655 ();
 sg13g2_decap_8 FILLER_166_1662 ();
 sg13g2_decap_8 FILLER_166_1669 ();
 sg13g2_decap_8 FILLER_166_1676 ();
 sg13g2_decap_8 FILLER_166_1683 ();
 sg13g2_decap_8 FILLER_166_1690 ();
 sg13g2_decap_8 FILLER_166_1697 ();
 sg13g2_decap_8 FILLER_166_1704 ();
 sg13g2_decap_8 FILLER_166_1711 ();
 sg13g2_decap_8 FILLER_166_1718 ();
 sg13g2_decap_8 FILLER_166_1725 ();
 sg13g2_decap_8 FILLER_166_1732 ();
 sg13g2_decap_8 FILLER_166_1739 ();
 sg13g2_decap_8 FILLER_166_1746 ();
 sg13g2_decap_8 FILLER_166_1753 ();
 sg13g2_decap_8 FILLER_166_1760 ();
 sg13g2_fill_1 FILLER_166_1767 ();
 sg13g2_decap_8 FILLER_167_0 ();
 sg13g2_decap_8 FILLER_167_7 ();
 sg13g2_decap_8 FILLER_167_14 ();
 sg13g2_decap_8 FILLER_167_21 ();
 sg13g2_decap_8 FILLER_167_28 ();
 sg13g2_decap_8 FILLER_167_35 ();
 sg13g2_decap_8 FILLER_167_42 ();
 sg13g2_decap_8 FILLER_167_49 ();
 sg13g2_decap_8 FILLER_167_56 ();
 sg13g2_decap_8 FILLER_167_63 ();
 sg13g2_decap_8 FILLER_167_70 ();
 sg13g2_decap_8 FILLER_167_77 ();
 sg13g2_decap_8 FILLER_167_84 ();
 sg13g2_decap_8 FILLER_167_91 ();
 sg13g2_decap_8 FILLER_167_98 ();
 sg13g2_decap_8 FILLER_167_105 ();
 sg13g2_decap_8 FILLER_167_112 ();
 sg13g2_decap_8 FILLER_167_119 ();
 sg13g2_decap_8 FILLER_167_126 ();
 sg13g2_decap_8 FILLER_167_133 ();
 sg13g2_decap_8 FILLER_167_140 ();
 sg13g2_decap_8 FILLER_167_147 ();
 sg13g2_decap_8 FILLER_167_154 ();
 sg13g2_decap_8 FILLER_167_161 ();
 sg13g2_decap_8 FILLER_167_168 ();
 sg13g2_decap_8 FILLER_167_175 ();
 sg13g2_decap_8 FILLER_167_199 ();
 sg13g2_decap_8 FILLER_167_206 ();
 sg13g2_decap_8 FILLER_167_213 ();
 sg13g2_decap_8 FILLER_167_220 ();
 sg13g2_decap_8 FILLER_167_227 ();
 sg13g2_decap_8 FILLER_167_234 ();
 sg13g2_fill_2 FILLER_167_241 ();
 sg13g2_decap_8 FILLER_167_267 ();
 sg13g2_fill_2 FILLER_167_274 ();
 sg13g2_fill_2 FILLER_167_281 ();
 sg13g2_fill_1 FILLER_167_283 ();
 sg13g2_decap_8 FILLER_167_299 ();
 sg13g2_fill_2 FILLER_167_306 ();
 sg13g2_fill_1 FILLER_167_312 ();
 sg13g2_decap_4 FILLER_167_323 ();
 sg13g2_fill_2 FILLER_167_334 ();
 sg13g2_decap_8 FILLER_167_340 ();
 sg13g2_decap_4 FILLER_167_347 ();
 sg13g2_fill_1 FILLER_167_351 ();
 sg13g2_decap_8 FILLER_167_375 ();
 sg13g2_decap_8 FILLER_167_382 ();
 sg13g2_decap_8 FILLER_167_389 ();
 sg13g2_decap_8 FILLER_167_396 ();
 sg13g2_fill_2 FILLER_167_403 ();
 sg13g2_fill_1 FILLER_167_405 ();
 sg13g2_decap_8 FILLER_167_410 ();
 sg13g2_fill_1 FILLER_167_417 ();
 sg13g2_decap_8 FILLER_167_422 ();
 sg13g2_decap_8 FILLER_167_429 ();
 sg13g2_decap_4 FILLER_167_436 ();
 sg13g2_fill_2 FILLER_167_440 ();
 sg13g2_decap_8 FILLER_167_447 ();
 sg13g2_fill_2 FILLER_167_454 ();
 sg13g2_fill_1 FILLER_167_456 ();
 sg13g2_decap_8 FILLER_167_465 ();
 sg13g2_decap_8 FILLER_167_472 ();
 sg13g2_decap_8 FILLER_167_479 ();
 sg13g2_decap_8 FILLER_167_486 ();
 sg13g2_decap_4 FILLER_167_493 ();
 sg13g2_fill_2 FILLER_167_497 ();
 sg13g2_fill_1 FILLER_167_507 ();
 sg13g2_fill_2 FILLER_167_520 ();
 sg13g2_decap_8 FILLER_167_541 ();
 sg13g2_decap_8 FILLER_167_548 ();
 sg13g2_decap_8 FILLER_167_555 ();
 sg13g2_fill_2 FILLER_167_562 ();
 sg13g2_fill_1 FILLER_167_564 ();
 sg13g2_decap_8 FILLER_167_574 ();
 sg13g2_decap_4 FILLER_167_581 ();
 sg13g2_fill_1 FILLER_167_585 ();
 sg13g2_fill_2 FILLER_167_594 ();
 sg13g2_fill_1 FILLER_167_596 ();
 sg13g2_decap_8 FILLER_167_608 ();
 sg13g2_decap_8 FILLER_167_615 ();
 sg13g2_decap_8 FILLER_167_622 ();
 sg13g2_decap_8 FILLER_167_629 ();
 sg13g2_decap_8 FILLER_167_636 ();
 sg13g2_decap_8 FILLER_167_643 ();
 sg13g2_fill_2 FILLER_167_650 ();
 sg13g2_decap_8 FILLER_167_662 ();
 sg13g2_decap_8 FILLER_167_669 ();
 sg13g2_decap_8 FILLER_167_676 ();
 sg13g2_decap_8 FILLER_167_683 ();
 sg13g2_decap_8 FILLER_167_690 ();
 sg13g2_decap_8 FILLER_167_697 ();
 sg13g2_decap_8 FILLER_167_704 ();
 sg13g2_decap_4 FILLER_167_711 ();
 sg13g2_decap_4 FILLER_167_719 ();
 sg13g2_fill_1 FILLER_167_723 ();
 sg13g2_decap_8 FILLER_167_750 ();
 sg13g2_decap_8 FILLER_167_757 ();
 sg13g2_decap_8 FILLER_167_764 ();
 sg13g2_decap_8 FILLER_167_771 ();
 sg13g2_fill_1 FILLER_167_778 ();
 sg13g2_fill_1 FILLER_167_787 ();
 sg13g2_decap_8 FILLER_167_792 ();
 sg13g2_decap_8 FILLER_167_799 ();
 sg13g2_decap_8 FILLER_167_806 ();
 sg13g2_decap_8 FILLER_167_813 ();
 sg13g2_decap_8 FILLER_167_820 ();
 sg13g2_decap_8 FILLER_167_827 ();
 sg13g2_decap_8 FILLER_167_837 ();
 sg13g2_decap_8 FILLER_167_844 ();
 sg13g2_fill_2 FILLER_167_851 ();
 sg13g2_decap_8 FILLER_167_858 ();
 sg13g2_decap_8 FILLER_167_865 ();
 sg13g2_decap_8 FILLER_167_872 ();
 sg13g2_decap_8 FILLER_167_879 ();
 sg13g2_decap_8 FILLER_167_886 ();
 sg13g2_decap_8 FILLER_167_893 ();
 sg13g2_decap_4 FILLER_167_900 ();
 sg13g2_fill_1 FILLER_167_904 ();
 sg13g2_decap_8 FILLER_167_910 ();
 sg13g2_decap_8 FILLER_167_917 ();
 sg13g2_decap_8 FILLER_167_924 ();
 sg13g2_decap_8 FILLER_167_931 ();
 sg13g2_decap_8 FILLER_167_938 ();
 sg13g2_decap_8 FILLER_167_945 ();
 sg13g2_decap_8 FILLER_167_952 ();
 sg13g2_decap_4 FILLER_167_959 ();
 sg13g2_decap_8 FILLER_167_982 ();
 sg13g2_decap_8 FILLER_167_989 ();
 sg13g2_fill_1 FILLER_167_996 ();
 sg13g2_fill_2 FILLER_167_1009 ();
 sg13g2_decap_8 FILLER_167_1027 ();
 sg13g2_decap_8 FILLER_167_1034 ();
 sg13g2_decap_8 FILLER_167_1041 ();
 sg13g2_decap_8 FILLER_167_1048 ();
 sg13g2_decap_8 FILLER_167_1055 ();
 sg13g2_decap_8 FILLER_167_1062 ();
 sg13g2_fill_1 FILLER_167_1077 ();
 sg13g2_decap_8 FILLER_167_1083 ();
 sg13g2_decap_8 FILLER_167_1090 ();
 sg13g2_decap_8 FILLER_167_1097 ();
 sg13g2_decap_8 FILLER_167_1104 ();
 sg13g2_decap_8 FILLER_167_1111 ();
 sg13g2_decap_8 FILLER_167_1118 ();
 sg13g2_decap_8 FILLER_167_1125 ();
 sg13g2_decap_8 FILLER_167_1132 ();
 sg13g2_decap_8 FILLER_167_1139 ();
 sg13g2_fill_2 FILLER_167_1150 ();
 sg13g2_fill_2 FILLER_167_1161 ();
 sg13g2_fill_1 FILLER_167_1163 ();
 sg13g2_decap_8 FILLER_167_1179 ();
 sg13g2_decap_8 FILLER_167_1186 ();
 sg13g2_decap_4 FILLER_167_1193 ();
 sg13g2_fill_1 FILLER_167_1197 ();
 sg13g2_fill_2 FILLER_167_1203 ();
 sg13g2_fill_1 FILLER_167_1205 ();
 sg13g2_decap_8 FILLER_167_1210 ();
 sg13g2_decap_8 FILLER_167_1217 ();
 sg13g2_fill_2 FILLER_167_1224 ();
 sg13g2_decap_8 FILLER_167_1243 ();
 sg13g2_fill_2 FILLER_167_1250 ();
 sg13g2_fill_1 FILLER_167_1252 ();
 sg13g2_decap_8 FILLER_167_1273 ();
 sg13g2_decap_8 FILLER_167_1280 ();
 sg13g2_decap_8 FILLER_167_1287 ();
 sg13g2_decap_8 FILLER_167_1294 ();
 sg13g2_decap_8 FILLER_167_1301 ();
 sg13g2_decap_8 FILLER_167_1308 ();
 sg13g2_decap_8 FILLER_167_1315 ();
 sg13g2_decap_8 FILLER_167_1322 ();
 sg13g2_decap_8 FILLER_167_1329 ();
 sg13g2_decap_8 FILLER_167_1336 ();
 sg13g2_decap_8 FILLER_167_1343 ();
 sg13g2_decap_8 FILLER_167_1350 ();
 sg13g2_decap_8 FILLER_167_1357 ();
 sg13g2_decap_8 FILLER_167_1364 ();
 sg13g2_decap_8 FILLER_167_1371 ();
 sg13g2_decap_8 FILLER_167_1378 ();
 sg13g2_decap_8 FILLER_167_1385 ();
 sg13g2_decap_8 FILLER_167_1392 ();
 sg13g2_decap_8 FILLER_167_1399 ();
 sg13g2_decap_8 FILLER_167_1406 ();
 sg13g2_decap_4 FILLER_167_1413 ();
 sg13g2_fill_2 FILLER_167_1417 ();
 sg13g2_decap_8 FILLER_167_1424 ();
 sg13g2_decap_8 FILLER_167_1431 ();
 sg13g2_decap_8 FILLER_167_1438 ();
 sg13g2_decap_8 FILLER_167_1445 ();
 sg13g2_decap_8 FILLER_167_1452 ();
 sg13g2_decap_8 FILLER_167_1459 ();
 sg13g2_decap_8 FILLER_167_1466 ();
 sg13g2_decap_8 FILLER_167_1473 ();
 sg13g2_decap_8 FILLER_167_1480 ();
 sg13g2_decap_8 FILLER_167_1487 ();
 sg13g2_decap_8 FILLER_167_1494 ();
 sg13g2_decap_8 FILLER_167_1501 ();
 sg13g2_decap_8 FILLER_167_1508 ();
 sg13g2_decap_8 FILLER_167_1515 ();
 sg13g2_decap_8 FILLER_167_1522 ();
 sg13g2_decap_8 FILLER_167_1529 ();
 sg13g2_decap_8 FILLER_167_1536 ();
 sg13g2_decap_8 FILLER_167_1543 ();
 sg13g2_decap_8 FILLER_167_1550 ();
 sg13g2_decap_8 FILLER_167_1557 ();
 sg13g2_decap_8 FILLER_167_1564 ();
 sg13g2_decap_8 FILLER_167_1571 ();
 sg13g2_decap_8 FILLER_167_1578 ();
 sg13g2_decap_8 FILLER_167_1585 ();
 sg13g2_decap_8 FILLER_167_1592 ();
 sg13g2_decap_8 FILLER_167_1599 ();
 sg13g2_decap_8 FILLER_167_1606 ();
 sg13g2_decap_8 FILLER_167_1613 ();
 sg13g2_decap_8 FILLER_167_1620 ();
 sg13g2_decap_8 FILLER_167_1627 ();
 sg13g2_decap_8 FILLER_167_1634 ();
 sg13g2_decap_8 FILLER_167_1641 ();
 sg13g2_decap_8 FILLER_167_1648 ();
 sg13g2_decap_8 FILLER_167_1655 ();
 sg13g2_decap_8 FILLER_167_1662 ();
 sg13g2_decap_8 FILLER_167_1669 ();
 sg13g2_decap_8 FILLER_167_1676 ();
 sg13g2_decap_8 FILLER_167_1683 ();
 sg13g2_decap_8 FILLER_167_1690 ();
 sg13g2_decap_8 FILLER_167_1697 ();
 sg13g2_decap_8 FILLER_167_1704 ();
 sg13g2_decap_8 FILLER_167_1711 ();
 sg13g2_decap_8 FILLER_167_1718 ();
 sg13g2_decap_8 FILLER_167_1725 ();
 sg13g2_decap_8 FILLER_167_1732 ();
 sg13g2_decap_8 FILLER_167_1739 ();
 sg13g2_decap_8 FILLER_167_1746 ();
 sg13g2_decap_8 FILLER_167_1753 ();
 sg13g2_decap_8 FILLER_167_1760 ();
 sg13g2_fill_1 FILLER_167_1767 ();
 sg13g2_decap_8 FILLER_168_0 ();
 sg13g2_decap_8 FILLER_168_7 ();
 sg13g2_decap_8 FILLER_168_14 ();
 sg13g2_decap_8 FILLER_168_21 ();
 sg13g2_decap_8 FILLER_168_28 ();
 sg13g2_decap_8 FILLER_168_35 ();
 sg13g2_decap_8 FILLER_168_42 ();
 sg13g2_decap_8 FILLER_168_49 ();
 sg13g2_decap_8 FILLER_168_56 ();
 sg13g2_decap_8 FILLER_168_63 ();
 sg13g2_decap_8 FILLER_168_70 ();
 sg13g2_decap_8 FILLER_168_77 ();
 sg13g2_decap_8 FILLER_168_84 ();
 sg13g2_decap_8 FILLER_168_91 ();
 sg13g2_decap_8 FILLER_168_98 ();
 sg13g2_decap_8 FILLER_168_105 ();
 sg13g2_decap_8 FILLER_168_112 ();
 sg13g2_decap_8 FILLER_168_119 ();
 sg13g2_decap_8 FILLER_168_126 ();
 sg13g2_decap_8 FILLER_168_133 ();
 sg13g2_decap_8 FILLER_168_140 ();
 sg13g2_decap_8 FILLER_168_147 ();
 sg13g2_decap_8 FILLER_168_154 ();
 sg13g2_decap_8 FILLER_168_161 ();
 sg13g2_decap_8 FILLER_168_168 ();
 sg13g2_decap_8 FILLER_168_178 ();
 sg13g2_decap_8 FILLER_168_185 ();
 sg13g2_decap_8 FILLER_168_192 ();
 sg13g2_decap_8 FILLER_168_199 ();
 sg13g2_decap_4 FILLER_168_206 ();
 sg13g2_fill_2 FILLER_168_210 ();
 sg13g2_decap_8 FILLER_168_222 ();
 sg13g2_decap_8 FILLER_168_229 ();
 sg13g2_decap_8 FILLER_168_236 ();
 sg13g2_decap_8 FILLER_168_247 ();
 sg13g2_decap_8 FILLER_168_274 ();
 sg13g2_decap_8 FILLER_168_281 ();
 sg13g2_decap_8 FILLER_168_288 ();
 sg13g2_decap_8 FILLER_168_295 ();
 sg13g2_decap_8 FILLER_168_302 ();
 sg13g2_decap_8 FILLER_168_309 ();
 sg13g2_decap_8 FILLER_168_316 ();
 sg13g2_decap_8 FILLER_168_323 ();
 sg13g2_decap_4 FILLER_168_330 ();
 sg13g2_fill_2 FILLER_168_339 ();
 sg13g2_fill_1 FILLER_168_348 ();
 sg13g2_fill_1 FILLER_168_354 ();
 sg13g2_fill_2 FILLER_168_363 ();
 sg13g2_fill_1 FILLER_168_365 ();
 sg13g2_decap_8 FILLER_168_384 ();
 sg13g2_decap_8 FILLER_168_391 ();
 sg13g2_decap_8 FILLER_168_398 ();
 sg13g2_fill_2 FILLER_168_405 ();
 sg13g2_fill_1 FILLER_168_407 ();
 sg13g2_fill_2 FILLER_168_416 ();
 sg13g2_decap_8 FILLER_168_431 ();
 sg13g2_fill_2 FILLER_168_438 ();
 sg13g2_fill_1 FILLER_168_440 ();
 sg13g2_decap_8 FILLER_168_444 ();
 sg13g2_decap_4 FILLER_168_451 ();
 sg13g2_decap_8 FILLER_168_471 ();
 sg13g2_decap_8 FILLER_168_478 ();
 sg13g2_decap_8 FILLER_168_485 ();
 sg13g2_decap_8 FILLER_168_492 ();
 sg13g2_decap_8 FILLER_168_499 ();
 sg13g2_fill_1 FILLER_168_506 ();
 sg13g2_fill_1 FILLER_168_511 ();
 sg13g2_decap_8 FILLER_168_536 ();
 sg13g2_decap_8 FILLER_168_543 ();
 sg13g2_decap_8 FILLER_168_550 ();
 sg13g2_decap_4 FILLER_168_557 ();
 sg13g2_fill_1 FILLER_168_561 ();
 sg13g2_fill_2 FILLER_168_566 ();
 sg13g2_fill_1 FILLER_168_568 ();
 sg13g2_decap_8 FILLER_168_572 ();
 sg13g2_decap_8 FILLER_168_579 ();
 sg13g2_decap_8 FILLER_168_586 ();
 sg13g2_decap_8 FILLER_168_593 ();
 sg13g2_decap_8 FILLER_168_600 ();
 sg13g2_decap_8 FILLER_168_607 ();
 sg13g2_decap_8 FILLER_168_614 ();
 sg13g2_decap_8 FILLER_168_621 ();
 sg13g2_fill_1 FILLER_168_628 ();
 sg13g2_decap_8 FILLER_168_665 ();
 sg13g2_decap_8 FILLER_168_672 ();
 sg13g2_decap_8 FILLER_168_679 ();
 sg13g2_decap_8 FILLER_168_686 ();
 sg13g2_decap_4 FILLER_168_693 ();
 sg13g2_fill_2 FILLER_168_697 ();
 sg13g2_fill_1 FILLER_168_703 ();
 sg13g2_fill_1 FILLER_168_718 ();
 sg13g2_decap_8 FILLER_168_729 ();
 sg13g2_decap_8 FILLER_168_736 ();
 sg13g2_decap_8 FILLER_168_743 ();
 sg13g2_decap_8 FILLER_168_750 ();
 sg13g2_decap_8 FILLER_168_757 ();
 sg13g2_decap_8 FILLER_168_764 ();
 sg13g2_decap_8 FILLER_168_771 ();
 sg13g2_fill_2 FILLER_168_778 ();
 sg13g2_decap_4 FILLER_168_800 ();
 sg13g2_fill_1 FILLER_168_804 ();
 sg13g2_fill_1 FILLER_168_810 ();
 sg13g2_decap_8 FILLER_168_816 ();
 sg13g2_fill_2 FILLER_168_823 ();
 sg13g2_fill_2 FILLER_168_835 ();
 sg13g2_fill_1 FILLER_168_863 ();
 sg13g2_decap_8 FILLER_168_872 ();
 sg13g2_decap_8 FILLER_168_879 ();
 sg13g2_decap_8 FILLER_168_886 ();
 sg13g2_decap_4 FILLER_168_893 ();
 sg13g2_fill_1 FILLER_168_897 ();
 sg13g2_decap_4 FILLER_168_910 ();
 sg13g2_decap_8 FILLER_168_926 ();
 sg13g2_decap_8 FILLER_168_933 ();
 sg13g2_decap_8 FILLER_168_940 ();
 sg13g2_decap_8 FILLER_168_947 ();
 sg13g2_decap_8 FILLER_168_954 ();
 sg13g2_decap_8 FILLER_168_961 ();
 sg13g2_decap_8 FILLER_168_968 ();
 sg13g2_decap_8 FILLER_168_975 ();
 sg13g2_decap_8 FILLER_168_982 ();
 sg13g2_decap_8 FILLER_168_989 ();
 sg13g2_decap_8 FILLER_168_996 ();
 sg13g2_decap_8 FILLER_168_1003 ();
 sg13g2_decap_8 FILLER_168_1010 ();
 sg13g2_decap_8 FILLER_168_1029 ();
 sg13g2_decap_8 FILLER_168_1036 ();
 sg13g2_decap_8 FILLER_168_1043 ();
 sg13g2_decap_8 FILLER_168_1050 ();
 sg13g2_decap_8 FILLER_168_1057 ();
 sg13g2_fill_2 FILLER_168_1064 ();
 sg13g2_fill_1 FILLER_168_1084 ();
 sg13g2_fill_2 FILLER_168_1093 ();
 sg13g2_decap_8 FILLER_168_1118 ();
 sg13g2_decap_8 FILLER_168_1125 ();
 sg13g2_decap_8 FILLER_168_1132 ();
 sg13g2_fill_2 FILLER_168_1139 ();
 sg13g2_fill_1 FILLER_168_1141 ();
 sg13g2_decap_8 FILLER_168_1154 ();
 sg13g2_decap_4 FILLER_168_1161 ();
 sg13g2_fill_1 FILLER_168_1165 ();
 sg13g2_decap_8 FILLER_168_1174 ();
 sg13g2_decap_8 FILLER_168_1181 ();
 sg13g2_decap_8 FILLER_168_1188 ();
 sg13g2_fill_2 FILLER_168_1195 ();
 sg13g2_decap_8 FILLER_168_1202 ();
 sg13g2_decap_8 FILLER_168_1209 ();
 sg13g2_decap_8 FILLER_168_1216 ();
 sg13g2_decap_8 FILLER_168_1223 ();
 sg13g2_decap_8 FILLER_168_1238 ();
 sg13g2_decap_8 FILLER_168_1245 ();
 sg13g2_fill_2 FILLER_168_1252 ();
 sg13g2_fill_1 FILLER_168_1254 ();
 sg13g2_decap_8 FILLER_168_1263 ();
 sg13g2_decap_8 FILLER_168_1270 ();
 sg13g2_decap_8 FILLER_168_1277 ();
 sg13g2_decap_8 FILLER_168_1284 ();
 sg13g2_decap_8 FILLER_168_1291 ();
 sg13g2_decap_8 FILLER_168_1298 ();
 sg13g2_decap_8 FILLER_168_1305 ();
 sg13g2_decap_8 FILLER_168_1312 ();
 sg13g2_decap_8 FILLER_168_1319 ();
 sg13g2_decap_8 FILLER_168_1326 ();
 sg13g2_decap_8 FILLER_168_1333 ();
 sg13g2_decap_8 FILLER_168_1340 ();
 sg13g2_decap_8 FILLER_168_1347 ();
 sg13g2_decap_8 FILLER_168_1354 ();
 sg13g2_decap_8 FILLER_168_1361 ();
 sg13g2_decap_8 FILLER_168_1368 ();
 sg13g2_decap_8 FILLER_168_1375 ();
 sg13g2_decap_8 FILLER_168_1382 ();
 sg13g2_decap_8 FILLER_168_1389 ();
 sg13g2_decap_8 FILLER_168_1396 ();
 sg13g2_decap_8 FILLER_168_1403 ();
 sg13g2_decap_8 FILLER_168_1410 ();
 sg13g2_decap_8 FILLER_168_1417 ();
 sg13g2_decap_8 FILLER_168_1424 ();
 sg13g2_decap_8 FILLER_168_1431 ();
 sg13g2_decap_8 FILLER_168_1438 ();
 sg13g2_decap_8 FILLER_168_1445 ();
 sg13g2_decap_8 FILLER_168_1452 ();
 sg13g2_decap_8 FILLER_168_1459 ();
 sg13g2_decap_8 FILLER_168_1466 ();
 sg13g2_decap_8 FILLER_168_1473 ();
 sg13g2_decap_8 FILLER_168_1480 ();
 sg13g2_decap_8 FILLER_168_1487 ();
 sg13g2_decap_8 FILLER_168_1494 ();
 sg13g2_decap_8 FILLER_168_1501 ();
 sg13g2_decap_8 FILLER_168_1508 ();
 sg13g2_decap_8 FILLER_168_1515 ();
 sg13g2_decap_8 FILLER_168_1522 ();
 sg13g2_decap_8 FILLER_168_1529 ();
 sg13g2_decap_8 FILLER_168_1536 ();
 sg13g2_decap_8 FILLER_168_1543 ();
 sg13g2_decap_8 FILLER_168_1550 ();
 sg13g2_decap_8 FILLER_168_1557 ();
 sg13g2_decap_8 FILLER_168_1564 ();
 sg13g2_decap_8 FILLER_168_1571 ();
 sg13g2_decap_8 FILLER_168_1578 ();
 sg13g2_decap_8 FILLER_168_1585 ();
 sg13g2_decap_8 FILLER_168_1592 ();
 sg13g2_decap_8 FILLER_168_1599 ();
 sg13g2_decap_8 FILLER_168_1606 ();
 sg13g2_decap_8 FILLER_168_1613 ();
 sg13g2_decap_8 FILLER_168_1620 ();
 sg13g2_decap_8 FILLER_168_1627 ();
 sg13g2_decap_8 FILLER_168_1634 ();
 sg13g2_decap_8 FILLER_168_1641 ();
 sg13g2_decap_8 FILLER_168_1648 ();
 sg13g2_decap_8 FILLER_168_1655 ();
 sg13g2_decap_8 FILLER_168_1662 ();
 sg13g2_decap_8 FILLER_168_1669 ();
 sg13g2_decap_8 FILLER_168_1676 ();
 sg13g2_decap_8 FILLER_168_1683 ();
 sg13g2_decap_8 FILLER_168_1690 ();
 sg13g2_decap_8 FILLER_168_1697 ();
 sg13g2_decap_8 FILLER_168_1704 ();
 sg13g2_decap_8 FILLER_168_1711 ();
 sg13g2_decap_8 FILLER_168_1718 ();
 sg13g2_decap_8 FILLER_168_1725 ();
 sg13g2_decap_8 FILLER_168_1732 ();
 sg13g2_decap_8 FILLER_168_1739 ();
 sg13g2_decap_8 FILLER_168_1746 ();
 sg13g2_decap_8 FILLER_168_1753 ();
 sg13g2_decap_8 FILLER_168_1760 ();
 sg13g2_fill_1 FILLER_168_1767 ();
 sg13g2_decap_8 FILLER_169_0 ();
 sg13g2_decap_8 FILLER_169_7 ();
 sg13g2_decap_8 FILLER_169_14 ();
 sg13g2_decap_8 FILLER_169_21 ();
 sg13g2_decap_8 FILLER_169_28 ();
 sg13g2_decap_8 FILLER_169_35 ();
 sg13g2_decap_8 FILLER_169_42 ();
 sg13g2_decap_8 FILLER_169_49 ();
 sg13g2_decap_8 FILLER_169_56 ();
 sg13g2_decap_8 FILLER_169_63 ();
 sg13g2_decap_8 FILLER_169_70 ();
 sg13g2_decap_8 FILLER_169_77 ();
 sg13g2_decap_8 FILLER_169_84 ();
 sg13g2_decap_8 FILLER_169_91 ();
 sg13g2_decap_8 FILLER_169_98 ();
 sg13g2_decap_8 FILLER_169_105 ();
 sg13g2_decap_8 FILLER_169_112 ();
 sg13g2_decap_8 FILLER_169_119 ();
 sg13g2_decap_8 FILLER_169_126 ();
 sg13g2_decap_8 FILLER_169_133 ();
 sg13g2_decap_8 FILLER_169_140 ();
 sg13g2_decap_8 FILLER_169_147 ();
 sg13g2_decap_8 FILLER_169_154 ();
 sg13g2_decap_8 FILLER_169_161 ();
 sg13g2_decap_8 FILLER_169_168 ();
 sg13g2_decap_8 FILLER_169_175 ();
 sg13g2_decap_8 FILLER_169_182 ();
 sg13g2_decap_8 FILLER_169_189 ();
 sg13g2_decap_8 FILLER_169_196 ();
 sg13g2_decap_8 FILLER_169_203 ();
 sg13g2_decap_8 FILLER_169_210 ();
 sg13g2_decap_8 FILLER_169_217 ();
 sg13g2_decap_4 FILLER_169_224 ();
 sg13g2_fill_2 FILLER_169_228 ();
 sg13g2_decap_8 FILLER_169_241 ();
 sg13g2_decap_8 FILLER_169_248 ();
 sg13g2_decap_8 FILLER_169_255 ();
 sg13g2_decap_8 FILLER_169_262 ();
 sg13g2_decap_8 FILLER_169_292 ();
 sg13g2_decap_8 FILLER_169_299 ();
 sg13g2_decap_8 FILLER_169_306 ();
 sg13g2_decap_8 FILLER_169_313 ();
 sg13g2_decap_8 FILLER_169_320 ();
 sg13g2_decap_4 FILLER_169_327 ();
 sg13g2_fill_2 FILLER_169_331 ();
 sg13g2_fill_2 FILLER_169_352 ();
 sg13g2_fill_1 FILLER_169_354 ();
 sg13g2_fill_2 FILLER_169_363 ();
 sg13g2_decap_8 FILLER_169_375 ();
 sg13g2_decap_8 FILLER_169_382 ();
 sg13g2_decap_8 FILLER_169_389 ();
 sg13g2_decap_8 FILLER_169_396 ();
 sg13g2_decap_8 FILLER_169_403 ();
 sg13g2_fill_2 FILLER_169_410 ();
 sg13g2_fill_1 FILLER_169_412 ();
 sg13g2_decap_8 FILLER_169_421 ();
 sg13g2_fill_1 FILLER_169_428 ();
 sg13g2_decap_8 FILLER_169_439 ();
 sg13g2_decap_8 FILLER_169_446 ();
 sg13g2_fill_1 FILLER_169_461 ();
 sg13g2_decap_8 FILLER_169_486 ();
 sg13g2_decap_8 FILLER_169_493 ();
 sg13g2_decap_8 FILLER_169_500 ();
 sg13g2_decap_8 FILLER_169_507 ();
 sg13g2_fill_2 FILLER_169_514 ();
 sg13g2_decap_8 FILLER_169_532 ();
 sg13g2_decap_8 FILLER_169_539 ();
 sg13g2_decap_8 FILLER_169_546 ();
 sg13g2_fill_1 FILLER_169_553 ();
 sg13g2_fill_2 FILLER_169_562 ();
 sg13g2_decap_4 FILLER_169_581 ();
 sg13g2_fill_1 FILLER_169_585 ();
 sg13g2_decap_8 FILLER_169_589 ();
 sg13g2_decap_8 FILLER_169_596 ();
 sg13g2_decap_8 FILLER_169_603 ();
 sg13g2_decap_8 FILLER_169_610 ();
 sg13g2_decap_8 FILLER_169_617 ();
 sg13g2_decap_8 FILLER_169_624 ();
 sg13g2_decap_8 FILLER_169_631 ();
 sg13g2_decap_8 FILLER_169_638 ();
 sg13g2_fill_2 FILLER_169_645 ();
 sg13g2_decap_4 FILLER_169_682 ();
 sg13g2_fill_2 FILLER_169_701 ();
 sg13g2_fill_1 FILLER_169_703 ();
 sg13g2_decap_8 FILLER_169_730 ();
 sg13g2_decap_8 FILLER_169_737 ();
 sg13g2_decap_8 FILLER_169_744 ();
 sg13g2_decap_8 FILLER_169_751 ();
 sg13g2_decap_8 FILLER_169_758 ();
 sg13g2_decap_8 FILLER_169_765 ();
 sg13g2_decap_8 FILLER_169_772 ();
 sg13g2_decap_4 FILLER_169_779 ();
 sg13g2_fill_1 FILLER_169_783 ();
 sg13g2_decap_8 FILLER_169_789 ();
 sg13g2_fill_2 FILLER_169_796 ();
 sg13g2_fill_1 FILLER_169_798 ();
 sg13g2_fill_1 FILLER_169_823 ();
 sg13g2_fill_2 FILLER_169_840 ();
 sg13g2_fill_2 FILLER_169_847 ();
 sg13g2_fill_1 FILLER_169_857 ();
 sg13g2_fill_1 FILLER_169_874 ();
 sg13g2_fill_1 FILLER_169_879 ();
 sg13g2_decap_8 FILLER_169_892 ();
 sg13g2_decap_8 FILLER_169_899 ();
 sg13g2_fill_1 FILLER_169_918 ();
 sg13g2_decap_8 FILLER_169_937 ();
 sg13g2_decap_8 FILLER_169_944 ();
 sg13g2_decap_8 FILLER_169_951 ();
 sg13g2_decap_8 FILLER_169_958 ();
 sg13g2_decap_8 FILLER_169_965 ();
 sg13g2_decap_8 FILLER_169_972 ();
 sg13g2_decap_8 FILLER_169_979 ();
 sg13g2_decap_8 FILLER_169_986 ();
 sg13g2_decap_8 FILLER_169_993 ();
 sg13g2_decap_8 FILLER_169_1000 ();
 sg13g2_decap_4 FILLER_169_1007 ();
 sg13g2_fill_1 FILLER_169_1011 ();
 sg13g2_decap_8 FILLER_169_1038 ();
 sg13g2_decap_8 FILLER_169_1045 ();
 sg13g2_decap_8 FILLER_169_1052 ();
 sg13g2_fill_2 FILLER_169_1071 ();
 sg13g2_fill_1 FILLER_169_1081 ();
 sg13g2_fill_2 FILLER_169_1092 ();
 sg13g2_fill_1 FILLER_169_1094 ();
 sg13g2_decap_8 FILLER_169_1103 ();
 sg13g2_decap_8 FILLER_169_1110 ();
 sg13g2_decap_4 FILLER_169_1117 ();
 sg13g2_fill_1 FILLER_169_1121 ();
 sg13g2_decap_8 FILLER_169_1131 ();
 sg13g2_decap_8 FILLER_169_1138 ();
 sg13g2_decap_8 FILLER_169_1145 ();
 sg13g2_decap_8 FILLER_169_1152 ();
 sg13g2_decap_8 FILLER_169_1159 ();
 sg13g2_decap_8 FILLER_169_1166 ();
 sg13g2_decap_8 FILLER_169_1173 ();
 sg13g2_decap_8 FILLER_169_1180 ();
 sg13g2_decap_8 FILLER_169_1187 ();
 sg13g2_fill_1 FILLER_169_1198 ();
 sg13g2_decap_8 FILLER_169_1207 ();
 sg13g2_decap_8 FILLER_169_1214 ();
 sg13g2_decap_8 FILLER_169_1221 ();
 sg13g2_decap_8 FILLER_169_1228 ();
 sg13g2_decap_8 FILLER_169_1235 ();
 sg13g2_decap_8 FILLER_169_1242 ();
 sg13g2_decap_8 FILLER_169_1249 ();
 sg13g2_decap_8 FILLER_169_1256 ();
 sg13g2_decap_8 FILLER_169_1263 ();
 sg13g2_decap_8 FILLER_169_1270 ();
 sg13g2_decap_8 FILLER_169_1277 ();
 sg13g2_decap_8 FILLER_169_1284 ();
 sg13g2_decap_8 FILLER_169_1291 ();
 sg13g2_decap_8 FILLER_169_1298 ();
 sg13g2_decap_8 FILLER_169_1305 ();
 sg13g2_decap_8 FILLER_169_1312 ();
 sg13g2_decap_8 FILLER_169_1319 ();
 sg13g2_decap_8 FILLER_169_1326 ();
 sg13g2_decap_8 FILLER_169_1333 ();
 sg13g2_decap_8 FILLER_169_1340 ();
 sg13g2_decap_8 FILLER_169_1347 ();
 sg13g2_decap_8 FILLER_169_1354 ();
 sg13g2_decap_8 FILLER_169_1361 ();
 sg13g2_decap_8 FILLER_169_1368 ();
 sg13g2_decap_8 FILLER_169_1375 ();
 sg13g2_decap_8 FILLER_169_1382 ();
 sg13g2_decap_8 FILLER_169_1389 ();
 sg13g2_decap_8 FILLER_169_1396 ();
 sg13g2_decap_8 FILLER_169_1403 ();
 sg13g2_decap_8 FILLER_169_1410 ();
 sg13g2_decap_8 FILLER_169_1417 ();
 sg13g2_decap_8 FILLER_169_1424 ();
 sg13g2_decap_8 FILLER_169_1431 ();
 sg13g2_decap_8 FILLER_169_1438 ();
 sg13g2_decap_8 FILLER_169_1445 ();
 sg13g2_decap_8 FILLER_169_1452 ();
 sg13g2_decap_8 FILLER_169_1459 ();
 sg13g2_decap_8 FILLER_169_1466 ();
 sg13g2_decap_8 FILLER_169_1473 ();
 sg13g2_decap_8 FILLER_169_1480 ();
 sg13g2_decap_8 FILLER_169_1487 ();
 sg13g2_decap_8 FILLER_169_1494 ();
 sg13g2_decap_8 FILLER_169_1501 ();
 sg13g2_decap_8 FILLER_169_1508 ();
 sg13g2_decap_8 FILLER_169_1515 ();
 sg13g2_decap_8 FILLER_169_1522 ();
 sg13g2_decap_8 FILLER_169_1529 ();
 sg13g2_decap_8 FILLER_169_1536 ();
 sg13g2_decap_8 FILLER_169_1543 ();
 sg13g2_decap_8 FILLER_169_1550 ();
 sg13g2_decap_8 FILLER_169_1557 ();
 sg13g2_decap_8 FILLER_169_1564 ();
 sg13g2_decap_8 FILLER_169_1571 ();
 sg13g2_decap_8 FILLER_169_1578 ();
 sg13g2_decap_8 FILLER_169_1585 ();
 sg13g2_decap_8 FILLER_169_1592 ();
 sg13g2_decap_8 FILLER_169_1599 ();
 sg13g2_decap_8 FILLER_169_1606 ();
 sg13g2_decap_8 FILLER_169_1613 ();
 sg13g2_decap_8 FILLER_169_1620 ();
 sg13g2_decap_8 FILLER_169_1627 ();
 sg13g2_decap_8 FILLER_169_1634 ();
 sg13g2_decap_8 FILLER_169_1641 ();
 sg13g2_decap_8 FILLER_169_1648 ();
 sg13g2_decap_8 FILLER_169_1655 ();
 sg13g2_decap_8 FILLER_169_1662 ();
 sg13g2_decap_8 FILLER_169_1669 ();
 sg13g2_decap_8 FILLER_169_1676 ();
 sg13g2_decap_8 FILLER_169_1683 ();
 sg13g2_decap_8 FILLER_169_1690 ();
 sg13g2_decap_8 FILLER_169_1697 ();
 sg13g2_decap_8 FILLER_169_1704 ();
 sg13g2_decap_8 FILLER_169_1711 ();
 sg13g2_decap_8 FILLER_169_1718 ();
 sg13g2_decap_8 FILLER_169_1725 ();
 sg13g2_decap_8 FILLER_169_1732 ();
 sg13g2_decap_8 FILLER_169_1739 ();
 sg13g2_decap_8 FILLER_169_1746 ();
 sg13g2_decap_8 FILLER_169_1753 ();
 sg13g2_decap_8 FILLER_169_1760 ();
 sg13g2_fill_1 FILLER_169_1767 ();
 sg13g2_decap_8 FILLER_170_0 ();
 sg13g2_decap_8 FILLER_170_7 ();
 sg13g2_decap_8 FILLER_170_14 ();
 sg13g2_decap_8 FILLER_170_21 ();
 sg13g2_decap_8 FILLER_170_28 ();
 sg13g2_decap_8 FILLER_170_35 ();
 sg13g2_decap_8 FILLER_170_42 ();
 sg13g2_decap_8 FILLER_170_49 ();
 sg13g2_decap_8 FILLER_170_56 ();
 sg13g2_decap_8 FILLER_170_63 ();
 sg13g2_decap_8 FILLER_170_70 ();
 sg13g2_decap_8 FILLER_170_77 ();
 sg13g2_decap_8 FILLER_170_84 ();
 sg13g2_decap_8 FILLER_170_91 ();
 sg13g2_decap_8 FILLER_170_98 ();
 sg13g2_decap_8 FILLER_170_105 ();
 sg13g2_decap_8 FILLER_170_112 ();
 sg13g2_decap_8 FILLER_170_119 ();
 sg13g2_decap_8 FILLER_170_126 ();
 sg13g2_decap_8 FILLER_170_133 ();
 sg13g2_decap_8 FILLER_170_140 ();
 sg13g2_decap_8 FILLER_170_147 ();
 sg13g2_decap_8 FILLER_170_154 ();
 sg13g2_decap_8 FILLER_170_161 ();
 sg13g2_decap_8 FILLER_170_168 ();
 sg13g2_fill_2 FILLER_170_175 ();
 sg13g2_fill_1 FILLER_170_177 ();
 sg13g2_decap_8 FILLER_170_197 ();
 sg13g2_decap_8 FILLER_170_204 ();
 sg13g2_decap_8 FILLER_170_211 ();
 sg13g2_fill_2 FILLER_170_218 ();
 sg13g2_decap_8 FILLER_170_223 ();
 sg13g2_decap_8 FILLER_170_230 ();
 sg13g2_decap_8 FILLER_170_237 ();
 sg13g2_decap_8 FILLER_170_244 ();
 sg13g2_decap_8 FILLER_170_251 ();
 sg13g2_decap_8 FILLER_170_258 ();
 sg13g2_fill_2 FILLER_170_265 ();
 sg13g2_fill_1 FILLER_170_267 ();
 sg13g2_fill_2 FILLER_170_274 ();
 sg13g2_fill_1 FILLER_170_276 ();
 sg13g2_fill_2 FILLER_170_282 ();
 sg13g2_decap_8 FILLER_170_300 ();
 sg13g2_decap_8 FILLER_170_307 ();
 sg13g2_decap_4 FILLER_170_314 ();
 sg13g2_fill_1 FILLER_170_318 ();
 sg13g2_decap_8 FILLER_170_331 ();
 sg13g2_fill_2 FILLER_170_338 ();
 sg13g2_fill_1 FILLER_170_340 ();
 sg13g2_decap_8 FILLER_170_350 ();
 sg13g2_decap_8 FILLER_170_357 ();
 sg13g2_decap_8 FILLER_170_364 ();
 sg13g2_decap_8 FILLER_170_371 ();
 sg13g2_decap_8 FILLER_170_378 ();
 sg13g2_decap_8 FILLER_170_385 ();
 sg13g2_decap_8 FILLER_170_392 ();
 sg13g2_decap_8 FILLER_170_399 ();
 sg13g2_decap_8 FILLER_170_416 ();
 sg13g2_decap_8 FILLER_170_423 ();
 sg13g2_decap_8 FILLER_170_438 ();
 sg13g2_decap_8 FILLER_170_445 ();
 sg13g2_decap_8 FILLER_170_452 ();
 sg13g2_decap_8 FILLER_170_459 ();
 sg13g2_decap_4 FILLER_170_474 ();
 sg13g2_fill_2 FILLER_170_478 ();
 sg13g2_decap_8 FILLER_170_488 ();
 sg13g2_decap_8 FILLER_170_495 ();
 sg13g2_decap_8 FILLER_170_502 ();
 sg13g2_decap_8 FILLER_170_509 ();
 sg13g2_fill_1 FILLER_170_516 ();
 sg13g2_decap_8 FILLER_170_534 ();
 sg13g2_decap_8 FILLER_170_541 ();
 sg13g2_decap_8 FILLER_170_548 ();
 sg13g2_decap_8 FILLER_170_555 ();
 sg13g2_fill_1 FILLER_170_566 ();
 sg13g2_decap_4 FILLER_170_572 ();
 sg13g2_fill_1 FILLER_170_584 ();
 sg13g2_decap_8 FILLER_170_593 ();
 sg13g2_decap_8 FILLER_170_600 ();
 sg13g2_decap_8 FILLER_170_607 ();
 sg13g2_decap_8 FILLER_170_614 ();
 sg13g2_decap_8 FILLER_170_621 ();
 sg13g2_decap_8 FILLER_170_628 ();
 sg13g2_decap_4 FILLER_170_635 ();
 sg13g2_fill_1 FILLER_170_639 ();
 sg13g2_decap_8 FILLER_170_644 ();
 sg13g2_fill_1 FILLER_170_651 ();
 sg13g2_decap_8 FILLER_170_669 ();
 sg13g2_decap_4 FILLER_170_676 ();
 sg13g2_fill_2 FILLER_170_680 ();
 sg13g2_decap_8 FILLER_170_708 ();
 sg13g2_decap_8 FILLER_170_715 ();
 sg13g2_decap_8 FILLER_170_722 ();
 sg13g2_decap_8 FILLER_170_729 ();
 sg13g2_decap_8 FILLER_170_736 ();
 sg13g2_decap_8 FILLER_170_743 ();
 sg13g2_decap_8 FILLER_170_750 ();
 sg13g2_decap_8 FILLER_170_757 ();
 sg13g2_decap_8 FILLER_170_764 ();
 sg13g2_fill_2 FILLER_170_771 ();
 sg13g2_fill_1 FILLER_170_773 ();
 sg13g2_decap_8 FILLER_170_782 ();
 sg13g2_decap_8 FILLER_170_789 ();
 sg13g2_decap_8 FILLER_170_796 ();
 sg13g2_decap_8 FILLER_170_803 ();
 sg13g2_decap_8 FILLER_170_810 ();
 sg13g2_decap_8 FILLER_170_817 ();
 sg13g2_decap_8 FILLER_170_824 ();
 sg13g2_decap_8 FILLER_170_831 ();
 sg13g2_decap_8 FILLER_170_838 ();
 sg13g2_fill_2 FILLER_170_849 ();
 sg13g2_fill_1 FILLER_170_851 ();
 sg13g2_decap_4 FILLER_170_860 ();
 sg13g2_decap_8 FILLER_170_868 ();
 sg13g2_decap_4 FILLER_170_875 ();
 sg13g2_fill_1 FILLER_170_879 ();
 sg13g2_decap_8 FILLER_170_892 ();
 sg13g2_decap_8 FILLER_170_899 ();
 sg13g2_fill_1 FILLER_170_906 ();
 sg13g2_decap_8 FILLER_170_935 ();
 sg13g2_decap_8 FILLER_170_942 ();
 sg13g2_decap_8 FILLER_170_949 ();
 sg13g2_decap_4 FILLER_170_956 ();
 sg13g2_fill_1 FILLER_170_960 ();
 sg13g2_decap_4 FILLER_170_976 ();
 sg13g2_fill_1 FILLER_170_980 ();
 sg13g2_decap_4 FILLER_170_985 ();
 sg13g2_fill_1 FILLER_170_989 ();
 sg13g2_decap_8 FILLER_170_999 ();
 sg13g2_decap_8 FILLER_170_1006 ();
 sg13g2_decap_8 FILLER_170_1013 ();
 sg13g2_fill_2 FILLER_170_1034 ();
 sg13g2_decap_8 FILLER_170_1040 ();
 sg13g2_decap_8 FILLER_170_1047 ();
 sg13g2_decap_8 FILLER_170_1054 ();
 sg13g2_fill_2 FILLER_170_1061 ();
 sg13g2_fill_1 FILLER_170_1063 ();
 sg13g2_decap_8 FILLER_170_1069 ();
 sg13g2_decap_4 FILLER_170_1076 ();
 sg13g2_fill_1 FILLER_170_1080 ();
 sg13g2_decap_8 FILLER_170_1101 ();
 sg13g2_decap_8 FILLER_170_1108 ();
 sg13g2_decap_8 FILLER_170_1115 ();
 sg13g2_decap_8 FILLER_170_1122 ();
 sg13g2_fill_2 FILLER_170_1129 ();
 sg13g2_fill_1 FILLER_170_1131 ();
 sg13g2_decap_8 FILLER_170_1148 ();
 sg13g2_decap_8 FILLER_170_1155 ();
 sg13g2_decap_8 FILLER_170_1162 ();
 sg13g2_decap_8 FILLER_170_1169 ();
 sg13g2_decap_8 FILLER_170_1176 ();
 sg13g2_fill_2 FILLER_170_1199 ();
 sg13g2_decap_8 FILLER_170_1209 ();
 sg13g2_decap_8 FILLER_170_1216 ();
 sg13g2_decap_8 FILLER_170_1223 ();
 sg13g2_decap_8 FILLER_170_1230 ();
 sg13g2_decap_8 FILLER_170_1237 ();
 sg13g2_decap_8 FILLER_170_1244 ();
 sg13g2_decap_8 FILLER_170_1251 ();
 sg13g2_decap_8 FILLER_170_1258 ();
 sg13g2_decap_8 FILLER_170_1265 ();
 sg13g2_decap_8 FILLER_170_1272 ();
 sg13g2_decap_8 FILLER_170_1279 ();
 sg13g2_decap_8 FILLER_170_1286 ();
 sg13g2_decap_8 FILLER_170_1293 ();
 sg13g2_decap_8 FILLER_170_1300 ();
 sg13g2_decap_8 FILLER_170_1307 ();
 sg13g2_decap_8 FILLER_170_1314 ();
 sg13g2_decap_8 FILLER_170_1321 ();
 sg13g2_decap_8 FILLER_170_1328 ();
 sg13g2_decap_8 FILLER_170_1335 ();
 sg13g2_decap_8 FILLER_170_1342 ();
 sg13g2_decap_8 FILLER_170_1349 ();
 sg13g2_decap_8 FILLER_170_1356 ();
 sg13g2_decap_8 FILLER_170_1363 ();
 sg13g2_decap_8 FILLER_170_1370 ();
 sg13g2_decap_8 FILLER_170_1377 ();
 sg13g2_decap_8 FILLER_170_1384 ();
 sg13g2_decap_8 FILLER_170_1391 ();
 sg13g2_decap_8 FILLER_170_1398 ();
 sg13g2_decap_8 FILLER_170_1405 ();
 sg13g2_decap_8 FILLER_170_1412 ();
 sg13g2_decap_8 FILLER_170_1419 ();
 sg13g2_decap_8 FILLER_170_1426 ();
 sg13g2_decap_8 FILLER_170_1433 ();
 sg13g2_decap_8 FILLER_170_1440 ();
 sg13g2_decap_8 FILLER_170_1447 ();
 sg13g2_decap_8 FILLER_170_1454 ();
 sg13g2_decap_8 FILLER_170_1461 ();
 sg13g2_decap_8 FILLER_170_1468 ();
 sg13g2_decap_8 FILLER_170_1475 ();
 sg13g2_decap_8 FILLER_170_1482 ();
 sg13g2_decap_8 FILLER_170_1489 ();
 sg13g2_decap_8 FILLER_170_1496 ();
 sg13g2_decap_8 FILLER_170_1503 ();
 sg13g2_decap_8 FILLER_170_1510 ();
 sg13g2_decap_8 FILLER_170_1517 ();
 sg13g2_decap_8 FILLER_170_1524 ();
 sg13g2_decap_8 FILLER_170_1531 ();
 sg13g2_decap_8 FILLER_170_1538 ();
 sg13g2_decap_8 FILLER_170_1545 ();
 sg13g2_decap_8 FILLER_170_1552 ();
 sg13g2_decap_8 FILLER_170_1559 ();
 sg13g2_decap_8 FILLER_170_1566 ();
 sg13g2_decap_8 FILLER_170_1573 ();
 sg13g2_decap_8 FILLER_170_1580 ();
 sg13g2_decap_8 FILLER_170_1587 ();
 sg13g2_decap_8 FILLER_170_1594 ();
 sg13g2_decap_8 FILLER_170_1601 ();
 sg13g2_decap_8 FILLER_170_1608 ();
 sg13g2_decap_8 FILLER_170_1615 ();
 sg13g2_decap_8 FILLER_170_1622 ();
 sg13g2_decap_8 FILLER_170_1629 ();
 sg13g2_decap_8 FILLER_170_1636 ();
 sg13g2_decap_8 FILLER_170_1643 ();
 sg13g2_decap_8 FILLER_170_1650 ();
 sg13g2_decap_8 FILLER_170_1657 ();
 sg13g2_decap_8 FILLER_170_1664 ();
 sg13g2_decap_8 FILLER_170_1671 ();
 sg13g2_decap_8 FILLER_170_1678 ();
 sg13g2_decap_8 FILLER_170_1685 ();
 sg13g2_decap_8 FILLER_170_1692 ();
 sg13g2_decap_8 FILLER_170_1699 ();
 sg13g2_decap_8 FILLER_170_1706 ();
 sg13g2_decap_8 FILLER_170_1713 ();
 sg13g2_decap_8 FILLER_170_1720 ();
 sg13g2_decap_8 FILLER_170_1727 ();
 sg13g2_decap_8 FILLER_170_1734 ();
 sg13g2_decap_8 FILLER_170_1741 ();
 sg13g2_decap_8 FILLER_170_1748 ();
 sg13g2_decap_8 FILLER_170_1755 ();
 sg13g2_decap_4 FILLER_170_1762 ();
 sg13g2_fill_2 FILLER_170_1766 ();
 sg13g2_decap_8 FILLER_171_0 ();
 sg13g2_decap_8 FILLER_171_7 ();
 sg13g2_decap_8 FILLER_171_14 ();
 sg13g2_decap_8 FILLER_171_21 ();
 sg13g2_decap_8 FILLER_171_28 ();
 sg13g2_decap_8 FILLER_171_35 ();
 sg13g2_decap_8 FILLER_171_42 ();
 sg13g2_decap_8 FILLER_171_49 ();
 sg13g2_decap_8 FILLER_171_56 ();
 sg13g2_decap_8 FILLER_171_63 ();
 sg13g2_decap_8 FILLER_171_70 ();
 sg13g2_decap_8 FILLER_171_77 ();
 sg13g2_decap_8 FILLER_171_84 ();
 sg13g2_decap_8 FILLER_171_91 ();
 sg13g2_decap_8 FILLER_171_98 ();
 sg13g2_decap_8 FILLER_171_105 ();
 sg13g2_decap_8 FILLER_171_112 ();
 sg13g2_decap_8 FILLER_171_119 ();
 sg13g2_decap_8 FILLER_171_126 ();
 sg13g2_decap_8 FILLER_171_133 ();
 sg13g2_decap_8 FILLER_171_140 ();
 sg13g2_decap_8 FILLER_171_147 ();
 sg13g2_decap_8 FILLER_171_154 ();
 sg13g2_decap_8 FILLER_171_161 ();
 sg13g2_decap_8 FILLER_171_168 ();
 sg13g2_decap_8 FILLER_171_175 ();
 sg13g2_decap_8 FILLER_171_182 ();
 sg13g2_decap_8 FILLER_171_189 ();
 sg13g2_fill_2 FILLER_171_196 ();
 sg13g2_decap_4 FILLER_171_203 ();
 sg13g2_fill_1 FILLER_171_207 ();
 sg13g2_decap_4 FILLER_171_219 ();
 sg13g2_decap_8 FILLER_171_234 ();
 sg13g2_decap_8 FILLER_171_241 ();
 sg13g2_decap_8 FILLER_171_248 ();
 sg13g2_fill_2 FILLER_171_255 ();
 sg13g2_fill_1 FILLER_171_257 ();
 sg13g2_decap_4 FILLER_171_294 ();
 sg13g2_decap_8 FILLER_171_303 ();
 sg13g2_fill_2 FILLER_171_310 ();
 sg13g2_decap_8 FILLER_171_334 ();
 sg13g2_decap_8 FILLER_171_341 ();
 sg13g2_decap_8 FILLER_171_348 ();
 sg13g2_decap_8 FILLER_171_355 ();
 sg13g2_decap_8 FILLER_171_362 ();
 sg13g2_decap_8 FILLER_171_369 ();
 sg13g2_decap_8 FILLER_171_376 ();
 sg13g2_decap_8 FILLER_171_383 ();
 sg13g2_decap_8 FILLER_171_390 ();
 sg13g2_decap_8 FILLER_171_397 ();
 sg13g2_fill_2 FILLER_171_404 ();
 sg13g2_fill_1 FILLER_171_414 ();
 sg13g2_decap_8 FILLER_171_423 ();
 sg13g2_decap_8 FILLER_171_430 ();
 sg13g2_decap_4 FILLER_171_437 ();
 sg13g2_fill_1 FILLER_171_441 ();
 sg13g2_decap_8 FILLER_171_446 ();
 sg13g2_decap_8 FILLER_171_453 ();
 sg13g2_decap_8 FILLER_171_460 ();
 sg13g2_decap_8 FILLER_171_467 ();
 sg13g2_decap_8 FILLER_171_474 ();
 sg13g2_decap_8 FILLER_171_481 ();
 sg13g2_decap_8 FILLER_171_488 ();
 sg13g2_decap_8 FILLER_171_495 ();
 sg13g2_decap_8 FILLER_171_502 ();
 sg13g2_decap_8 FILLER_171_509 ();
 sg13g2_fill_2 FILLER_171_516 ();
 sg13g2_fill_2 FILLER_171_526 ();
 sg13g2_decap_8 FILLER_171_532 ();
 sg13g2_decap_4 FILLER_171_539 ();
 sg13g2_fill_1 FILLER_171_543 ();
 sg13g2_decap_8 FILLER_171_549 ();
 sg13g2_decap_8 FILLER_171_556 ();
 sg13g2_decap_8 FILLER_171_563 ();
 sg13g2_decap_4 FILLER_171_570 ();
 sg13g2_fill_2 FILLER_171_574 ();
 sg13g2_fill_2 FILLER_171_580 ();
 sg13g2_fill_1 FILLER_171_587 ();
 sg13g2_decap_8 FILLER_171_604 ();
 sg13g2_decap_8 FILLER_171_611 ();
 sg13g2_decap_8 FILLER_171_618 ();
 sg13g2_decap_8 FILLER_171_625 ();
 sg13g2_decap_8 FILLER_171_632 ();
 sg13g2_decap_8 FILLER_171_639 ();
 sg13g2_decap_8 FILLER_171_646 ();
 sg13g2_decap_8 FILLER_171_653 ();
 sg13g2_decap_8 FILLER_171_660 ();
 sg13g2_decap_8 FILLER_171_667 ();
 sg13g2_decap_8 FILLER_171_674 ();
 sg13g2_decap_8 FILLER_171_681 ();
 sg13g2_decap_4 FILLER_171_688 ();
 sg13g2_fill_1 FILLER_171_692 ();
 sg13g2_decap_8 FILLER_171_697 ();
 sg13g2_decap_8 FILLER_171_704 ();
 sg13g2_decap_8 FILLER_171_711 ();
 sg13g2_decap_8 FILLER_171_718 ();
 sg13g2_decap_8 FILLER_171_725 ();
 sg13g2_decap_8 FILLER_171_732 ();
 sg13g2_decap_8 FILLER_171_739 ();
 sg13g2_decap_8 FILLER_171_746 ();
 sg13g2_decap_8 FILLER_171_753 ();
 sg13g2_decap_8 FILLER_171_760 ();
 sg13g2_decap_4 FILLER_171_767 ();
 sg13g2_fill_2 FILLER_171_771 ();
 sg13g2_decap_8 FILLER_171_789 ();
 sg13g2_decap_8 FILLER_171_796 ();
 sg13g2_decap_4 FILLER_171_803 ();
 sg13g2_decap_8 FILLER_171_815 ();
 sg13g2_decap_8 FILLER_171_822 ();
 sg13g2_decap_8 FILLER_171_829 ();
 sg13g2_decap_4 FILLER_171_836 ();
 sg13g2_fill_1 FILLER_171_840 ();
 sg13g2_decap_8 FILLER_171_849 ();
 sg13g2_decap_8 FILLER_171_856 ();
 sg13g2_decap_8 FILLER_171_863 ();
 sg13g2_decap_4 FILLER_171_870 ();
 sg13g2_fill_2 FILLER_171_874 ();
 sg13g2_decap_8 FILLER_171_894 ();
 sg13g2_decap_8 FILLER_171_901 ();
 sg13g2_decap_8 FILLER_171_908 ();
 sg13g2_decap_8 FILLER_171_915 ();
 sg13g2_decap_8 FILLER_171_922 ();
 sg13g2_decap_8 FILLER_171_929 ();
 sg13g2_decap_8 FILLER_171_936 ();
 sg13g2_decap_8 FILLER_171_943 ();
 sg13g2_decap_8 FILLER_171_950 ();
 sg13g2_decap_8 FILLER_171_957 ();
 sg13g2_decap_8 FILLER_171_992 ();
 sg13g2_decap_8 FILLER_171_999 ();
 sg13g2_fill_2 FILLER_171_1006 ();
 sg13g2_fill_1 FILLER_171_1008 ();
 sg13g2_decap_8 FILLER_171_1018 ();
 sg13g2_fill_2 FILLER_171_1025 ();
 sg13g2_fill_2 FILLER_171_1031 ();
 sg13g2_fill_1 FILLER_171_1033 ();
 sg13g2_fill_2 FILLER_171_1038 ();
 sg13g2_decap_8 FILLER_171_1045 ();
 sg13g2_decap_8 FILLER_171_1052 ();
 sg13g2_decap_8 FILLER_171_1059 ();
 sg13g2_decap_8 FILLER_171_1066 ();
 sg13g2_decap_8 FILLER_171_1073 ();
 sg13g2_decap_8 FILLER_171_1080 ();
 sg13g2_decap_8 FILLER_171_1087 ();
 sg13g2_decap_8 FILLER_171_1094 ();
 sg13g2_decap_8 FILLER_171_1101 ();
 sg13g2_decap_8 FILLER_171_1108 ();
 sg13g2_decap_8 FILLER_171_1115 ();
 sg13g2_fill_2 FILLER_171_1122 ();
 sg13g2_decap_8 FILLER_171_1157 ();
 sg13g2_decap_8 FILLER_171_1164 ();
 sg13g2_decap_8 FILLER_171_1171 ();
 sg13g2_fill_1 FILLER_171_1191 ();
 sg13g2_decap_8 FILLER_171_1209 ();
 sg13g2_decap_8 FILLER_171_1216 ();
 sg13g2_decap_8 FILLER_171_1223 ();
 sg13g2_decap_8 FILLER_171_1230 ();
 sg13g2_decap_8 FILLER_171_1237 ();
 sg13g2_decap_8 FILLER_171_1244 ();
 sg13g2_decap_8 FILLER_171_1251 ();
 sg13g2_decap_8 FILLER_171_1258 ();
 sg13g2_decap_8 FILLER_171_1265 ();
 sg13g2_decap_8 FILLER_171_1272 ();
 sg13g2_decap_8 FILLER_171_1279 ();
 sg13g2_decap_8 FILLER_171_1286 ();
 sg13g2_decap_8 FILLER_171_1293 ();
 sg13g2_decap_8 FILLER_171_1300 ();
 sg13g2_decap_8 FILLER_171_1307 ();
 sg13g2_decap_8 FILLER_171_1314 ();
 sg13g2_decap_8 FILLER_171_1321 ();
 sg13g2_decap_8 FILLER_171_1328 ();
 sg13g2_decap_8 FILLER_171_1335 ();
 sg13g2_decap_8 FILLER_171_1342 ();
 sg13g2_decap_8 FILLER_171_1349 ();
 sg13g2_decap_8 FILLER_171_1356 ();
 sg13g2_decap_8 FILLER_171_1363 ();
 sg13g2_decap_8 FILLER_171_1370 ();
 sg13g2_decap_8 FILLER_171_1377 ();
 sg13g2_decap_8 FILLER_171_1384 ();
 sg13g2_decap_8 FILLER_171_1391 ();
 sg13g2_decap_8 FILLER_171_1398 ();
 sg13g2_decap_8 FILLER_171_1405 ();
 sg13g2_decap_8 FILLER_171_1412 ();
 sg13g2_decap_8 FILLER_171_1419 ();
 sg13g2_decap_8 FILLER_171_1426 ();
 sg13g2_decap_8 FILLER_171_1433 ();
 sg13g2_decap_8 FILLER_171_1440 ();
 sg13g2_decap_8 FILLER_171_1447 ();
 sg13g2_decap_8 FILLER_171_1454 ();
 sg13g2_decap_8 FILLER_171_1461 ();
 sg13g2_decap_8 FILLER_171_1468 ();
 sg13g2_decap_8 FILLER_171_1475 ();
 sg13g2_decap_8 FILLER_171_1482 ();
 sg13g2_decap_8 FILLER_171_1489 ();
 sg13g2_decap_8 FILLER_171_1496 ();
 sg13g2_decap_8 FILLER_171_1503 ();
 sg13g2_decap_8 FILLER_171_1510 ();
 sg13g2_decap_8 FILLER_171_1517 ();
 sg13g2_decap_8 FILLER_171_1524 ();
 sg13g2_decap_8 FILLER_171_1531 ();
 sg13g2_decap_8 FILLER_171_1538 ();
 sg13g2_decap_8 FILLER_171_1545 ();
 sg13g2_decap_8 FILLER_171_1552 ();
 sg13g2_decap_8 FILLER_171_1559 ();
 sg13g2_decap_8 FILLER_171_1566 ();
 sg13g2_decap_8 FILLER_171_1573 ();
 sg13g2_decap_8 FILLER_171_1580 ();
 sg13g2_decap_8 FILLER_171_1587 ();
 sg13g2_decap_8 FILLER_171_1594 ();
 sg13g2_decap_8 FILLER_171_1601 ();
 sg13g2_decap_8 FILLER_171_1608 ();
 sg13g2_decap_8 FILLER_171_1615 ();
 sg13g2_decap_8 FILLER_171_1622 ();
 sg13g2_decap_8 FILLER_171_1629 ();
 sg13g2_decap_8 FILLER_171_1636 ();
 sg13g2_decap_8 FILLER_171_1643 ();
 sg13g2_decap_8 FILLER_171_1650 ();
 sg13g2_decap_8 FILLER_171_1657 ();
 sg13g2_decap_8 FILLER_171_1664 ();
 sg13g2_decap_8 FILLER_171_1671 ();
 sg13g2_decap_8 FILLER_171_1678 ();
 sg13g2_decap_8 FILLER_171_1685 ();
 sg13g2_decap_8 FILLER_171_1692 ();
 sg13g2_decap_8 FILLER_171_1699 ();
 sg13g2_decap_8 FILLER_171_1706 ();
 sg13g2_decap_8 FILLER_171_1713 ();
 sg13g2_decap_8 FILLER_171_1720 ();
 sg13g2_decap_8 FILLER_171_1727 ();
 sg13g2_decap_8 FILLER_171_1734 ();
 sg13g2_decap_8 FILLER_171_1741 ();
 sg13g2_decap_8 FILLER_171_1748 ();
 sg13g2_decap_8 FILLER_171_1755 ();
 sg13g2_decap_4 FILLER_171_1762 ();
 sg13g2_fill_2 FILLER_171_1766 ();
 sg13g2_decap_8 FILLER_172_0 ();
 sg13g2_decap_8 FILLER_172_7 ();
 sg13g2_decap_8 FILLER_172_14 ();
 sg13g2_decap_8 FILLER_172_21 ();
 sg13g2_decap_8 FILLER_172_28 ();
 sg13g2_decap_8 FILLER_172_35 ();
 sg13g2_decap_8 FILLER_172_42 ();
 sg13g2_decap_8 FILLER_172_49 ();
 sg13g2_decap_8 FILLER_172_56 ();
 sg13g2_decap_8 FILLER_172_63 ();
 sg13g2_decap_8 FILLER_172_70 ();
 sg13g2_decap_8 FILLER_172_77 ();
 sg13g2_decap_8 FILLER_172_84 ();
 sg13g2_decap_8 FILLER_172_91 ();
 sg13g2_decap_8 FILLER_172_98 ();
 sg13g2_decap_8 FILLER_172_105 ();
 sg13g2_decap_8 FILLER_172_112 ();
 sg13g2_decap_8 FILLER_172_119 ();
 sg13g2_decap_8 FILLER_172_126 ();
 sg13g2_decap_8 FILLER_172_133 ();
 sg13g2_decap_8 FILLER_172_140 ();
 sg13g2_decap_8 FILLER_172_147 ();
 sg13g2_decap_8 FILLER_172_154 ();
 sg13g2_decap_8 FILLER_172_161 ();
 sg13g2_decap_8 FILLER_172_168 ();
 sg13g2_decap_8 FILLER_172_175 ();
 sg13g2_fill_2 FILLER_172_182 ();
 sg13g2_decap_4 FILLER_172_189 ();
 sg13g2_fill_1 FILLER_172_193 ();
 sg13g2_decap_8 FILLER_172_199 ();
 sg13g2_decap_8 FILLER_172_206 ();
 sg13g2_decap_8 FILLER_172_213 ();
 sg13g2_decap_8 FILLER_172_220 ();
 sg13g2_decap_8 FILLER_172_227 ();
 sg13g2_decap_8 FILLER_172_234 ();
 sg13g2_decap_8 FILLER_172_241 ();
 sg13g2_decap_8 FILLER_172_248 ();
 sg13g2_decap_8 FILLER_172_255 ();
 sg13g2_decap_4 FILLER_172_262 ();
 sg13g2_fill_2 FILLER_172_266 ();
 sg13g2_decap_4 FILLER_172_279 ();
 sg13g2_decap_8 FILLER_172_288 ();
 sg13g2_decap_8 FILLER_172_295 ();
 sg13g2_decap_8 FILLER_172_302 ();
 sg13g2_decap_4 FILLER_172_309 ();
 sg13g2_fill_1 FILLER_172_318 ();
 sg13g2_decap_8 FILLER_172_330 ();
 sg13g2_decap_8 FILLER_172_337 ();
 sg13g2_decap_8 FILLER_172_344 ();
 sg13g2_decap_8 FILLER_172_351 ();
 sg13g2_decap_4 FILLER_172_358 ();
 sg13g2_fill_1 FILLER_172_362 ();
 sg13g2_decap_8 FILLER_172_389 ();
 sg13g2_decap_8 FILLER_172_396 ();
 sg13g2_decap_8 FILLER_172_403 ();
 sg13g2_decap_4 FILLER_172_410 ();
 sg13g2_fill_2 FILLER_172_414 ();
 sg13g2_decap_8 FILLER_172_420 ();
 sg13g2_decap_8 FILLER_172_427 ();
 sg13g2_fill_2 FILLER_172_434 ();
 sg13g2_fill_1 FILLER_172_448 ();
 sg13g2_decap_8 FILLER_172_454 ();
 sg13g2_decap_8 FILLER_172_461 ();
 sg13g2_decap_4 FILLER_172_468 ();
 sg13g2_fill_2 FILLER_172_472 ();
 sg13g2_decap_8 FILLER_172_495 ();
 sg13g2_decap_8 FILLER_172_502 ();
 sg13g2_decap_8 FILLER_172_509 ();
 sg13g2_decap_8 FILLER_172_516 ();
 sg13g2_decap_8 FILLER_172_523 ();
 sg13g2_fill_1 FILLER_172_539 ();
 sg13g2_decap_8 FILLER_172_560 ();
 sg13g2_decap_8 FILLER_172_567 ();
 sg13g2_decap_8 FILLER_172_574 ();
 sg13g2_fill_2 FILLER_172_581 ();
 sg13g2_decap_8 FILLER_172_599 ();
 sg13g2_decap_8 FILLER_172_606 ();
 sg13g2_decap_8 FILLER_172_613 ();
 sg13g2_decap_8 FILLER_172_620 ();
 sg13g2_decap_8 FILLER_172_627 ();
 sg13g2_decap_8 FILLER_172_634 ();
 sg13g2_decap_8 FILLER_172_641 ();
 sg13g2_decap_8 FILLER_172_648 ();
 sg13g2_decap_8 FILLER_172_655 ();
 sg13g2_decap_8 FILLER_172_662 ();
 sg13g2_decap_8 FILLER_172_669 ();
 sg13g2_decap_8 FILLER_172_676 ();
 sg13g2_decap_8 FILLER_172_683 ();
 sg13g2_decap_8 FILLER_172_690 ();
 sg13g2_decap_8 FILLER_172_697 ();
 sg13g2_decap_8 FILLER_172_704 ();
 sg13g2_decap_8 FILLER_172_711 ();
 sg13g2_decap_8 FILLER_172_718 ();
 sg13g2_decap_8 FILLER_172_725 ();
 sg13g2_decap_8 FILLER_172_732 ();
 sg13g2_decap_8 FILLER_172_739 ();
 sg13g2_decap_8 FILLER_172_746 ();
 sg13g2_decap_8 FILLER_172_753 ();
 sg13g2_decap_8 FILLER_172_760 ();
 sg13g2_decap_4 FILLER_172_767 ();
 sg13g2_fill_2 FILLER_172_771 ();
 sg13g2_decap_8 FILLER_172_781 ();
 sg13g2_decap_8 FILLER_172_788 ();
 sg13g2_decap_8 FILLER_172_795 ();
 sg13g2_decap_8 FILLER_172_802 ();
 sg13g2_decap_8 FILLER_172_809 ();
 sg13g2_decap_8 FILLER_172_816 ();
 sg13g2_decap_8 FILLER_172_823 ();
 sg13g2_decap_8 FILLER_172_830 ();
 sg13g2_decap_8 FILLER_172_837 ();
 sg13g2_decap_8 FILLER_172_844 ();
 sg13g2_decap_8 FILLER_172_851 ();
 sg13g2_decap_8 FILLER_172_858 ();
 sg13g2_decap_8 FILLER_172_865 ();
 sg13g2_decap_8 FILLER_172_872 ();
 sg13g2_decap_8 FILLER_172_879 ();
 sg13g2_decap_8 FILLER_172_886 ();
 sg13g2_decap_4 FILLER_172_893 ();
 sg13g2_fill_1 FILLER_172_897 ();
 sg13g2_decap_8 FILLER_172_921 ();
 sg13g2_decap_8 FILLER_172_928 ();
 sg13g2_decap_8 FILLER_172_935 ();
 sg13g2_decap_8 FILLER_172_942 ();
 sg13g2_decap_8 FILLER_172_949 ();
 sg13g2_decap_8 FILLER_172_956 ();
 sg13g2_decap_8 FILLER_172_963 ();
 sg13g2_decap_8 FILLER_172_970 ();
 sg13g2_decap_8 FILLER_172_977 ();
 sg13g2_decap_8 FILLER_172_984 ();
 sg13g2_decap_8 FILLER_172_991 ();
 sg13g2_decap_8 FILLER_172_998 ();
 sg13g2_decap_8 FILLER_172_1005 ();
 sg13g2_decap_4 FILLER_172_1012 ();
 sg13g2_fill_1 FILLER_172_1016 ();
 sg13g2_decap_8 FILLER_172_1025 ();
 sg13g2_decap_4 FILLER_172_1032 ();
 sg13g2_fill_2 FILLER_172_1036 ();
 sg13g2_decap_8 FILLER_172_1050 ();
 sg13g2_decap_8 FILLER_172_1057 ();
 sg13g2_decap_8 FILLER_172_1064 ();
 sg13g2_fill_1 FILLER_172_1071 ();
 sg13g2_decap_8 FILLER_172_1083 ();
 sg13g2_decap_8 FILLER_172_1090 ();
 sg13g2_decap_8 FILLER_172_1097 ();
 sg13g2_decap_8 FILLER_172_1104 ();
 sg13g2_decap_8 FILLER_172_1111 ();
 sg13g2_decap_8 FILLER_172_1118 ();
 sg13g2_decap_8 FILLER_172_1125 ();
 sg13g2_fill_2 FILLER_172_1132 ();
 sg13g2_decap_8 FILLER_172_1152 ();
 sg13g2_decap_8 FILLER_172_1159 ();
 sg13g2_decap_8 FILLER_172_1166 ();
 sg13g2_decap_8 FILLER_172_1177 ();
 sg13g2_decap_4 FILLER_172_1184 ();
 sg13g2_fill_1 FILLER_172_1188 ();
 sg13g2_decap_8 FILLER_172_1201 ();
 sg13g2_decap_8 FILLER_172_1208 ();
 sg13g2_decap_8 FILLER_172_1215 ();
 sg13g2_decap_8 FILLER_172_1222 ();
 sg13g2_decap_8 FILLER_172_1229 ();
 sg13g2_decap_8 FILLER_172_1236 ();
 sg13g2_decap_8 FILLER_172_1243 ();
 sg13g2_decap_8 FILLER_172_1250 ();
 sg13g2_decap_8 FILLER_172_1257 ();
 sg13g2_decap_8 FILLER_172_1264 ();
 sg13g2_decap_8 FILLER_172_1271 ();
 sg13g2_decap_8 FILLER_172_1278 ();
 sg13g2_decap_8 FILLER_172_1285 ();
 sg13g2_decap_8 FILLER_172_1292 ();
 sg13g2_decap_8 FILLER_172_1299 ();
 sg13g2_decap_8 FILLER_172_1306 ();
 sg13g2_decap_8 FILLER_172_1313 ();
 sg13g2_decap_8 FILLER_172_1320 ();
 sg13g2_decap_8 FILLER_172_1327 ();
 sg13g2_decap_8 FILLER_172_1334 ();
 sg13g2_decap_8 FILLER_172_1341 ();
 sg13g2_decap_8 FILLER_172_1348 ();
 sg13g2_decap_8 FILLER_172_1355 ();
 sg13g2_decap_8 FILLER_172_1362 ();
 sg13g2_decap_8 FILLER_172_1369 ();
 sg13g2_decap_8 FILLER_172_1376 ();
 sg13g2_decap_8 FILLER_172_1383 ();
 sg13g2_decap_8 FILLER_172_1390 ();
 sg13g2_decap_8 FILLER_172_1397 ();
 sg13g2_decap_8 FILLER_172_1404 ();
 sg13g2_decap_8 FILLER_172_1411 ();
 sg13g2_decap_8 FILLER_172_1418 ();
 sg13g2_decap_8 FILLER_172_1425 ();
 sg13g2_decap_8 FILLER_172_1432 ();
 sg13g2_decap_8 FILLER_172_1439 ();
 sg13g2_decap_8 FILLER_172_1446 ();
 sg13g2_decap_8 FILLER_172_1453 ();
 sg13g2_decap_8 FILLER_172_1460 ();
 sg13g2_decap_8 FILLER_172_1467 ();
 sg13g2_decap_8 FILLER_172_1474 ();
 sg13g2_decap_8 FILLER_172_1481 ();
 sg13g2_decap_8 FILLER_172_1488 ();
 sg13g2_decap_8 FILLER_172_1495 ();
 sg13g2_decap_8 FILLER_172_1502 ();
 sg13g2_decap_8 FILLER_172_1509 ();
 sg13g2_decap_8 FILLER_172_1516 ();
 sg13g2_decap_8 FILLER_172_1523 ();
 sg13g2_decap_8 FILLER_172_1530 ();
 sg13g2_decap_8 FILLER_172_1537 ();
 sg13g2_decap_8 FILLER_172_1544 ();
 sg13g2_decap_8 FILLER_172_1551 ();
 sg13g2_decap_8 FILLER_172_1558 ();
 sg13g2_decap_8 FILLER_172_1565 ();
 sg13g2_decap_8 FILLER_172_1572 ();
 sg13g2_decap_8 FILLER_172_1579 ();
 sg13g2_decap_8 FILLER_172_1586 ();
 sg13g2_decap_8 FILLER_172_1593 ();
 sg13g2_decap_8 FILLER_172_1600 ();
 sg13g2_decap_8 FILLER_172_1607 ();
 sg13g2_decap_8 FILLER_172_1614 ();
 sg13g2_decap_8 FILLER_172_1621 ();
 sg13g2_decap_8 FILLER_172_1628 ();
 sg13g2_decap_8 FILLER_172_1635 ();
 sg13g2_decap_8 FILLER_172_1642 ();
 sg13g2_decap_8 FILLER_172_1649 ();
 sg13g2_decap_8 FILLER_172_1656 ();
 sg13g2_decap_8 FILLER_172_1663 ();
 sg13g2_decap_8 FILLER_172_1670 ();
 sg13g2_decap_8 FILLER_172_1677 ();
 sg13g2_decap_8 FILLER_172_1684 ();
 sg13g2_decap_8 FILLER_172_1691 ();
 sg13g2_decap_8 FILLER_172_1698 ();
 sg13g2_decap_8 FILLER_172_1705 ();
 sg13g2_decap_8 FILLER_172_1712 ();
 sg13g2_decap_8 FILLER_172_1719 ();
 sg13g2_decap_8 FILLER_172_1726 ();
 sg13g2_decap_8 FILLER_172_1733 ();
 sg13g2_decap_8 FILLER_172_1740 ();
 sg13g2_decap_8 FILLER_172_1747 ();
 sg13g2_decap_8 FILLER_172_1754 ();
 sg13g2_decap_8 FILLER_172_1761 ();
 sg13g2_decap_8 FILLER_173_0 ();
 sg13g2_decap_8 FILLER_173_7 ();
 sg13g2_decap_8 FILLER_173_14 ();
 sg13g2_decap_8 FILLER_173_21 ();
 sg13g2_decap_8 FILLER_173_28 ();
 sg13g2_decap_8 FILLER_173_35 ();
 sg13g2_decap_8 FILLER_173_42 ();
 sg13g2_decap_8 FILLER_173_49 ();
 sg13g2_decap_8 FILLER_173_56 ();
 sg13g2_decap_8 FILLER_173_63 ();
 sg13g2_decap_8 FILLER_173_70 ();
 sg13g2_decap_8 FILLER_173_77 ();
 sg13g2_decap_8 FILLER_173_84 ();
 sg13g2_decap_8 FILLER_173_91 ();
 sg13g2_decap_8 FILLER_173_98 ();
 sg13g2_decap_8 FILLER_173_105 ();
 sg13g2_decap_8 FILLER_173_112 ();
 sg13g2_decap_8 FILLER_173_119 ();
 sg13g2_decap_8 FILLER_173_126 ();
 sg13g2_decap_8 FILLER_173_133 ();
 sg13g2_decap_8 FILLER_173_140 ();
 sg13g2_decap_8 FILLER_173_147 ();
 sg13g2_decap_4 FILLER_173_154 ();
 sg13g2_fill_2 FILLER_173_158 ();
 sg13g2_decap_8 FILLER_173_164 ();
 sg13g2_decap_8 FILLER_173_171 ();
 sg13g2_decap_8 FILLER_173_178 ();
 sg13g2_decap_8 FILLER_173_185 ();
 sg13g2_decap_8 FILLER_173_192 ();
 sg13g2_fill_2 FILLER_173_199 ();
 sg13g2_fill_2 FILLER_173_212 ();
 sg13g2_decap_8 FILLER_173_220 ();
 sg13g2_decap_8 FILLER_173_227 ();
 sg13g2_decap_4 FILLER_173_234 ();
 sg13g2_fill_2 FILLER_173_238 ();
 sg13g2_decap_8 FILLER_173_245 ();
 sg13g2_decap_8 FILLER_173_252 ();
 sg13g2_decap_8 FILLER_173_264 ();
 sg13g2_decap_8 FILLER_173_271 ();
 sg13g2_decap_8 FILLER_173_278 ();
 sg13g2_decap_8 FILLER_173_285 ();
 sg13g2_decap_8 FILLER_173_292 ();
 sg13g2_decap_8 FILLER_173_299 ();
 sg13g2_decap_8 FILLER_173_306 ();
 sg13g2_decap_8 FILLER_173_313 ();
 sg13g2_decap_8 FILLER_173_320 ();
 sg13g2_decap_8 FILLER_173_327 ();
 sg13g2_decap_8 FILLER_173_334 ();
 sg13g2_decap_8 FILLER_173_341 ();
 sg13g2_decap_8 FILLER_173_348 ();
 sg13g2_decap_8 FILLER_173_355 ();
 sg13g2_fill_2 FILLER_173_362 ();
 sg13g2_decap_8 FILLER_173_395 ();
 sg13g2_decap_8 FILLER_173_402 ();
 sg13g2_decap_8 FILLER_173_409 ();
 sg13g2_decap_8 FILLER_173_416 ();
 sg13g2_decap_8 FILLER_173_423 ();
 sg13g2_decap_8 FILLER_173_430 ();
 sg13g2_decap_4 FILLER_173_437 ();
 sg13g2_decap_8 FILLER_173_449 ();
 sg13g2_decap_8 FILLER_173_456 ();
 sg13g2_decap_4 FILLER_173_463 ();
 sg13g2_fill_1 FILLER_173_467 ();
 sg13g2_decap_8 FILLER_173_481 ();
 sg13g2_decap_8 FILLER_173_488 ();
 sg13g2_decap_8 FILLER_173_495 ();
 sg13g2_decap_8 FILLER_173_502 ();
 sg13g2_fill_2 FILLER_173_509 ();
 sg13g2_decap_4 FILLER_173_516 ();
 sg13g2_decap_8 FILLER_173_528 ();
 sg13g2_decap_8 FILLER_173_535 ();
 sg13g2_fill_1 FILLER_173_542 ();
 sg13g2_decap_8 FILLER_173_551 ();
 sg13g2_decap_8 FILLER_173_558 ();
 sg13g2_decap_8 FILLER_173_565 ();
 sg13g2_decap_8 FILLER_173_572 ();
 sg13g2_decap_8 FILLER_173_579 ();
 sg13g2_decap_8 FILLER_173_586 ();
 sg13g2_decap_8 FILLER_173_593 ();
 sg13g2_decap_8 FILLER_173_600 ();
 sg13g2_decap_8 FILLER_173_607 ();
 sg13g2_decap_8 FILLER_173_614 ();
 sg13g2_decap_8 FILLER_173_621 ();
 sg13g2_decap_8 FILLER_173_628 ();
 sg13g2_decap_8 FILLER_173_635 ();
 sg13g2_decap_8 FILLER_173_642 ();
 sg13g2_decap_8 FILLER_173_649 ();
 sg13g2_decap_8 FILLER_173_656 ();
 sg13g2_decap_8 FILLER_173_663 ();
 sg13g2_decap_8 FILLER_173_670 ();
 sg13g2_fill_2 FILLER_173_681 ();
 sg13g2_fill_1 FILLER_173_683 ();
 sg13g2_decap_8 FILLER_173_689 ();
 sg13g2_decap_8 FILLER_173_696 ();
 sg13g2_decap_8 FILLER_173_703 ();
 sg13g2_decap_8 FILLER_173_710 ();
 sg13g2_decap_8 FILLER_173_717 ();
 sg13g2_decap_8 FILLER_173_735 ();
 sg13g2_decap_8 FILLER_173_742 ();
 sg13g2_decap_8 FILLER_173_765 ();
 sg13g2_decap_8 FILLER_173_772 ();
 sg13g2_decap_8 FILLER_173_779 ();
 sg13g2_decap_8 FILLER_173_786 ();
 sg13g2_decap_8 FILLER_173_793 ();
 sg13g2_decap_8 FILLER_173_800 ();
 sg13g2_decap_8 FILLER_173_807 ();
 sg13g2_decap_8 FILLER_173_814 ();
 sg13g2_decap_8 FILLER_173_821 ();
 sg13g2_fill_1 FILLER_173_828 ();
 sg13g2_decap_8 FILLER_173_834 ();
 sg13g2_decap_8 FILLER_173_841 ();
 sg13g2_decap_8 FILLER_173_848 ();
 sg13g2_decap_8 FILLER_173_855 ();
 sg13g2_decap_8 FILLER_173_862 ();
 sg13g2_decap_8 FILLER_173_869 ();
 sg13g2_decap_8 FILLER_173_876 ();
 sg13g2_decap_8 FILLER_173_883 ();
 sg13g2_fill_2 FILLER_173_890 ();
 sg13g2_fill_1 FILLER_173_892 ();
 sg13g2_decap_8 FILLER_173_917 ();
 sg13g2_decap_8 FILLER_173_924 ();
 sg13g2_decap_8 FILLER_173_931 ();
 sg13g2_decap_8 FILLER_173_938 ();
 sg13g2_decap_8 FILLER_173_945 ();
 sg13g2_decap_8 FILLER_173_952 ();
 sg13g2_decap_8 FILLER_173_959 ();
 sg13g2_decap_4 FILLER_173_966 ();
 sg13g2_fill_1 FILLER_173_970 ();
 sg13g2_decap_8 FILLER_173_974 ();
 sg13g2_decap_8 FILLER_173_981 ();
 sg13g2_decap_8 FILLER_173_988 ();
 sg13g2_decap_8 FILLER_173_995 ();
 sg13g2_decap_8 FILLER_173_1002 ();
 sg13g2_decap_8 FILLER_173_1009 ();
 sg13g2_fill_1 FILLER_173_1016 ();
 sg13g2_decap_8 FILLER_173_1038 ();
 sg13g2_decap_8 FILLER_173_1045 ();
 sg13g2_decap_8 FILLER_173_1052 ();
 sg13g2_decap_8 FILLER_173_1059 ();
 sg13g2_decap_8 FILLER_173_1066 ();
 sg13g2_decap_8 FILLER_173_1073 ();
 sg13g2_decap_8 FILLER_173_1080 ();
 sg13g2_decap_8 FILLER_173_1087 ();
 sg13g2_decap_8 FILLER_173_1094 ();
 sg13g2_decap_8 FILLER_173_1101 ();
 sg13g2_decap_8 FILLER_173_1108 ();
 sg13g2_decap_8 FILLER_173_1115 ();
 sg13g2_decap_4 FILLER_173_1122 ();
 sg13g2_fill_2 FILLER_173_1126 ();
 sg13g2_decap_8 FILLER_173_1153 ();
 sg13g2_decap_8 FILLER_173_1160 ();
 sg13g2_decap_8 FILLER_173_1167 ();
 sg13g2_decap_4 FILLER_173_1174 ();
 sg13g2_fill_2 FILLER_173_1178 ();
 sg13g2_decap_8 FILLER_173_1184 ();
 sg13g2_decap_8 FILLER_173_1191 ();
 sg13g2_decap_8 FILLER_173_1198 ();
 sg13g2_decap_8 FILLER_173_1205 ();
 sg13g2_decap_8 FILLER_173_1212 ();
 sg13g2_decap_8 FILLER_173_1219 ();
 sg13g2_decap_8 FILLER_173_1226 ();
 sg13g2_decap_8 FILLER_173_1233 ();
 sg13g2_decap_8 FILLER_173_1240 ();
 sg13g2_decap_8 FILLER_173_1247 ();
 sg13g2_decap_8 FILLER_173_1254 ();
 sg13g2_decap_8 FILLER_173_1261 ();
 sg13g2_decap_8 FILLER_173_1268 ();
 sg13g2_decap_8 FILLER_173_1275 ();
 sg13g2_decap_8 FILLER_173_1282 ();
 sg13g2_decap_8 FILLER_173_1289 ();
 sg13g2_decap_8 FILLER_173_1296 ();
 sg13g2_decap_8 FILLER_173_1303 ();
 sg13g2_decap_8 FILLER_173_1310 ();
 sg13g2_decap_8 FILLER_173_1317 ();
 sg13g2_decap_8 FILLER_173_1324 ();
 sg13g2_decap_8 FILLER_173_1331 ();
 sg13g2_decap_8 FILLER_173_1338 ();
 sg13g2_decap_8 FILLER_173_1345 ();
 sg13g2_decap_8 FILLER_173_1352 ();
 sg13g2_decap_8 FILLER_173_1359 ();
 sg13g2_decap_8 FILLER_173_1366 ();
 sg13g2_decap_8 FILLER_173_1373 ();
 sg13g2_decap_8 FILLER_173_1380 ();
 sg13g2_decap_8 FILLER_173_1387 ();
 sg13g2_decap_8 FILLER_173_1394 ();
 sg13g2_decap_8 FILLER_173_1401 ();
 sg13g2_decap_8 FILLER_173_1408 ();
 sg13g2_decap_8 FILLER_173_1415 ();
 sg13g2_decap_8 FILLER_173_1422 ();
 sg13g2_decap_8 FILLER_173_1429 ();
 sg13g2_decap_8 FILLER_173_1436 ();
 sg13g2_decap_8 FILLER_173_1443 ();
 sg13g2_decap_8 FILLER_173_1450 ();
 sg13g2_decap_8 FILLER_173_1457 ();
 sg13g2_decap_8 FILLER_173_1464 ();
 sg13g2_decap_8 FILLER_173_1471 ();
 sg13g2_decap_8 FILLER_173_1478 ();
 sg13g2_decap_8 FILLER_173_1485 ();
 sg13g2_decap_8 FILLER_173_1492 ();
 sg13g2_decap_8 FILLER_173_1499 ();
 sg13g2_decap_8 FILLER_173_1506 ();
 sg13g2_decap_8 FILLER_173_1513 ();
 sg13g2_decap_8 FILLER_173_1520 ();
 sg13g2_decap_8 FILLER_173_1527 ();
 sg13g2_decap_8 FILLER_173_1534 ();
 sg13g2_decap_8 FILLER_173_1541 ();
 sg13g2_decap_8 FILLER_173_1548 ();
 sg13g2_decap_8 FILLER_173_1555 ();
 sg13g2_decap_8 FILLER_173_1562 ();
 sg13g2_decap_8 FILLER_173_1569 ();
 sg13g2_decap_8 FILLER_173_1576 ();
 sg13g2_decap_8 FILLER_173_1583 ();
 sg13g2_decap_8 FILLER_173_1590 ();
 sg13g2_decap_8 FILLER_173_1597 ();
 sg13g2_decap_8 FILLER_173_1604 ();
 sg13g2_decap_8 FILLER_173_1611 ();
 sg13g2_decap_8 FILLER_173_1618 ();
 sg13g2_decap_8 FILLER_173_1625 ();
 sg13g2_decap_8 FILLER_173_1632 ();
 sg13g2_decap_8 FILLER_173_1639 ();
 sg13g2_decap_8 FILLER_173_1646 ();
 sg13g2_decap_8 FILLER_173_1653 ();
 sg13g2_decap_8 FILLER_173_1660 ();
 sg13g2_decap_8 FILLER_173_1667 ();
 sg13g2_decap_8 FILLER_173_1674 ();
 sg13g2_decap_8 FILLER_173_1681 ();
 sg13g2_decap_8 FILLER_173_1688 ();
 sg13g2_decap_8 FILLER_173_1695 ();
 sg13g2_decap_8 FILLER_173_1702 ();
 sg13g2_decap_8 FILLER_173_1709 ();
 sg13g2_decap_8 FILLER_173_1716 ();
 sg13g2_decap_8 FILLER_173_1723 ();
 sg13g2_decap_8 FILLER_173_1730 ();
 sg13g2_decap_8 FILLER_173_1737 ();
 sg13g2_decap_8 FILLER_173_1744 ();
 sg13g2_decap_8 FILLER_173_1751 ();
 sg13g2_decap_8 FILLER_173_1758 ();
 sg13g2_fill_2 FILLER_173_1765 ();
 sg13g2_fill_1 FILLER_173_1767 ();
 sg13g2_decap_8 FILLER_174_0 ();
 sg13g2_decap_8 FILLER_174_7 ();
 sg13g2_decap_8 FILLER_174_14 ();
 sg13g2_decap_8 FILLER_174_21 ();
 sg13g2_decap_8 FILLER_174_28 ();
 sg13g2_decap_8 FILLER_174_35 ();
 sg13g2_decap_8 FILLER_174_42 ();
 sg13g2_decap_8 FILLER_174_49 ();
 sg13g2_decap_8 FILLER_174_56 ();
 sg13g2_decap_8 FILLER_174_63 ();
 sg13g2_decap_8 FILLER_174_70 ();
 sg13g2_decap_8 FILLER_174_77 ();
 sg13g2_decap_8 FILLER_174_84 ();
 sg13g2_decap_8 FILLER_174_91 ();
 sg13g2_decap_8 FILLER_174_98 ();
 sg13g2_decap_8 FILLER_174_105 ();
 sg13g2_decap_8 FILLER_174_112 ();
 sg13g2_decap_8 FILLER_174_119 ();
 sg13g2_decap_8 FILLER_174_126 ();
 sg13g2_decap_8 FILLER_174_133 ();
 sg13g2_decap_8 FILLER_174_140 ();
 sg13g2_decap_8 FILLER_174_147 ();
 sg13g2_decap_8 FILLER_174_154 ();
 sg13g2_decap_8 FILLER_174_161 ();
 sg13g2_decap_8 FILLER_174_168 ();
 sg13g2_fill_2 FILLER_174_175 ();
 sg13g2_fill_1 FILLER_174_177 ();
 sg13g2_fill_2 FILLER_174_198 ();
 sg13g2_decap_4 FILLER_174_216 ();
 sg13g2_decap_8 FILLER_174_223 ();
 sg13g2_fill_1 FILLER_174_230 ();
 sg13g2_fill_2 FILLER_174_243 ();
 sg13g2_decap_8 FILLER_174_255 ();
 sg13g2_decap_4 FILLER_174_262 ();
 sg13g2_fill_1 FILLER_174_266 ();
 sg13g2_decap_8 FILLER_174_271 ();
 sg13g2_decap_8 FILLER_174_278 ();
 sg13g2_decap_8 FILLER_174_285 ();
 sg13g2_decap_8 FILLER_174_292 ();
 sg13g2_decap_8 FILLER_174_299 ();
 sg13g2_decap_8 FILLER_174_306 ();
 sg13g2_decap_8 FILLER_174_313 ();
 sg13g2_decap_8 FILLER_174_320 ();
 sg13g2_decap_8 FILLER_174_327 ();
 sg13g2_decap_8 FILLER_174_334 ();
 sg13g2_decap_8 FILLER_174_341 ();
 sg13g2_decap_8 FILLER_174_348 ();
 sg13g2_decap_8 FILLER_174_355 ();
 sg13g2_fill_2 FILLER_174_362 ();
 sg13g2_fill_1 FILLER_174_368 ();
 sg13g2_fill_1 FILLER_174_387 ();
 sg13g2_decap_8 FILLER_174_397 ();
 sg13g2_decap_8 FILLER_174_404 ();
 sg13g2_decap_8 FILLER_174_411 ();
 sg13g2_decap_8 FILLER_174_418 ();
 sg13g2_decap_8 FILLER_174_425 ();
 sg13g2_decap_8 FILLER_174_432 ();
 sg13g2_decap_8 FILLER_174_439 ();
 sg13g2_decap_8 FILLER_174_446 ();
 sg13g2_decap_4 FILLER_174_453 ();
 sg13g2_fill_1 FILLER_174_457 ();
 sg13g2_decap_4 FILLER_174_462 ();
 sg13g2_fill_2 FILLER_174_466 ();
 sg13g2_decap_8 FILLER_174_475 ();
 sg13g2_decap_8 FILLER_174_482 ();
 sg13g2_decap_8 FILLER_174_489 ();
 sg13g2_decap_8 FILLER_174_496 ();
 sg13g2_decap_4 FILLER_174_503 ();
 sg13g2_decap_8 FILLER_174_522 ();
 sg13g2_decap_8 FILLER_174_529 ();
 sg13g2_decap_8 FILLER_174_536 ();
 sg13g2_fill_2 FILLER_174_543 ();
 sg13g2_decap_8 FILLER_174_562 ();
 sg13g2_decap_8 FILLER_174_569 ();
 sg13g2_decap_8 FILLER_174_576 ();
 sg13g2_decap_8 FILLER_174_583 ();
 sg13g2_decap_8 FILLER_174_590 ();
 sg13g2_decap_8 FILLER_174_597 ();
 sg13g2_decap_4 FILLER_174_604 ();
 sg13g2_fill_2 FILLER_174_608 ();
 sg13g2_decap_8 FILLER_174_617 ();
 sg13g2_fill_1 FILLER_174_624 ();
 sg13g2_decap_8 FILLER_174_633 ();
 sg13g2_decap_8 FILLER_174_640 ();
 sg13g2_decap_8 FILLER_174_647 ();
 sg13g2_decap_8 FILLER_174_654 ();
 sg13g2_decap_8 FILLER_174_661 ();
 sg13g2_fill_1 FILLER_174_668 ();
 sg13g2_decap_8 FILLER_174_689 ();
 sg13g2_decap_8 FILLER_174_696 ();
 sg13g2_decap_8 FILLER_174_703 ();
 sg13g2_decap_8 FILLER_174_710 ();
 sg13g2_decap_4 FILLER_174_717 ();
 sg13g2_fill_1 FILLER_174_721 ();
 sg13g2_fill_2 FILLER_174_738 ();
 sg13g2_fill_1 FILLER_174_740 ();
 sg13g2_decap_8 FILLER_174_772 ();
 sg13g2_decap_8 FILLER_174_779 ();
 sg13g2_decap_8 FILLER_174_786 ();
 sg13g2_decap_8 FILLER_174_793 ();
 sg13g2_decap_8 FILLER_174_800 ();
 sg13g2_decap_8 FILLER_174_807 ();
 sg13g2_decap_4 FILLER_174_814 ();
 sg13g2_decap_4 FILLER_174_823 ();
 sg13g2_decap_8 FILLER_174_835 ();
 sg13g2_decap_8 FILLER_174_842 ();
 sg13g2_decap_8 FILLER_174_849 ();
 sg13g2_decap_8 FILLER_174_856 ();
 sg13g2_decap_8 FILLER_174_863 ();
 sg13g2_decap_8 FILLER_174_870 ();
 sg13g2_decap_8 FILLER_174_877 ();
 sg13g2_fill_2 FILLER_174_884 ();
 sg13g2_fill_1 FILLER_174_886 ();
 sg13g2_decap_8 FILLER_174_912 ();
 sg13g2_fill_2 FILLER_174_919 ();
 sg13g2_fill_1 FILLER_174_921 ();
 sg13g2_decap_8 FILLER_174_927 ();
 sg13g2_decap_8 FILLER_174_934 ();
 sg13g2_decap_8 FILLER_174_941 ();
 sg13g2_decap_8 FILLER_174_948 ();
 sg13g2_decap_8 FILLER_174_955 ();
 sg13g2_decap_4 FILLER_174_962 ();
 sg13g2_fill_1 FILLER_174_966 ();
 sg13g2_decap_8 FILLER_174_971 ();
 sg13g2_decap_8 FILLER_174_978 ();
 sg13g2_decap_8 FILLER_174_985 ();
 sg13g2_decap_8 FILLER_174_992 ();
 sg13g2_decap_8 FILLER_174_999 ();
 sg13g2_decap_8 FILLER_174_1006 ();
 sg13g2_fill_2 FILLER_174_1013 ();
 sg13g2_fill_1 FILLER_174_1015 ();
 sg13g2_fill_1 FILLER_174_1020 ();
 sg13g2_decap_8 FILLER_174_1025 ();
 sg13g2_decap_8 FILLER_174_1032 ();
 sg13g2_decap_8 FILLER_174_1039 ();
 sg13g2_fill_2 FILLER_174_1046 ();
 sg13g2_decap_8 FILLER_174_1051 ();
 sg13g2_decap_8 FILLER_174_1058 ();
 sg13g2_decap_8 FILLER_174_1065 ();
 sg13g2_decap_8 FILLER_174_1072 ();
 sg13g2_decap_8 FILLER_174_1079 ();
 sg13g2_decap_8 FILLER_174_1086 ();
 sg13g2_decap_8 FILLER_174_1093 ();
 sg13g2_decap_8 FILLER_174_1100 ();
 sg13g2_decap_4 FILLER_174_1107 ();
 sg13g2_fill_1 FILLER_174_1111 ();
 sg13g2_fill_2 FILLER_174_1117 ();
 sg13g2_decap_8 FILLER_174_1124 ();
 sg13g2_decap_4 FILLER_174_1131 ();
 sg13g2_fill_2 FILLER_174_1140 ();
 sg13g2_decap_8 FILLER_174_1146 ();
 sg13g2_decap_8 FILLER_174_1153 ();
 sg13g2_decap_8 FILLER_174_1160 ();
 sg13g2_fill_1 FILLER_174_1167 ();
 sg13g2_decap_8 FILLER_174_1176 ();
 sg13g2_decap_8 FILLER_174_1183 ();
 sg13g2_decap_8 FILLER_174_1190 ();
 sg13g2_decap_8 FILLER_174_1197 ();
 sg13g2_decap_8 FILLER_174_1204 ();
 sg13g2_decap_8 FILLER_174_1211 ();
 sg13g2_decap_8 FILLER_174_1218 ();
 sg13g2_decap_8 FILLER_174_1225 ();
 sg13g2_decap_8 FILLER_174_1232 ();
 sg13g2_decap_8 FILLER_174_1239 ();
 sg13g2_decap_8 FILLER_174_1246 ();
 sg13g2_decap_8 FILLER_174_1253 ();
 sg13g2_decap_8 FILLER_174_1260 ();
 sg13g2_decap_8 FILLER_174_1267 ();
 sg13g2_decap_8 FILLER_174_1274 ();
 sg13g2_decap_8 FILLER_174_1281 ();
 sg13g2_decap_8 FILLER_174_1288 ();
 sg13g2_decap_8 FILLER_174_1295 ();
 sg13g2_decap_8 FILLER_174_1302 ();
 sg13g2_decap_8 FILLER_174_1309 ();
 sg13g2_decap_8 FILLER_174_1316 ();
 sg13g2_decap_8 FILLER_174_1323 ();
 sg13g2_decap_8 FILLER_174_1330 ();
 sg13g2_decap_8 FILLER_174_1337 ();
 sg13g2_decap_8 FILLER_174_1344 ();
 sg13g2_decap_8 FILLER_174_1351 ();
 sg13g2_decap_8 FILLER_174_1358 ();
 sg13g2_decap_8 FILLER_174_1365 ();
 sg13g2_decap_8 FILLER_174_1372 ();
 sg13g2_decap_8 FILLER_174_1379 ();
 sg13g2_decap_8 FILLER_174_1386 ();
 sg13g2_decap_8 FILLER_174_1393 ();
 sg13g2_decap_8 FILLER_174_1400 ();
 sg13g2_decap_8 FILLER_174_1407 ();
 sg13g2_decap_8 FILLER_174_1414 ();
 sg13g2_decap_8 FILLER_174_1421 ();
 sg13g2_decap_8 FILLER_174_1428 ();
 sg13g2_decap_8 FILLER_174_1435 ();
 sg13g2_decap_8 FILLER_174_1442 ();
 sg13g2_decap_8 FILLER_174_1449 ();
 sg13g2_decap_8 FILLER_174_1456 ();
 sg13g2_decap_8 FILLER_174_1463 ();
 sg13g2_decap_8 FILLER_174_1470 ();
 sg13g2_decap_8 FILLER_174_1477 ();
 sg13g2_decap_8 FILLER_174_1484 ();
 sg13g2_decap_8 FILLER_174_1491 ();
 sg13g2_decap_8 FILLER_174_1498 ();
 sg13g2_decap_8 FILLER_174_1505 ();
 sg13g2_decap_8 FILLER_174_1512 ();
 sg13g2_decap_8 FILLER_174_1519 ();
 sg13g2_decap_8 FILLER_174_1526 ();
 sg13g2_decap_8 FILLER_174_1533 ();
 sg13g2_decap_8 FILLER_174_1540 ();
 sg13g2_decap_8 FILLER_174_1547 ();
 sg13g2_decap_8 FILLER_174_1554 ();
 sg13g2_decap_8 FILLER_174_1561 ();
 sg13g2_decap_8 FILLER_174_1568 ();
 sg13g2_decap_8 FILLER_174_1575 ();
 sg13g2_decap_8 FILLER_174_1582 ();
 sg13g2_decap_8 FILLER_174_1589 ();
 sg13g2_decap_8 FILLER_174_1596 ();
 sg13g2_decap_8 FILLER_174_1603 ();
 sg13g2_decap_8 FILLER_174_1610 ();
 sg13g2_decap_8 FILLER_174_1617 ();
 sg13g2_decap_8 FILLER_174_1624 ();
 sg13g2_decap_8 FILLER_174_1631 ();
 sg13g2_decap_8 FILLER_174_1638 ();
 sg13g2_decap_8 FILLER_174_1645 ();
 sg13g2_decap_8 FILLER_174_1652 ();
 sg13g2_decap_8 FILLER_174_1659 ();
 sg13g2_decap_8 FILLER_174_1666 ();
 sg13g2_decap_8 FILLER_174_1673 ();
 sg13g2_decap_8 FILLER_174_1680 ();
 sg13g2_decap_8 FILLER_174_1687 ();
 sg13g2_decap_8 FILLER_174_1694 ();
 sg13g2_decap_8 FILLER_174_1701 ();
 sg13g2_decap_8 FILLER_174_1708 ();
 sg13g2_decap_8 FILLER_174_1715 ();
 sg13g2_decap_8 FILLER_174_1722 ();
 sg13g2_decap_8 FILLER_174_1729 ();
 sg13g2_decap_8 FILLER_174_1736 ();
 sg13g2_decap_8 FILLER_174_1743 ();
 sg13g2_decap_8 FILLER_174_1750 ();
 sg13g2_decap_8 FILLER_174_1757 ();
 sg13g2_decap_4 FILLER_174_1764 ();
 sg13g2_decap_8 FILLER_175_0 ();
 sg13g2_decap_8 FILLER_175_7 ();
 sg13g2_decap_8 FILLER_175_14 ();
 sg13g2_decap_8 FILLER_175_21 ();
 sg13g2_decap_8 FILLER_175_28 ();
 sg13g2_decap_8 FILLER_175_35 ();
 sg13g2_decap_8 FILLER_175_42 ();
 sg13g2_decap_8 FILLER_175_49 ();
 sg13g2_decap_8 FILLER_175_56 ();
 sg13g2_decap_8 FILLER_175_63 ();
 sg13g2_decap_8 FILLER_175_70 ();
 sg13g2_decap_8 FILLER_175_77 ();
 sg13g2_decap_8 FILLER_175_84 ();
 sg13g2_decap_8 FILLER_175_91 ();
 sg13g2_decap_8 FILLER_175_98 ();
 sg13g2_decap_8 FILLER_175_105 ();
 sg13g2_decap_8 FILLER_175_112 ();
 sg13g2_decap_8 FILLER_175_119 ();
 sg13g2_decap_8 FILLER_175_126 ();
 sg13g2_decap_8 FILLER_175_133 ();
 sg13g2_decap_8 FILLER_175_140 ();
 sg13g2_decap_8 FILLER_175_147 ();
 sg13g2_decap_8 FILLER_175_154 ();
 sg13g2_decap_8 FILLER_175_161 ();
 sg13g2_decap_8 FILLER_175_168 ();
 sg13g2_decap_4 FILLER_175_175 ();
 sg13g2_fill_2 FILLER_175_187 ();
 sg13g2_fill_2 FILLER_175_200 ();
 sg13g2_fill_2 FILLER_175_226 ();
 sg13g2_decap_8 FILLER_175_234 ();
 sg13g2_decap_8 FILLER_175_241 ();
 sg13g2_decap_8 FILLER_175_248 ();
 sg13g2_decap_8 FILLER_175_255 ();
 sg13g2_fill_2 FILLER_175_262 ();
 sg13g2_decap_4 FILLER_175_269 ();
 sg13g2_fill_1 FILLER_175_273 ();
 sg13g2_fill_2 FILLER_175_277 ();
 sg13g2_decap_8 FILLER_175_289 ();
 sg13g2_decap_8 FILLER_175_296 ();
 sg13g2_decap_8 FILLER_175_303 ();
 sg13g2_decap_8 FILLER_175_310 ();
 sg13g2_decap_8 FILLER_175_317 ();
 sg13g2_decap_8 FILLER_175_324 ();
 sg13g2_decap_8 FILLER_175_331 ();
 sg13g2_decap_8 FILLER_175_338 ();
 sg13g2_decap_8 FILLER_175_345 ();
 sg13g2_decap_8 FILLER_175_352 ();
 sg13g2_decap_8 FILLER_175_359 ();
 sg13g2_decap_8 FILLER_175_366 ();
 sg13g2_decap_4 FILLER_175_373 ();
 sg13g2_fill_2 FILLER_175_377 ();
 sg13g2_decap_8 FILLER_175_387 ();
 sg13g2_decap_8 FILLER_175_394 ();
 sg13g2_decap_8 FILLER_175_401 ();
 sg13g2_decap_8 FILLER_175_408 ();
 sg13g2_decap_8 FILLER_175_415 ();
 sg13g2_decap_8 FILLER_175_422 ();
 sg13g2_decap_8 FILLER_175_429 ();
 sg13g2_decap_8 FILLER_175_436 ();
 sg13g2_fill_2 FILLER_175_443 ();
 sg13g2_fill_1 FILLER_175_445 ();
 sg13g2_decap_8 FILLER_175_479 ();
 sg13g2_decap_8 FILLER_175_486 ();
 sg13g2_decap_8 FILLER_175_493 ();
 sg13g2_decap_4 FILLER_175_500 ();
 sg13g2_fill_2 FILLER_175_504 ();
 sg13g2_decap_8 FILLER_175_515 ();
 sg13g2_decap_8 FILLER_175_522 ();
 sg13g2_decap_8 FILLER_175_529 ();
 sg13g2_decap_8 FILLER_175_536 ();
 sg13g2_decap_4 FILLER_175_543 ();
 sg13g2_decap_8 FILLER_175_559 ();
 sg13g2_decap_8 FILLER_175_566 ();
 sg13g2_decap_8 FILLER_175_573 ();
 sg13g2_decap_4 FILLER_175_580 ();
 sg13g2_fill_2 FILLER_175_589 ();
 sg13g2_fill_2 FILLER_175_598 ();
 sg13g2_fill_2 FILLER_175_617 ();
 sg13g2_fill_1 FILLER_175_619 ();
 sg13g2_decap_8 FILLER_175_630 ();
 sg13g2_decap_8 FILLER_175_637 ();
 sg13g2_decap_8 FILLER_175_644 ();
 sg13g2_decap_8 FILLER_175_651 ();
 sg13g2_fill_2 FILLER_175_658 ();
 sg13g2_decap_8 FILLER_175_694 ();
 sg13g2_decap_8 FILLER_175_701 ();
 sg13g2_decap_4 FILLER_175_708 ();
 sg13g2_fill_1 FILLER_175_712 ();
 sg13g2_decap_4 FILLER_175_741 ();
 sg13g2_fill_1 FILLER_175_745 ();
 sg13g2_fill_1 FILLER_175_756 ();
 sg13g2_decap_8 FILLER_175_775 ();
 sg13g2_decap_8 FILLER_175_782 ();
 sg13g2_decap_8 FILLER_175_789 ();
 sg13g2_decap_8 FILLER_175_796 ();
 sg13g2_decap_8 FILLER_175_803 ();
 sg13g2_fill_2 FILLER_175_826 ();
 sg13g2_fill_1 FILLER_175_828 ();
 sg13g2_decap_8 FILLER_175_841 ();
 sg13g2_decap_8 FILLER_175_848 ();
 sg13g2_decap_8 FILLER_175_855 ();
 sg13g2_decap_8 FILLER_175_862 ();
 sg13g2_decap_8 FILLER_175_869 ();
 sg13g2_decap_8 FILLER_175_876 ();
 sg13g2_decap_8 FILLER_175_901 ();
 sg13g2_decap_8 FILLER_175_908 ();
 sg13g2_decap_4 FILLER_175_915 ();
 sg13g2_decap_8 FILLER_175_925 ();
 sg13g2_decap_8 FILLER_175_932 ();
 sg13g2_decap_8 FILLER_175_939 ();
 sg13g2_decap_4 FILLER_175_946 ();
 sg13g2_fill_1 FILLER_175_950 ();
 sg13g2_decap_8 FILLER_175_986 ();
 sg13g2_decap_8 FILLER_175_993 ();
 sg13g2_decap_8 FILLER_175_1000 ();
 sg13g2_fill_2 FILLER_175_1007 ();
 sg13g2_fill_1 FILLER_175_1009 ();
 sg13g2_decap_8 FILLER_175_1018 ();
 sg13g2_decap_4 FILLER_175_1025 ();
 sg13g2_fill_1 FILLER_175_1029 ();
 sg13g2_decap_8 FILLER_175_1034 ();
 sg13g2_decap_8 FILLER_175_1041 ();
 sg13g2_decap_8 FILLER_175_1074 ();
 sg13g2_decap_8 FILLER_175_1081 ();
 sg13g2_decap_8 FILLER_175_1088 ();
 sg13g2_decap_8 FILLER_175_1095 ();
 sg13g2_fill_2 FILLER_175_1102 ();
 sg13g2_decap_8 FILLER_175_1136 ();
 sg13g2_decap_8 FILLER_175_1143 ();
 sg13g2_decap_8 FILLER_175_1150 ();
 sg13g2_decap_4 FILLER_175_1157 ();
 sg13g2_fill_1 FILLER_175_1161 ();
 sg13g2_decap_8 FILLER_175_1165 ();
 sg13g2_fill_1 FILLER_175_1172 ();
 sg13g2_decap_8 FILLER_175_1189 ();
 sg13g2_decap_8 FILLER_175_1196 ();
 sg13g2_decap_8 FILLER_175_1203 ();
 sg13g2_decap_8 FILLER_175_1210 ();
 sg13g2_decap_8 FILLER_175_1217 ();
 sg13g2_decap_8 FILLER_175_1224 ();
 sg13g2_decap_8 FILLER_175_1231 ();
 sg13g2_decap_8 FILLER_175_1238 ();
 sg13g2_decap_8 FILLER_175_1245 ();
 sg13g2_decap_8 FILLER_175_1252 ();
 sg13g2_decap_8 FILLER_175_1259 ();
 sg13g2_decap_8 FILLER_175_1266 ();
 sg13g2_decap_8 FILLER_175_1273 ();
 sg13g2_decap_8 FILLER_175_1280 ();
 sg13g2_decap_8 FILLER_175_1287 ();
 sg13g2_decap_8 FILLER_175_1294 ();
 sg13g2_decap_8 FILLER_175_1301 ();
 sg13g2_decap_8 FILLER_175_1308 ();
 sg13g2_decap_8 FILLER_175_1315 ();
 sg13g2_decap_8 FILLER_175_1322 ();
 sg13g2_decap_8 FILLER_175_1329 ();
 sg13g2_decap_8 FILLER_175_1336 ();
 sg13g2_decap_8 FILLER_175_1343 ();
 sg13g2_decap_8 FILLER_175_1350 ();
 sg13g2_decap_8 FILLER_175_1357 ();
 sg13g2_decap_8 FILLER_175_1364 ();
 sg13g2_decap_8 FILLER_175_1371 ();
 sg13g2_decap_8 FILLER_175_1378 ();
 sg13g2_decap_8 FILLER_175_1385 ();
 sg13g2_decap_8 FILLER_175_1392 ();
 sg13g2_decap_8 FILLER_175_1399 ();
 sg13g2_decap_8 FILLER_175_1406 ();
 sg13g2_decap_8 FILLER_175_1413 ();
 sg13g2_decap_8 FILLER_175_1420 ();
 sg13g2_decap_8 FILLER_175_1427 ();
 sg13g2_decap_8 FILLER_175_1434 ();
 sg13g2_decap_8 FILLER_175_1441 ();
 sg13g2_decap_8 FILLER_175_1448 ();
 sg13g2_decap_8 FILLER_175_1455 ();
 sg13g2_decap_8 FILLER_175_1462 ();
 sg13g2_decap_8 FILLER_175_1469 ();
 sg13g2_decap_8 FILLER_175_1476 ();
 sg13g2_decap_8 FILLER_175_1483 ();
 sg13g2_decap_8 FILLER_175_1490 ();
 sg13g2_decap_8 FILLER_175_1497 ();
 sg13g2_decap_8 FILLER_175_1504 ();
 sg13g2_decap_8 FILLER_175_1511 ();
 sg13g2_decap_8 FILLER_175_1518 ();
 sg13g2_decap_8 FILLER_175_1525 ();
 sg13g2_decap_8 FILLER_175_1532 ();
 sg13g2_decap_8 FILLER_175_1539 ();
 sg13g2_decap_8 FILLER_175_1546 ();
 sg13g2_decap_8 FILLER_175_1553 ();
 sg13g2_decap_8 FILLER_175_1560 ();
 sg13g2_decap_8 FILLER_175_1567 ();
 sg13g2_decap_8 FILLER_175_1574 ();
 sg13g2_decap_8 FILLER_175_1581 ();
 sg13g2_decap_8 FILLER_175_1588 ();
 sg13g2_decap_8 FILLER_175_1595 ();
 sg13g2_decap_8 FILLER_175_1602 ();
 sg13g2_decap_8 FILLER_175_1609 ();
 sg13g2_decap_8 FILLER_175_1616 ();
 sg13g2_decap_8 FILLER_175_1623 ();
 sg13g2_decap_8 FILLER_175_1630 ();
 sg13g2_decap_8 FILLER_175_1637 ();
 sg13g2_decap_8 FILLER_175_1644 ();
 sg13g2_decap_8 FILLER_175_1651 ();
 sg13g2_decap_8 FILLER_175_1658 ();
 sg13g2_decap_8 FILLER_175_1665 ();
 sg13g2_decap_8 FILLER_175_1672 ();
 sg13g2_decap_8 FILLER_175_1679 ();
 sg13g2_decap_8 FILLER_175_1686 ();
 sg13g2_decap_8 FILLER_175_1693 ();
 sg13g2_decap_8 FILLER_175_1700 ();
 sg13g2_decap_8 FILLER_175_1707 ();
 sg13g2_decap_8 FILLER_175_1714 ();
 sg13g2_decap_8 FILLER_175_1721 ();
 sg13g2_decap_8 FILLER_175_1728 ();
 sg13g2_decap_8 FILLER_175_1735 ();
 sg13g2_decap_8 FILLER_175_1742 ();
 sg13g2_decap_8 FILLER_175_1749 ();
 sg13g2_decap_8 FILLER_175_1756 ();
 sg13g2_decap_4 FILLER_175_1763 ();
 sg13g2_fill_1 FILLER_175_1767 ();
 sg13g2_decap_8 FILLER_176_0 ();
 sg13g2_decap_8 FILLER_176_7 ();
 sg13g2_decap_8 FILLER_176_14 ();
 sg13g2_decap_8 FILLER_176_21 ();
 sg13g2_decap_8 FILLER_176_28 ();
 sg13g2_decap_8 FILLER_176_35 ();
 sg13g2_decap_8 FILLER_176_42 ();
 sg13g2_decap_8 FILLER_176_49 ();
 sg13g2_decap_8 FILLER_176_56 ();
 sg13g2_decap_8 FILLER_176_63 ();
 sg13g2_decap_8 FILLER_176_70 ();
 sg13g2_decap_8 FILLER_176_77 ();
 sg13g2_decap_8 FILLER_176_84 ();
 sg13g2_decap_8 FILLER_176_91 ();
 sg13g2_decap_8 FILLER_176_98 ();
 sg13g2_decap_8 FILLER_176_105 ();
 sg13g2_decap_8 FILLER_176_112 ();
 sg13g2_decap_8 FILLER_176_119 ();
 sg13g2_decap_8 FILLER_176_126 ();
 sg13g2_decap_8 FILLER_176_133 ();
 sg13g2_decap_8 FILLER_176_140 ();
 sg13g2_decap_8 FILLER_176_147 ();
 sg13g2_decap_8 FILLER_176_154 ();
 sg13g2_decap_8 FILLER_176_161 ();
 sg13g2_decap_8 FILLER_176_168 ();
 sg13g2_decap_8 FILLER_176_175 ();
 sg13g2_fill_2 FILLER_176_182 ();
 sg13g2_fill_1 FILLER_176_204 ();
 sg13g2_decap_4 FILLER_176_216 ();
 sg13g2_decap_8 FILLER_176_226 ();
 sg13g2_decap_4 FILLER_176_249 ();
 sg13g2_fill_2 FILLER_176_253 ();
 sg13g2_decap_4 FILLER_176_259 ();
 sg13g2_decap_8 FILLER_176_298 ();
 sg13g2_decap_8 FILLER_176_305 ();
 sg13g2_decap_8 FILLER_176_312 ();
 sg13g2_decap_8 FILLER_176_319 ();
 sg13g2_decap_8 FILLER_176_341 ();
 sg13g2_decap_8 FILLER_176_352 ();
 sg13g2_decap_8 FILLER_176_359 ();
 sg13g2_decap_8 FILLER_176_366 ();
 sg13g2_decap_8 FILLER_176_373 ();
 sg13g2_decap_8 FILLER_176_380 ();
 sg13g2_decap_8 FILLER_176_387 ();
 sg13g2_fill_2 FILLER_176_394 ();
 sg13g2_fill_1 FILLER_176_396 ();
 sg13g2_decap_8 FILLER_176_410 ();
 sg13g2_decap_8 FILLER_176_417 ();
 sg13g2_decap_8 FILLER_176_424 ();
 sg13g2_decap_8 FILLER_176_431 ();
 sg13g2_decap_8 FILLER_176_484 ();
 sg13g2_decap_8 FILLER_176_491 ();
 sg13g2_decap_8 FILLER_176_498 ();
 sg13g2_decap_8 FILLER_176_518 ();
 sg13g2_decap_8 FILLER_176_525 ();
 sg13g2_decap_8 FILLER_176_532 ();
 sg13g2_decap_8 FILLER_176_539 ();
 sg13g2_decap_8 FILLER_176_546 ();
 sg13g2_decap_4 FILLER_176_553 ();
 sg13g2_fill_1 FILLER_176_557 ();
 sg13g2_decap_8 FILLER_176_562 ();
 sg13g2_decap_4 FILLER_176_569 ();
 sg13g2_fill_2 FILLER_176_573 ();
 sg13g2_fill_1 FILLER_176_591 ();
 sg13g2_fill_1 FILLER_176_612 ();
 sg13g2_decap_8 FILLER_176_638 ();
 sg13g2_decap_8 FILLER_176_645 ();
 sg13g2_decap_8 FILLER_176_652 ();
 sg13g2_decap_8 FILLER_176_659 ();
 sg13g2_decap_4 FILLER_176_666 ();
 sg13g2_fill_1 FILLER_176_670 ();
 sg13g2_decap_8 FILLER_176_684 ();
 sg13g2_decap_8 FILLER_176_691 ();
 sg13g2_decap_8 FILLER_176_698 ();
 sg13g2_decap_4 FILLER_176_705 ();
 sg13g2_fill_1 FILLER_176_709 ();
 sg13g2_fill_2 FILLER_176_721 ();
 sg13g2_fill_2 FILLER_176_727 ();
 sg13g2_decap_4 FILLER_176_737 ();
 sg13g2_fill_1 FILLER_176_741 ();
 sg13g2_decap_8 FILLER_176_784 ();
 sg13g2_decap_8 FILLER_176_791 ();
 sg13g2_decap_8 FILLER_176_798 ();
 sg13g2_decap_4 FILLER_176_805 ();
 sg13g2_fill_2 FILLER_176_809 ();
 sg13g2_decap_4 FILLER_176_816 ();
 sg13g2_decap_4 FILLER_176_825 ();
 sg13g2_fill_1 FILLER_176_829 ();
 sg13g2_decap_8 FILLER_176_833 ();
 sg13g2_fill_1 FILLER_176_840 ();
 sg13g2_decap_8 FILLER_176_846 ();
 sg13g2_decap_8 FILLER_176_853 ();
 sg13g2_decap_8 FILLER_176_860 ();
 sg13g2_decap_8 FILLER_176_867 ();
 sg13g2_decap_8 FILLER_176_874 ();
 sg13g2_decap_8 FILLER_176_881 ();
 sg13g2_decap_8 FILLER_176_888 ();
 sg13g2_decap_8 FILLER_176_895 ();
 sg13g2_decap_8 FILLER_176_902 ();
 sg13g2_decap_4 FILLER_176_909 ();
 sg13g2_decap_8 FILLER_176_929 ();
 sg13g2_decap_8 FILLER_176_936 ();
 sg13g2_decap_8 FILLER_176_943 ();
 sg13g2_decap_8 FILLER_176_950 ();
 sg13g2_decap_4 FILLER_176_957 ();
 sg13g2_fill_1 FILLER_176_966 ();
 sg13g2_decap_8 FILLER_176_998 ();
 sg13g2_decap_8 FILLER_176_1005 ();
 sg13g2_decap_8 FILLER_176_1012 ();
 sg13g2_fill_2 FILLER_176_1019 ();
 sg13g2_fill_1 FILLER_176_1021 ();
 sg13g2_fill_2 FILLER_176_1027 ();
 sg13g2_fill_2 FILLER_176_1037 ();
 sg13g2_fill_1 FILLER_176_1050 ();
 sg13g2_fill_2 FILLER_176_1090 ();
 sg13g2_fill_1 FILLER_176_1106 ();
 sg13g2_fill_1 FILLER_176_1119 ();
 sg13g2_decap_8 FILLER_176_1137 ();
 sg13g2_decap_8 FILLER_176_1144 ();
 sg13g2_decap_8 FILLER_176_1151 ();
 sg13g2_decap_8 FILLER_176_1158 ();
 sg13g2_decap_8 FILLER_176_1165 ();
 sg13g2_decap_8 FILLER_176_1172 ();
 sg13g2_decap_8 FILLER_176_1179 ();
 sg13g2_decap_8 FILLER_176_1186 ();
 sg13g2_decap_8 FILLER_176_1193 ();
 sg13g2_decap_8 FILLER_176_1200 ();
 sg13g2_decap_8 FILLER_176_1207 ();
 sg13g2_decap_8 FILLER_176_1214 ();
 sg13g2_decap_8 FILLER_176_1221 ();
 sg13g2_decap_8 FILLER_176_1228 ();
 sg13g2_decap_8 FILLER_176_1235 ();
 sg13g2_decap_8 FILLER_176_1242 ();
 sg13g2_decap_8 FILLER_176_1249 ();
 sg13g2_decap_8 FILLER_176_1256 ();
 sg13g2_decap_8 FILLER_176_1263 ();
 sg13g2_decap_8 FILLER_176_1270 ();
 sg13g2_decap_8 FILLER_176_1277 ();
 sg13g2_decap_8 FILLER_176_1284 ();
 sg13g2_decap_8 FILLER_176_1291 ();
 sg13g2_decap_8 FILLER_176_1298 ();
 sg13g2_decap_8 FILLER_176_1305 ();
 sg13g2_decap_8 FILLER_176_1312 ();
 sg13g2_decap_8 FILLER_176_1319 ();
 sg13g2_decap_8 FILLER_176_1326 ();
 sg13g2_decap_8 FILLER_176_1333 ();
 sg13g2_decap_8 FILLER_176_1340 ();
 sg13g2_decap_8 FILLER_176_1347 ();
 sg13g2_decap_8 FILLER_176_1354 ();
 sg13g2_decap_8 FILLER_176_1361 ();
 sg13g2_decap_8 FILLER_176_1368 ();
 sg13g2_decap_8 FILLER_176_1375 ();
 sg13g2_decap_8 FILLER_176_1382 ();
 sg13g2_decap_8 FILLER_176_1389 ();
 sg13g2_decap_8 FILLER_176_1396 ();
 sg13g2_decap_8 FILLER_176_1403 ();
 sg13g2_decap_8 FILLER_176_1410 ();
 sg13g2_decap_8 FILLER_176_1417 ();
 sg13g2_decap_8 FILLER_176_1424 ();
 sg13g2_decap_8 FILLER_176_1431 ();
 sg13g2_decap_8 FILLER_176_1438 ();
 sg13g2_decap_8 FILLER_176_1445 ();
 sg13g2_decap_8 FILLER_176_1452 ();
 sg13g2_decap_8 FILLER_176_1459 ();
 sg13g2_decap_8 FILLER_176_1466 ();
 sg13g2_decap_8 FILLER_176_1473 ();
 sg13g2_decap_8 FILLER_176_1480 ();
 sg13g2_decap_8 FILLER_176_1487 ();
 sg13g2_decap_8 FILLER_176_1494 ();
 sg13g2_decap_8 FILLER_176_1501 ();
 sg13g2_decap_8 FILLER_176_1508 ();
 sg13g2_decap_8 FILLER_176_1515 ();
 sg13g2_decap_8 FILLER_176_1522 ();
 sg13g2_decap_8 FILLER_176_1529 ();
 sg13g2_decap_8 FILLER_176_1536 ();
 sg13g2_decap_8 FILLER_176_1543 ();
 sg13g2_decap_8 FILLER_176_1550 ();
 sg13g2_decap_8 FILLER_176_1557 ();
 sg13g2_decap_8 FILLER_176_1564 ();
 sg13g2_decap_8 FILLER_176_1571 ();
 sg13g2_decap_8 FILLER_176_1578 ();
 sg13g2_decap_8 FILLER_176_1585 ();
 sg13g2_decap_8 FILLER_176_1592 ();
 sg13g2_decap_8 FILLER_176_1599 ();
 sg13g2_decap_8 FILLER_176_1606 ();
 sg13g2_decap_8 FILLER_176_1613 ();
 sg13g2_decap_8 FILLER_176_1620 ();
 sg13g2_decap_8 FILLER_176_1627 ();
 sg13g2_decap_8 FILLER_176_1634 ();
 sg13g2_decap_8 FILLER_176_1641 ();
 sg13g2_decap_8 FILLER_176_1648 ();
 sg13g2_decap_8 FILLER_176_1655 ();
 sg13g2_decap_8 FILLER_176_1662 ();
 sg13g2_decap_8 FILLER_176_1669 ();
 sg13g2_decap_8 FILLER_176_1676 ();
 sg13g2_decap_8 FILLER_176_1683 ();
 sg13g2_decap_8 FILLER_176_1690 ();
 sg13g2_decap_8 FILLER_176_1697 ();
 sg13g2_decap_8 FILLER_176_1704 ();
 sg13g2_decap_8 FILLER_176_1711 ();
 sg13g2_decap_8 FILLER_176_1718 ();
 sg13g2_decap_8 FILLER_176_1725 ();
 sg13g2_decap_8 FILLER_176_1732 ();
 sg13g2_decap_8 FILLER_176_1739 ();
 sg13g2_decap_8 FILLER_176_1746 ();
 sg13g2_decap_8 FILLER_176_1753 ();
 sg13g2_decap_8 FILLER_176_1760 ();
 sg13g2_fill_1 FILLER_176_1767 ();
 sg13g2_decap_8 FILLER_177_0 ();
 sg13g2_decap_8 FILLER_177_7 ();
 sg13g2_decap_8 FILLER_177_14 ();
 sg13g2_decap_8 FILLER_177_21 ();
 sg13g2_decap_8 FILLER_177_28 ();
 sg13g2_decap_8 FILLER_177_35 ();
 sg13g2_decap_8 FILLER_177_42 ();
 sg13g2_decap_8 FILLER_177_49 ();
 sg13g2_decap_8 FILLER_177_56 ();
 sg13g2_decap_8 FILLER_177_63 ();
 sg13g2_decap_8 FILLER_177_70 ();
 sg13g2_decap_8 FILLER_177_77 ();
 sg13g2_decap_8 FILLER_177_84 ();
 sg13g2_decap_8 FILLER_177_91 ();
 sg13g2_decap_8 FILLER_177_98 ();
 sg13g2_decap_8 FILLER_177_105 ();
 sg13g2_decap_8 FILLER_177_112 ();
 sg13g2_decap_8 FILLER_177_119 ();
 sg13g2_decap_8 FILLER_177_126 ();
 sg13g2_decap_8 FILLER_177_133 ();
 sg13g2_decap_8 FILLER_177_140 ();
 sg13g2_decap_8 FILLER_177_147 ();
 sg13g2_decap_8 FILLER_177_154 ();
 sg13g2_decap_8 FILLER_177_161 ();
 sg13g2_decap_8 FILLER_177_168 ();
 sg13g2_decap_8 FILLER_177_175 ();
 sg13g2_decap_8 FILLER_177_210 ();
 sg13g2_decap_8 FILLER_177_217 ();
 sg13g2_decap_8 FILLER_177_224 ();
 sg13g2_decap_8 FILLER_177_231 ();
 sg13g2_fill_2 FILLER_177_238 ();
 sg13g2_decap_8 FILLER_177_245 ();
 sg13g2_decap_4 FILLER_177_252 ();
 sg13g2_fill_1 FILLER_177_256 ();
 sg13g2_decap_8 FILLER_177_298 ();
 sg13g2_decap_8 FILLER_177_305 ();
 sg13g2_decap_8 FILLER_177_312 ();
 sg13g2_decap_4 FILLER_177_319 ();
 sg13g2_fill_2 FILLER_177_323 ();
 sg13g2_decap_8 FILLER_177_351 ();
 sg13g2_decap_8 FILLER_177_358 ();
 sg13g2_decap_4 FILLER_177_365 ();
 sg13g2_fill_2 FILLER_177_369 ();
 sg13g2_decap_8 FILLER_177_420 ();
 sg13g2_decap_8 FILLER_177_427 ();
 sg13g2_decap_8 FILLER_177_434 ();
 sg13g2_decap_8 FILLER_177_441 ();
 sg13g2_fill_2 FILLER_177_460 ();
 sg13g2_decap_8 FILLER_177_476 ();
 sg13g2_decap_8 FILLER_177_483 ();
 sg13g2_decap_8 FILLER_177_490 ();
 sg13g2_decap_4 FILLER_177_497 ();
 sg13g2_decap_8 FILLER_177_506 ();
 sg13g2_decap_8 FILLER_177_521 ();
 sg13g2_decap_8 FILLER_177_528 ();
 sg13g2_decap_8 FILLER_177_535 ();
 sg13g2_decap_8 FILLER_177_542 ();
 sg13g2_fill_2 FILLER_177_549 ();
 sg13g2_decap_4 FILLER_177_580 ();
 sg13g2_fill_1 FILLER_177_584 ();
 sg13g2_fill_2 FILLER_177_589 ();
 sg13g2_fill_1 FILLER_177_591 ();
 sg13g2_fill_2 FILLER_177_597 ();
 sg13g2_fill_1 FILLER_177_599 ();
 sg13g2_decap_4 FILLER_177_605 ();
 sg13g2_fill_2 FILLER_177_609 ();
 sg13g2_decap_8 FILLER_177_647 ();
 sg13g2_fill_2 FILLER_177_654 ();
 sg13g2_fill_1 FILLER_177_656 ();
 sg13g2_decap_4 FILLER_177_678 ();
 sg13g2_decap_8 FILLER_177_688 ();
 sg13g2_decap_8 FILLER_177_695 ();
 sg13g2_decap_8 FILLER_177_702 ();
 sg13g2_decap_4 FILLER_177_709 ();
 sg13g2_fill_1 FILLER_177_713 ();
 sg13g2_decap_8 FILLER_177_734 ();
 sg13g2_decap_8 FILLER_177_741 ();
 sg13g2_decap_8 FILLER_177_748 ();
 sg13g2_decap_8 FILLER_177_788 ();
 sg13g2_decap_8 FILLER_177_795 ();
 sg13g2_decap_4 FILLER_177_802 ();
 sg13g2_fill_2 FILLER_177_825 ();
 sg13g2_fill_1 FILLER_177_827 ();
 sg13g2_decap_4 FILLER_177_840 ();
 sg13g2_fill_1 FILLER_177_844 ();
 sg13g2_decap_8 FILLER_177_880 ();
 sg13g2_fill_2 FILLER_177_887 ();
 sg13g2_fill_1 FILLER_177_889 ();
 sg13g2_decap_8 FILLER_177_898 ();
 sg13g2_fill_1 FILLER_177_905 ();
 sg13g2_fill_2 FILLER_177_911 ();
 sg13g2_fill_1 FILLER_177_913 ();
 sg13g2_fill_2 FILLER_177_922 ();
 sg13g2_decap_4 FILLER_177_932 ();
 sg13g2_fill_2 FILLER_177_936 ();
 sg13g2_decap_8 FILLER_177_955 ();
 sg13g2_decap_4 FILLER_177_962 ();
 sg13g2_fill_2 FILLER_177_966 ();
 sg13g2_fill_1 FILLER_177_973 ();
 sg13g2_fill_2 FILLER_177_993 ();
 sg13g2_fill_1 FILLER_177_995 ();
 sg13g2_decap_8 FILLER_177_1011 ();
 sg13g2_decap_4 FILLER_177_1018 ();
 sg13g2_fill_2 FILLER_177_1022 ();
 sg13g2_decap_4 FILLER_177_1042 ();
 sg13g2_decap_8 FILLER_177_1071 ();
 sg13g2_decap_4 FILLER_177_1078 ();
 sg13g2_fill_2 FILLER_177_1082 ();
 sg13g2_decap_8 FILLER_177_1092 ();
 sg13g2_decap_8 FILLER_177_1099 ();
 sg13g2_decap_4 FILLER_177_1106 ();
 sg13g2_fill_1 FILLER_177_1115 ();
 sg13g2_decap_8 FILLER_177_1139 ();
 sg13g2_decap_8 FILLER_177_1146 ();
 sg13g2_decap_8 FILLER_177_1153 ();
 sg13g2_decap_8 FILLER_177_1160 ();
 sg13g2_decap_8 FILLER_177_1167 ();
 sg13g2_decap_8 FILLER_177_1174 ();
 sg13g2_decap_8 FILLER_177_1181 ();
 sg13g2_decap_8 FILLER_177_1188 ();
 sg13g2_decap_8 FILLER_177_1195 ();
 sg13g2_decap_8 FILLER_177_1202 ();
 sg13g2_decap_8 FILLER_177_1209 ();
 sg13g2_decap_8 FILLER_177_1216 ();
 sg13g2_decap_8 FILLER_177_1223 ();
 sg13g2_decap_8 FILLER_177_1230 ();
 sg13g2_decap_8 FILLER_177_1237 ();
 sg13g2_decap_8 FILLER_177_1244 ();
 sg13g2_decap_8 FILLER_177_1251 ();
 sg13g2_decap_8 FILLER_177_1258 ();
 sg13g2_decap_8 FILLER_177_1265 ();
 sg13g2_decap_8 FILLER_177_1272 ();
 sg13g2_decap_8 FILLER_177_1279 ();
 sg13g2_decap_8 FILLER_177_1286 ();
 sg13g2_decap_8 FILLER_177_1293 ();
 sg13g2_decap_8 FILLER_177_1300 ();
 sg13g2_decap_8 FILLER_177_1307 ();
 sg13g2_decap_8 FILLER_177_1314 ();
 sg13g2_decap_8 FILLER_177_1321 ();
 sg13g2_decap_8 FILLER_177_1328 ();
 sg13g2_decap_8 FILLER_177_1335 ();
 sg13g2_decap_8 FILLER_177_1342 ();
 sg13g2_decap_8 FILLER_177_1349 ();
 sg13g2_decap_8 FILLER_177_1356 ();
 sg13g2_decap_8 FILLER_177_1363 ();
 sg13g2_decap_8 FILLER_177_1370 ();
 sg13g2_decap_8 FILLER_177_1377 ();
 sg13g2_decap_8 FILLER_177_1384 ();
 sg13g2_decap_8 FILLER_177_1391 ();
 sg13g2_decap_8 FILLER_177_1398 ();
 sg13g2_decap_8 FILLER_177_1405 ();
 sg13g2_decap_8 FILLER_177_1412 ();
 sg13g2_decap_8 FILLER_177_1419 ();
 sg13g2_decap_8 FILLER_177_1426 ();
 sg13g2_decap_8 FILLER_177_1433 ();
 sg13g2_decap_8 FILLER_177_1440 ();
 sg13g2_decap_8 FILLER_177_1447 ();
 sg13g2_decap_8 FILLER_177_1454 ();
 sg13g2_decap_8 FILLER_177_1461 ();
 sg13g2_decap_8 FILLER_177_1468 ();
 sg13g2_decap_8 FILLER_177_1475 ();
 sg13g2_decap_8 FILLER_177_1482 ();
 sg13g2_decap_8 FILLER_177_1489 ();
 sg13g2_decap_8 FILLER_177_1496 ();
 sg13g2_decap_8 FILLER_177_1503 ();
 sg13g2_decap_8 FILLER_177_1510 ();
 sg13g2_decap_8 FILLER_177_1517 ();
 sg13g2_decap_8 FILLER_177_1524 ();
 sg13g2_decap_8 FILLER_177_1531 ();
 sg13g2_decap_8 FILLER_177_1538 ();
 sg13g2_decap_8 FILLER_177_1545 ();
 sg13g2_decap_8 FILLER_177_1552 ();
 sg13g2_decap_8 FILLER_177_1559 ();
 sg13g2_decap_8 FILLER_177_1566 ();
 sg13g2_decap_8 FILLER_177_1573 ();
 sg13g2_decap_8 FILLER_177_1580 ();
 sg13g2_decap_8 FILLER_177_1587 ();
 sg13g2_decap_8 FILLER_177_1594 ();
 sg13g2_decap_8 FILLER_177_1601 ();
 sg13g2_decap_8 FILLER_177_1608 ();
 sg13g2_decap_8 FILLER_177_1615 ();
 sg13g2_decap_8 FILLER_177_1622 ();
 sg13g2_decap_8 FILLER_177_1629 ();
 sg13g2_decap_8 FILLER_177_1636 ();
 sg13g2_decap_8 FILLER_177_1643 ();
 sg13g2_decap_8 FILLER_177_1650 ();
 sg13g2_decap_8 FILLER_177_1657 ();
 sg13g2_decap_8 FILLER_177_1664 ();
 sg13g2_decap_8 FILLER_177_1671 ();
 sg13g2_decap_8 FILLER_177_1678 ();
 sg13g2_decap_8 FILLER_177_1685 ();
 sg13g2_decap_8 FILLER_177_1692 ();
 sg13g2_decap_8 FILLER_177_1699 ();
 sg13g2_decap_8 FILLER_177_1706 ();
 sg13g2_decap_8 FILLER_177_1713 ();
 sg13g2_decap_8 FILLER_177_1720 ();
 sg13g2_decap_8 FILLER_177_1727 ();
 sg13g2_decap_8 FILLER_177_1734 ();
 sg13g2_decap_8 FILLER_177_1741 ();
 sg13g2_decap_8 FILLER_177_1748 ();
 sg13g2_decap_8 FILLER_177_1755 ();
 sg13g2_decap_4 FILLER_177_1762 ();
 sg13g2_fill_2 FILLER_177_1766 ();
 sg13g2_decap_8 FILLER_178_0 ();
 sg13g2_decap_8 FILLER_178_7 ();
 sg13g2_decap_8 FILLER_178_14 ();
 sg13g2_decap_8 FILLER_178_21 ();
 sg13g2_decap_8 FILLER_178_28 ();
 sg13g2_decap_8 FILLER_178_35 ();
 sg13g2_decap_8 FILLER_178_42 ();
 sg13g2_decap_8 FILLER_178_49 ();
 sg13g2_decap_8 FILLER_178_56 ();
 sg13g2_decap_8 FILLER_178_63 ();
 sg13g2_decap_8 FILLER_178_70 ();
 sg13g2_decap_8 FILLER_178_77 ();
 sg13g2_decap_8 FILLER_178_84 ();
 sg13g2_decap_8 FILLER_178_91 ();
 sg13g2_decap_8 FILLER_178_98 ();
 sg13g2_decap_8 FILLER_178_105 ();
 sg13g2_decap_8 FILLER_178_112 ();
 sg13g2_decap_8 FILLER_178_119 ();
 sg13g2_decap_8 FILLER_178_126 ();
 sg13g2_decap_8 FILLER_178_133 ();
 sg13g2_decap_8 FILLER_178_140 ();
 sg13g2_decap_8 FILLER_178_147 ();
 sg13g2_decap_8 FILLER_178_154 ();
 sg13g2_decap_8 FILLER_178_161 ();
 sg13g2_decap_8 FILLER_178_168 ();
 sg13g2_decap_8 FILLER_178_175 ();
 sg13g2_decap_8 FILLER_178_182 ();
 sg13g2_decap_8 FILLER_178_189 ();
 sg13g2_decap_4 FILLER_178_196 ();
 sg13g2_fill_2 FILLER_178_200 ();
 sg13g2_decap_4 FILLER_178_207 ();
 sg13g2_decap_8 FILLER_178_216 ();
 sg13g2_decap_8 FILLER_178_223 ();
 sg13g2_decap_8 FILLER_178_230 ();
 sg13g2_decap_8 FILLER_178_237 ();
 sg13g2_decap_8 FILLER_178_244 ();
 sg13g2_decap_8 FILLER_178_251 ();
 sg13g2_fill_2 FILLER_178_258 ();
 sg13g2_fill_1 FILLER_178_260 ();
 sg13g2_fill_1 FILLER_178_267 ();
 sg13g2_decap_8 FILLER_178_287 ();
 sg13g2_decap_8 FILLER_178_294 ();
 sg13g2_decap_8 FILLER_178_301 ();
 sg13g2_decap_8 FILLER_178_308 ();
 sg13g2_decap_8 FILLER_178_315 ();
 sg13g2_decap_8 FILLER_178_322 ();
 sg13g2_fill_2 FILLER_178_329 ();
 sg13g2_fill_1 FILLER_178_340 ();
 sg13g2_decap_4 FILLER_178_367 ();
 sg13g2_decap_8 FILLER_178_380 ();
 sg13g2_decap_4 FILLER_178_387 ();
 sg13g2_fill_1 FILLER_178_391 ();
 sg13g2_decap_8 FILLER_178_396 ();
 sg13g2_decap_4 FILLER_178_403 ();
 sg13g2_decap_8 FILLER_178_416 ();
 sg13g2_decap_8 FILLER_178_423 ();
 sg13g2_decap_8 FILLER_178_430 ();
 sg13g2_decap_8 FILLER_178_437 ();
 sg13g2_decap_8 FILLER_178_444 ();
 sg13g2_decap_8 FILLER_178_451 ();
 sg13g2_decap_8 FILLER_178_458 ();
 sg13g2_fill_2 FILLER_178_465 ();
 sg13g2_fill_1 FILLER_178_467 ();
 sg13g2_decap_8 FILLER_178_488 ();
 sg13g2_fill_1 FILLER_178_495 ();
 sg13g2_decap_8 FILLER_178_516 ();
 sg13g2_decap_8 FILLER_178_523 ();
 sg13g2_decap_8 FILLER_178_530 ();
 sg13g2_decap_8 FILLER_178_537 ();
 sg13g2_decap_8 FILLER_178_544 ();
 sg13g2_decap_8 FILLER_178_551 ();
 sg13g2_decap_8 FILLER_178_558 ();
 sg13g2_decap_8 FILLER_178_565 ();
 sg13g2_decap_4 FILLER_178_572 ();
 sg13g2_decap_4 FILLER_178_584 ();
 sg13g2_fill_1 FILLER_178_588 ();
 sg13g2_decap_8 FILLER_178_594 ();
 sg13g2_decap_8 FILLER_178_601 ();
 sg13g2_decap_8 FILLER_178_608 ();
 sg13g2_fill_2 FILLER_178_615 ();
 sg13g2_decap_4 FILLER_178_621 ();
 sg13g2_fill_2 FILLER_178_625 ();
 sg13g2_decap_8 FILLER_178_635 ();
 sg13g2_decap_8 FILLER_178_642 ();
 sg13g2_decap_8 FILLER_178_649 ();
 sg13g2_fill_1 FILLER_178_656 ();
 sg13g2_decap_8 FILLER_178_676 ();
 sg13g2_decap_8 FILLER_178_683 ();
 sg13g2_decap_4 FILLER_178_690 ();
 sg13g2_fill_1 FILLER_178_694 ();
 sg13g2_decap_8 FILLER_178_731 ();
 sg13g2_decap_8 FILLER_178_738 ();
 sg13g2_decap_8 FILLER_178_745 ();
 sg13g2_decap_8 FILLER_178_752 ();
 sg13g2_fill_2 FILLER_178_759 ();
 sg13g2_decap_8 FILLER_178_786 ();
 sg13g2_decap_8 FILLER_178_793 ();
 sg13g2_fill_1 FILLER_178_800 ();
 sg13g2_decap_8 FILLER_178_842 ();
 sg13g2_decap_8 FILLER_178_849 ();
 sg13g2_decap_8 FILLER_178_891 ();
 sg13g2_decap_8 FILLER_178_898 ();
 sg13g2_decap_8 FILLER_178_910 ();
 sg13g2_decap_8 FILLER_178_917 ();
 sg13g2_fill_2 FILLER_178_924 ();
 sg13g2_fill_1 FILLER_178_926 ();
 sg13g2_decap_8 FILLER_178_951 ();
 sg13g2_decap_8 FILLER_178_958 ();
 sg13g2_decap_8 FILLER_178_965 ();
 sg13g2_decap_8 FILLER_178_972 ();
 sg13g2_decap_4 FILLER_178_979 ();
 sg13g2_fill_1 FILLER_178_983 ();
 sg13g2_fill_1 FILLER_178_989 ();
 sg13g2_decap_8 FILLER_178_994 ();
 sg13g2_decap_8 FILLER_178_1001 ();
 sg13g2_decap_8 FILLER_178_1008 ();
 sg13g2_decap_8 FILLER_178_1015 ();
 sg13g2_decap_8 FILLER_178_1022 ();
 sg13g2_fill_1 FILLER_178_1029 ();
 sg13g2_decap_8 FILLER_178_1041 ();
 sg13g2_decap_8 FILLER_178_1048 ();
 sg13g2_decap_8 FILLER_178_1055 ();
 sg13g2_decap_8 FILLER_178_1062 ();
 sg13g2_decap_8 FILLER_178_1069 ();
 sg13g2_decap_8 FILLER_178_1076 ();
 sg13g2_decap_8 FILLER_178_1083 ();
 sg13g2_decap_8 FILLER_178_1090 ();
 sg13g2_decap_8 FILLER_178_1097 ();
 sg13g2_decap_8 FILLER_178_1104 ();
 sg13g2_decap_8 FILLER_178_1111 ();
 sg13g2_decap_8 FILLER_178_1118 ();
 sg13g2_decap_4 FILLER_178_1125 ();
 sg13g2_decap_8 FILLER_178_1133 ();
 sg13g2_decap_8 FILLER_178_1140 ();
 sg13g2_decap_8 FILLER_178_1147 ();
 sg13g2_decap_8 FILLER_178_1154 ();
 sg13g2_decap_8 FILLER_178_1161 ();
 sg13g2_decap_8 FILLER_178_1168 ();
 sg13g2_decap_8 FILLER_178_1175 ();
 sg13g2_decap_8 FILLER_178_1182 ();
 sg13g2_decap_8 FILLER_178_1189 ();
 sg13g2_decap_8 FILLER_178_1196 ();
 sg13g2_decap_8 FILLER_178_1203 ();
 sg13g2_decap_8 FILLER_178_1210 ();
 sg13g2_decap_8 FILLER_178_1217 ();
 sg13g2_decap_8 FILLER_178_1224 ();
 sg13g2_decap_8 FILLER_178_1231 ();
 sg13g2_decap_8 FILLER_178_1238 ();
 sg13g2_decap_8 FILLER_178_1245 ();
 sg13g2_decap_8 FILLER_178_1252 ();
 sg13g2_decap_8 FILLER_178_1259 ();
 sg13g2_decap_8 FILLER_178_1266 ();
 sg13g2_decap_8 FILLER_178_1273 ();
 sg13g2_decap_8 FILLER_178_1280 ();
 sg13g2_decap_8 FILLER_178_1287 ();
 sg13g2_decap_8 FILLER_178_1294 ();
 sg13g2_decap_8 FILLER_178_1301 ();
 sg13g2_decap_8 FILLER_178_1308 ();
 sg13g2_decap_8 FILLER_178_1315 ();
 sg13g2_decap_8 FILLER_178_1322 ();
 sg13g2_decap_8 FILLER_178_1329 ();
 sg13g2_decap_8 FILLER_178_1336 ();
 sg13g2_decap_8 FILLER_178_1343 ();
 sg13g2_decap_8 FILLER_178_1350 ();
 sg13g2_decap_8 FILLER_178_1357 ();
 sg13g2_decap_8 FILLER_178_1364 ();
 sg13g2_decap_8 FILLER_178_1371 ();
 sg13g2_decap_8 FILLER_178_1378 ();
 sg13g2_decap_8 FILLER_178_1385 ();
 sg13g2_decap_8 FILLER_178_1392 ();
 sg13g2_decap_8 FILLER_178_1399 ();
 sg13g2_decap_8 FILLER_178_1406 ();
 sg13g2_decap_8 FILLER_178_1413 ();
 sg13g2_decap_8 FILLER_178_1420 ();
 sg13g2_decap_8 FILLER_178_1427 ();
 sg13g2_decap_8 FILLER_178_1434 ();
 sg13g2_decap_8 FILLER_178_1441 ();
 sg13g2_decap_8 FILLER_178_1448 ();
 sg13g2_decap_8 FILLER_178_1455 ();
 sg13g2_decap_8 FILLER_178_1462 ();
 sg13g2_decap_8 FILLER_178_1469 ();
 sg13g2_decap_8 FILLER_178_1476 ();
 sg13g2_decap_8 FILLER_178_1483 ();
 sg13g2_decap_8 FILLER_178_1490 ();
 sg13g2_decap_8 FILLER_178_1497 ();
 sg13g2_decap_8 FILLER_178_1504 ();
 sg13g2_decap_8 FILLER_178_1511 ();
 sg13g2_decap_8 FILLER_178_1518 ();
 sg13g2_decap_8 FILLER_178_1525 ();
 sg13g2_decap_8 FILLER_178_1532 ();
 sg13g2_decap_8 FILLER_178_1539 ();
 sg13g2_decap_8 FILLER_178_1546 ();
 sg13g2_decap_8 FILLER_178_1553 ();
 sg13g2_decap_8 FILLER_178_1560 ();
 sg13g2_decap_8 FILLER_178_1567 ();
 sg13g2_decap_8 FILLER_178_1574 ();
 sg13g2_decap_8 FILLER_178_1581 ();
 sg13g2_decap_8 FILLER_178_1588 ();
 sg13g2_decap_8 FILLER_178_1595 ();
 sg13g2_decap_8 FILLER_178_1602 ();
 sg13g2_decap_8 FILLER_178_1609 ();
 sg13g2_decap_8 FILLER_178_1616 ();
 sg13g2_decap_8 FILLER_178_1623 ();
 sg13g2_decap_8 FILLER_178_1630 ();
 sg13g2_decap_8 FILLER_178_1637 ();
 sg13g2_decap_8 FILLER_178_1644 ();
 sg13g2_decap_8 FILLER_178_1651 ();
 sg13g2_decap_8 FILLER_178_1658 ();
 sg13g2_decap_8 FILLER_178_1665 ();
 sg13g2_decap_8 FILLER_178_1672 ();
 sg13g2_decap_8 FILLER_178_1679 ();
 sg13g2_decap_8 FILLER_178_1686 ();
 sg13g2_decap_8 FILLER_178_1693 ();
 sg13g2_decap_8 FILLER_178_1700 ();
 sg13g2_decap_8 FILLER_178_1707 ();
 sg13g2_decap_8 FILLER_178_1714 ();
 sg13g2_decap_8 FILLER_178_1721 ();
 sg13g2_decap_8 FILLER_178_1728 ();
 sg13g2_decap_8 FILLER_178_1735 ();
 sg13g2_decap_8 FILLER_178_1742 ();
 sg13g2_decap_8 FILLER_178_1749 ();
 sg13g2_decap_8 FILLER_178_1756 ();
 sg13g2_decap_4 FILLER_178_1763 ();
 sg13g2_fill_1 FILLER_178_1767 ();
 sg13g2_decap_8 FILLER_179_0 ();
 sg13g2_decap_8 FILLER_179_7 ();
 sg13g2_decap_8 FILLER_179_14 ();
 sg13g2_decap_8 FILLER_179_21 ();
 sg13g2_decap_8 FILLER_179_28 ();
 sg13g2_decap_8 FILLER_179_35 ();
 sg13g2_decap_8 FILLER_179_42 ();
 sg13g2_decap_8 FILLER_179_49 ();
 sg13g2_decap_8 FILLER_179_56 ();
 sg13g2_decap_8 FILLER_179_63 ();
 sg13g2_decap_8 FILLER_179_70 ();
 sg13g2_decap_8 FILLER_179_77 ();
 sg13g2_decap_8 FILLER_179_84 ();
 sg13g2_decap_8 FILLER_179_91 ();
 sg13g2_decap_8 FILLER_179_98 ();
 sg13g2_decap_8 FILLER_179_105 ();
 sg13g2_decap_8 FILLER_179_112 ();
 sg13g2_decap_8 FILLER_179_119 ();
 sg13g2_decap_8 FILLER_179_126 ();
 sg13g2_decap_8 FILLER_179_133 ();
 sg13g2_decap_8 FILLER_179_140 ();
 sg13g2_decap_8 FILLER_179_147 ();
 sg13g2_decap_8 FILLER_179_154 ();
 sg13g2_decap_8 FILLER_179_161 ();
 sg13g2_decap_8 FILLER_179_168 ();
 sg13g2_decap_8 FILLER_179_175 ();
 sg13g2_decap_8 FILLER_179_182 ();
 sg13g2_decap_8 FILLER_179_189 ();
 sg13g2_decap_8 FILLER_179_196 ();
 sg13g2_fill_2 FILLER_179_203 ();
 sg13g2_fill_1 FILLER_179_205 ();
 sg13g2_decap_8 FILLER_179_227 ();
 sg13g2_fill_2 FILLER_179_234 ();
 sg13g2_fill_1 FILLER_179_236 ();
 sg13g2_decap_8 FILLER_179_240 ();
 sg13g2_fill_2 FILLER_179_247 ();
 sg13g2_decap_8 FILLER_179_254 ();
 sg13g2_decap_8 FILLER_179_261 ();
 sg13g2_decap_8 FILLER_179_268 ();
 sg13g2_fill_2 FILLER_179_275 ();
 sg13g2_decap_8 FILLER_179_280 ();
 sg13g2_fill_2 FILLER_179_287 ();
 sg13g2_decap_8 FILLER_179_301 ();
 sg13g2_decap_8 FILLER_179_308 ();
 sg13g2_decap_8 FILLER_179_315 ();
 sg13g2_decap_8 FILLER_179_322 ();
 sg13g2_decap_4 FILLER_179_329 ();
 sg13g2_fill_2 FILLER_179_333 ();
 sg13g2_decap_4 FILLER_179_339 ();
 sg13g2_fill_1 FILLER_179_343 ();
 sg13g2_decap_4 FILLER_179_358 ();
 sg13g2_fill_1 FILLER_179_362 ();
 sg13g2_decap_8 FILLER_179_368 ();
 sg13g2_decap_8 FILLER_179_375 ();
 sg13g2_decap_8 FILLER_179_382 ();
 sg13g2_decap_8 FILLER_179_389 ();
 sg13g2_decap_8 FILLER_179_396 ();
 sg13g2_decap_8 FILLER_179_403 ();
 sg13g2_decap_8 FILLER_179_410 ();
 sg13g2_decap_8 FILLER_179_417 ();
 sg13g2_decap_8 FILLER_179_424 ();
 sg13g2_decap_8 FILLER_179_431 ();
 sg13g2_decap_8 FILLER_179_438 ();
 sg13g2_decap_8 FILLER_179_445 ();
 sg13g2_decap_8 FILLER_179_452 ();
 sg13g2_decap_8 FILLER_179_459 ();
 sg13g2_decap_8 FILLER_179_466 ();
 sg13g2_fill_1 FILLER_179_473 ();
 sg13g2_decap_8 FILLER_179_478 ();
 sg13g2_decap_8 FILLER_179_497 ();
 sg13g2_decap_8 FILLER_179_504 ();
 sg13g2_fill_2 FILLER_179_511 ();
 sg13g2_decap_8 FILLER_179_518 ();
 sg13g2_decap_8 FILLER_179_525 ();
 sg13g2_decap_8 FILLER_179_532 ();
 sg13g2_decap_8 FILLER_179_539 ();
 sg13g2_decap_4 FILLER_179_550 ();
 sg13g2_fill_2 FILLER_179_564 ();
 sg13g2_decap_8 FILLER_179_582 ();
 sg13g2_decap_8 FILLER_179_589 ();
 sg13g2_decap_8 FILLER_179_596 ();
 sg13g2_decap_8 FILLER_179_603 ();
 sg13g2_decap_8 FILLER_179_610 ();
 sg13g2_decap_8 FILLER_179_617 ();
 sg13g2_decap_8 FILLER_179_624 ();
 sg13g2_decap_8 FILLER_179_631 ();
 sg13g2_decap_8 FILLER_179_638 ();
 sg13g2_decap_4 FILLER_179_645 ();
 sg13g2_decap_8 FILLER_179_653 ();
 sg13g2_decap_4 FILLER_179_660 ();
 sg13g2_fill_2 FILLER_179_664 ();
 sg13g2_decap_8 FILLER_179_670 ();
 sg13g2_decap_8 FILLER_179_677 ();
 sg13g2_decap_4 FILLER_179_684 ();
 sg13g2_fill_2 FILLER_179_688 ();
 sg13g2_decap_8 FILLER_179_726 ();
 sg13g2_decap_8 FILLER_179_733 ();
 sg13g2_decap_8 FILLER_179_740 ();
 sg13g2_decap_8 FILLER_179_747 ();
 sg13g2_decap_8 FILLER_179_754 ();
 sg13g2_decap_8 FILLER_179_761 ();
 sg13g2_fill_2 FILLER_179_768 ();
 sg13g2_fill_1 FILLER_179_770 ();
 sg13g2_decap_8 FILLER_179_779 ();
 sg13g2_decap_8 FILLER_179_786 ();
 sg13g2_decap_8 FILLER_179_793 ();
 sg13g2_decap_8 FILLER_179_800 ();
 sg13g2_decap_4 FILLER_179_807 ();
 sg13g2_decap_8 FILLER_179_830 ();
 sg13g2_decap_8 FILLER_179_837 ();
 sg13g2_decap_8 FILLER_179_844 ();
 sg13g2_decap_8 FILLER_179_851 ();
 sg13g2_decap_8 FILLER_179_858 ();
 sg13g2_decap_4 FILLER_179_870 ();
 sg13g2_fill_2 FILLER_179_874 ();
 sg13g2_decap_8 FILLER_179_884 ();
 sg13g2_decap_8 FILLER_179_891 ();
 sg13g2_decap_8 FILLER_179_898 ();
 sg13g2_decap_8 FILLER_179_905 ();
 sg13g2_decap_8 FILLER_179_912 ();
 sg13g2_decap_8 FILLER_179_919 ();
 sg13g2_decap_8 FILLER_179_926 ();
 sg13g2_fill_2 FILLER_179_933 ();
 sg13g2_fill_1 FILLER_179_935 ();
 sg13g2_fill_2 FILLER_179_939 ();
 sg13g2_decap_8 FILLER_179_949 ();
 sg13g2_decap_8 FILLER_179_956 ();
 sg13g2_decap_8 FILLER_179_963 ();
 sg13g2_decap_8 FILLER_179_970 ();
 sg13g2_decap_8 FILLER_179_977 ();
 sg13g2_decap_8 FILLER_179_984 ();
 sg13g2_decap_8 FILLER_179_991 ();
 sg13g2_decap_8 FILLER_179_998 ();
 sg13g2_decap_8 FILLER_179_1005 ();
 sg13g2_decap_8 FILLER_179_1012 ();
 sg13g2_decap_8 FILLER_179_1019 ();
 sg13g2_decap_8 FILLER_179_1026 ();
 sg13g2_decap_8 FILLER_179_1033 ();
 sg13g2_decap_8 FILLER_179_1040 ();
 sg13g2_decap_8 FILLER_179_1047 ();
 sg13g2_decap_8 FILLER_179_1054 ();
 sg13g2_decap_8 FILLER_179_1061 ();
 sg13g2_decap_8 FILLER_179_1068 ();
 sg13g2_decap_8 FILLER_179_1075 ();
 sg13g2_decap_8 FILLER_179_1082 ();
 sg13g2_decap_8 FILLER_179_1089 ();
 sg13g2_decap_8 FILLER_179_1096 ();
 sg13g2_decap_8 FILLER_179_1103 ();
 sg13g2_decap_8 FILLER_179_1110 ();
 sg13g2_decap_8 FILLER_179_1117 ();
 sg13g2_decap_8 FILLER_179_1124 ();
 sg13g2_decap_8 FILLER_179_1131 ();
 sg13g2_decap_8 FILLER_179_1138 ();
 sg13g2_decap_8 FILLER_179_1145 ();
 sg13g2_decap_8 FILLER_179_1152 ();
 sg13g2_decap_8 FILLER_179_1159 ();
 sg13g2_decap_8 FILLER_179_1166 ();
 sg13g2_decap_8 FILLER_179_1173 ();
 sg13g2_decap_8 FILLER_179_1180 ();
 sg13g2_decap_8 FILLER_179_1187 ();
 sg13g2_decap_8 FILLER_179_1194 ();
 sg13g2_decap_8 FILLER_179_1201 ();
 sg13g2_decap_8 FILLER_179_1208 ();
 sg13g2_decap_8 FILLER_179_1215 ();
 sg13g2_decap_8 FILLER_179_1222 ();
 sg13g2_decap_8 FILLER_179_1229 ();
 sg13g2_decap_8 FILLER_179_1236 ();
 sg13g2_decap_8 FILLER_179_1243 ();
 sg13g2_decap_8 FILLER_179_1250 ();
 sg13g2_decap_8 FILLER_179_1257 ();
 sg13g2_decap_8 FILLER_179_1264 ();
 sg13g2_decap_8 FILLER_179_1271 ();
 sg13g2_decap_8 FILLER_179_1278 ();
 sg13g2_decap_8 FILLER_179_1285 ();
 sg13g2_decap_8 FILLER_179_1292 ();
 sg13g2_decap_8 FILLER_179_1299 ();
 sg13g2_decap_8 FILLER_179_1306 ();
 sg13g2_decap_8 FILLER_179_1313 ();
 sg13g2_decap_8 FILLER_179_1320 ();
 sg13g2_decap_8 FILLER_179_1327 ();
 sg13g2_decap_8 FILLER_179_1334 ();
 sg13g2_decap_8 FILLER_179_1341 ();
 sg13g2_decap_8 FILLER_179_1348 ();
 sg13g2_decap_8 FILLER_179_1355 ();
 sg13g2_decap_8 FILLER_179_1362 ();
 sg13g2_decap_8 FILLER_179_1369 ();
 sg13g2_decap_8 FILLER_179_1376 ();
 sg13g2_decap_8 FILLER_179_1383 ();
 sg13g2_decap_8 FILLER_179_1390 ();
 sg13g2_decap_8 FILLER_179_1397 ();
 sg13g2_decap_8 FILLER_179_1404 ();
 sg13g2_decap_8 FILLER_179_1411 ();
 sg13g2_decap_8 FILLER_179_1418 ();
 sg13g2_decap_8 FILLER_179_1425 ();
 sg13g2_decap_8 FILLER_179_1432 ();
 sg13g2_decap_8 FILLER_179_1439 ();
 sg13g2_decap_8 FILLER_179_1446 ();
 sg13g2_decap_8 FILLER_179_1453 ();
 sg13g2_decap_8 FILLER_179_1460 ();
 sg13g2_decap_8 FILLER_179_1467 ();
 sg13g2_decap_8 FILLER_179_1474 ();
 sg13g2_decap_8 FILLER_179_1481 ();
 sg13g2_decap_8 FILLER_179_1488 ();
 sg13g2_decap_8 FILLER_179_1495 ();
 sg13g2_decap_8 FILLER_179_1502 ();
 sg13g2_decap_8 FILLER_179_1509 ();
 sg13g2_decap_8 FILLER_179_1516 ();
 sg13g2_decap_8 FILLER_179_1523 ();
 sg13g2_decap_8 FILLER_179_1530 ();
 sg13g2_decap_8 FILLER_179_1537 ();
 sg13g2_decap_8 FILLER_179_1544 ();
 sg13g2_decap_8 FILLER_179_1551 ();
 sg13g2_decap_8 FILLER_179_1558 ();
 sg13g2_decap_8 FILLER_179_1565 ();
 sg13g2_decap_8 FILLER_179_1572 ();
 sg13g2_decap_8 FILLER_179_1579 ();
 sg13g2_decap_8 FILLER_179_1586 ();
 sg13g2_decap_8 FILLER_179_1593 ();
 sg13g2_decap_8 FILLER_179_1600 ();
 sg13g2_decap_8 FILLER_179_1607 ();
 sg13g2_decap_8 FILLER_179_1614 ();
 sg13g2_decap_8 FILLER_179_1621 ();
 sg13g2_decap_8 FILLER_179_1628 ();
 sg13g2_decap_8 FILLER_179_1635 ();
 sg13g2_decap_8 FILLER_179_1642 ();
 sg13g2_decap_8 FILLER_179_1649 ();
 sg13g2_decap_8 FILLER_179_1656 ();
 sg13g2_decap_8 FILLER_179_1663 ();
 sg13g2_decap_8 FILLER_179_1670 ();
 sg13g2_decap_8 FILLER_179_1677 ();
 sg13g2_decap_8 FILLER_179_1684 ();
 sg13g2_decap_8 FILLER_179_1691 ();
 sg13g2_decap_8 FILLER_179_1698 ();
 sg13g2_decap_8 FILLER_179_1705 ();
 sg13g2_decap_8 FILLER_179_1712 ();
 sg13g2_decap_8 FILLER_179_1719 ();
 sg13g2_decap_8 FILLER_179_1726 ();
 sg13g2_decap_8 FILLER_179_1733 ();
 sg13g2_decap_8 FILLER_179_1740 ();
 sg13g2_decap_8 FILLER_179_1747 ();
 sg13g2_decap_8 FILLER_179_1754 ();
 sg13g2_decap_8 FILLER_179_1761 ();
 sg13g2_decap_8 FILLER_180_0 ();
 sg13g2_decap_8 FILLER_180_7 ();
 sg13g2_decap_8 FILLER_180_14 ();
 sg13g2_decap_8 FILLER_180_21 ();
 sg13g2_decap_8 FILLER_180_28 ();
 sg13g2_decap_8 FILLER_180_35 ();
 sg13g2_decap_8 FILLER_180_42 ();
 sg13g2_decap_8 FILLER_180_49 ();
 sg13g2_decap_8 FILLER_180_56 ();
 sg13g2_decap_8 FILLER_180_63 ();
 sg13g2_decap_8 FILLER_180_70 ();
 sg13g2_decap_8 FILLER_180_77 ();
 sg13g2_decap_8 FILLER_180_84 ();
 sg13g2_decap_8 FILLER_180_91 ();
 sg13g2_decap_8 FILLER_180_98 ();
 sg13g2_decap_8 FILLER_180_105 ();
 sg13g2_decap_8 FILLER_180_112 ();
 sg13g2_decap_8 FILLER_180_119 ();
 sg13g2_decap_8 FILLER_180_126 ();
 sg13g2_decap_8 FILLER_180_133 ();
 sg13g2_decap_8 FILLER_180_140 ();
 sg13g2_decap_8 FILLER_180_147 ();
 sg13g2_decap_8 FILLER_180_154 ();
 sg13g2_decap_8 FILLER_180_161 ();
 sg13g2_decap_8 FILLER_180_168 ();
 sg13g2_decap_8 FILLER_180_175 ();
 sg13g2_decap_8 FILLER_180_182 ();
 sg13g2_decap_8 FILLER_180_189 ();
 sg13g2_fill_1 FILLER_180_196 ();
 sg13g2_decap_8 FILLER_180_232 ();
 sg13g2_decap_8 FILLER_180_239 ();
 sg13g2_decap_8 FILLER_180_246 ();
 sg13g2_decap_8 FILLER_180_253 ();
 sg13g2_decap_8 FILLER_180_260 ();
 sg13g2_decap_8 FILLER_180_267 ();
 sg13g2_decap_8 FILLER_180_274 ();
 sg13g2_decap_8 FILLER_180_281 ();
 sg13g2_decap_8 FILLER_180_288 ();
 sg13g2_decap_8 FILLER_180_295 ();
 sg13g2_decap_8 FILLER_180_302 ();
 sg13g2_decap_8 FILLER_180_309 ();
 sg13g2_decap_8 FILLER_180_316 ();
 sg13g2_decap_8 FILLER_180_323 ();
 sg13g2_decap_8 FILLER_180_330 ();
 sg13g2_decap_8 FILLER_180_337 ();
 sg13g2_decap_8 FILLER_180_349 ();
 sg13g2_decap_8 FILLER_180_356 ();
 sg13g2_decap_8 FILLER_180_363 ();
 sg13g2_decap_8 FILLER_180_370 ();
 sg13g2_decap_8 FILLER_180_377 ();
 sg13g2_decap_8 FILLER_180_384 ();
 sg13g2_decap_8 FILLER_180_391 ();
 sg13g2_decap_8 FILLER_180_398 ();
 sg13g2_decap_4 FILLER_180_430 ();
 sg13g2_decap_8 FILLER_180_440 ();
 sg13g2_decap_8 FILLER_180_447 ();
 sg13g2_decap_8 FILLER_180_454 ();
 sg13g2_decap_8 FILLER_180_461 ();
 sg13g2_decap_8 FILLER_180_468 ();
 sg13g2_decap_8 FILLER_180_475 ();
 sg13g2_decap_8 FILLER_180_482 ();
 sg13g2_decap_8 FILLER_180_489 ();
 sg13g2_decap_8 FILLER_180_496 ();
 sg13g2_fill_2 FILLER_180_503 ();
 sg13g2_fill_2 FILLER_180_520 ();
 sg13g2_fill_1 FILLER_180_522 ();
 sg13g2_decap_4 FILLER_180_528 ();
 sg13g2_fill_2 FILLER_180_537 ();
 sg13g2_fill_1 FILLER_180_552 ();
 sg13g2_decap_8 FILLER_180_558 ();
 sg13g2_decap_8 FILLER_180_565 ();
 sg13g2_decap_8 FILLER_180_572 ();
 sg13g2_decap_8 FILLER_180_579 ();
 sg13g2_decap_8 FILLER_180_586 ();
 sg13g2_decap_8 FILLER_180_593 ();
 sg13g2_decap_8 FILLER_180_600 ();
 sg13g2_decap_8 FILLER_180_607 ();
 sg13g2_decap_8 FILLER_180_614 ();
 sg13g2_decap_8 FILLER_180_621 ();
 sg13g2_decap_8 FILLER_180_628 ();
 sg13g2_decap_8 FILLER_180_635 ();
 sg13g2_decap_8 FILLER_180_642 ();
 sg13g2_decap_8 FILLER_180_649 ();
 sg13g2_decap_8 FILLER_180_656 ();
 sg13g2_decap_8 FILLER_180_663 ();
 sg13g2_decap_8 FILLER_180_670 ();
 sg13g2_decap_8 FILLER_180_677 ();
 sg13g2_decap_8 FILLER_180_684 ();
 sg13g2_decap_8 FILLER_180_691 ();
 sg13g2_fill_2 FILLER_180_698 ();
 sg13g2_fill_1 FILLER_180_707 ();
 sg13g2_decap_8 FILLER_180_718 ();
 sg13g2_decap_8 FILLER_180_725 ();
 sg13g2_decap_8 FILLER_180_732 ();
 sg13g2_decap_8 FILLER_180_739 ();
 sg13g2_decap_8 FILLER_180_746 ();
 sg13g2_decap_8 FILLER_180_753 ();
 sg13g2_decap_8 FILLER_180_760 ();
 sg13g2_decap_8 FILLER_180_767 ();
 sg13g2_decap_8 FILLER_180_774 ();
 sg13g2_decap_8 FILLER_180_781 ();
 sg13g2_decap_8 FILLER_180_788 ();
 sg13g2_decap_8 FILLER_180_795 ();
 sg13g2_decap_8 FILLER_180_802 ();
 sg13g2_decap_8 FILLER_180_809 ();
 sg13g2_fill_2 FILLER_180_816 ();
 sg13g2_fill_1 FILLER_180_818 ();
 sg13g2_decap_8 FILLER_180_824 ();
 sg13g2_decap_8 FILLER_180_831 ();
 sg13g2_decap_8 FILLER_180_838 ();
 sg13g2_decap_8 FILLER_180_845 ();
 sg13g2_decap_8 FILLER_180_852 ();
 sg13g2_decap_8 FILLER_180_859 ();
 sg13g2_decap_8 FILLER_180_866 ();
 sg13g2_decap_8 FILLER_180_873 ();
 sg13g2_decap_8 FILLER_180_880 ();
 sg13g2_decap_8 FILLER_180_887 ();
 sg13g2_decap_8 FILLER_180_894 ();
 sg13g2_decap_8 FILLER_180_901 ();
 sg13g2_decap_8 FILLER_180_908 ();
 sg13g2_decap_8 FILLER_180_915 ();
 sg13g2_decap_8 FILLER_180_922 ();
 sg13g2_decap_8 FILLER_180_929 ();
 sg13g2_decap_8 FILLER_180_936 ();
 sg13g2_decap_8 FILLER_180_943 ();
 sg13g2_decap_8 FILLER_180_950 ();
 sg13g2_decap_8 FILLER_180_957 ();
 sg13g2_decap_8 FILLER_180_964 ();
 sg13g2_decap_8 FILLER_180_971 ();
 sg13g2_decap_8 FILLER_180_978 ();
 sg13g2_decap_8 FILLER_180_985 ();
 sg13g2_decap_8 FILLER_180_992 ();
 sg13g2_decap_8 FILLER_180_999 ();
 sg13g2_decap_8 FILLER_180_1006 ();
 sg13g2_decap_8 FILLER_180_1013 ();
 sg13g2_decap_8 FILLER_180_1020 ();
 sg13g2_decap_8 FILLER_180_1027 ();
 sg13g2_decap_8 FILLER_180_1034 ();
 sg13g2_decap_8 FILLER_180_1041 ();
 sg13g2_decap_8 FILLER_180_1048 ();
 sg13g2_decap_8 FILLER_180_1055 ();
 sg13g2_decap_8 FILLER_180_1062 ();
 sg13g2_decap_8 FILLER_180_1069 ();
 sg13g2_decap_8 FILLER_180_1076 ();
 sg13g2_decap_8 FILLER_180_1083 ();
 sg13g2_decap_8 FILLER_180_1090 ();
 sg13g2_decap_8 FILLER_180_1097 ();
 sg13g2_decap_8 FILLER_180_1104 ();
 sg13g2_decap_8 FILLER_180_1111 ();
 sg13g2_decap_8 FILLER_180_1118 ();
 sg13g2_decap_8 FILLER_180_1125 ();
 sg13g2_decap_8 FILLER_180_1132 ();
 sg13g2_decap_8 FILLER_180_1139 ();
 sg13g2_decap_8 FILLER_180_1146 ();
 sg13g2_decap_8 FILLER_180_1153 ();
 sg13g2_decap_8 FILLER_180_1160 ();
 sg13g2_decap_8 FILLER_180_1167 ();
 sg13g2_decap_8 FILLER_180_1174 ();
 sg13g2_decap_8 FILLER_180_1181 ();
 sg13g2_decap_8 FILLER_180_1188 ();
 sg13g2_decap_8 FILLER_180_1195 ();
 sg13g2_decap_8 FILLER_180_1202 ();
 sg13g2_decap_8 FILLER_180_1209 ();
 sg13g2_decap_8 FILLER_180_1216 ();
 sg13g2_decap_8 FILLER_180_1223 ();
 sg13g2_decap_8 FILLER_180_1230 ();
 sg13g2_decap_8 FILLER_180_1237 ();
 sg13g2_decap_8 FILLER_180_1244 ();
 sg13g2_decap_8 FILLER_180_1251 ();
 sg13g2_decap_8 FILLER_180_1258 ();
 sg13g2_decap_8 FILLER_180_1265 ();
 sg13g2_decap_8 FILLER_180_1272 ();
 sg13g2_decap_8 FILLER_180_1279 ();
 sg13g2_decap_8 FILLER_180_1286 ();
 sg13g2_decap_8 FILLER_180_1293 ();
 sg13g2_decap_8 FILLER_180_1300 ();
 sg13g2_decap_8 FILLER_180_1307 ();
 sg13g2_decap_8 FILLER_180_1314 ();
 sg13g2_decap_8 FILLER_180_1321 ();
 sg13g2_decap_8 FILLER_180_1328 ();
 sg13g2_decap_8 FILLER_180_1335 ();
 sg13g2_decap_8 FILLER_180_1342 ();
 sg13g2_decap_8 FILLER_180_1349 ();
 sg13g2_decap_8 FILLER_180_1356 ();
 sg13g2_decap_8 FILLER_180_1363 ();
 sg13g2_decap_8 FILLER_180_1370 ();
 sg13g2_decap_8 FILLER_180_1377 ();
 sg13g2_decap_8 FILLER_180_1384 ();
 sg13g2_decap_8 FILLER_180_1391 ();
 sg13g2_decap_8 FILLER_180_1398 ();
 sg13g2_decap_8 FILLER_180_1405 ();
 sg13g2_decap_8 FILLER_180_1412 ();
 sg13g2_decap_8 FILLER_180_1419 ();
 sg13g2_decap_8 FILLER_180_1426 ();
 sg13g2_decap_8 FILLER_180_1433 ();
 sg13g2_decap_8 FILLER_180_1440 ();
 sg13g2_decap_8 FILLER_180_1447 ();
 sg13g2_decap_8 FILLER_180_1454 ();
 sg13g2_decap_8 FILLER_180_1461 ();
 sg13g2_decap_8 FILLER_180_1468 ();
 sg13g2_decap_8 FILLER_180_1475 ();
 sg13g2_decap_8 FILLER_180_1482 ();
 sg13g2_decap_8 FILLER_180_1489 ();
 sg13g2_decap_8 FILLER_180_1496 ();
 sg13g2_decap_8 FILLER_180_1503 ();
 sg13g2_decap_8 FILLER_180_1510 ();
 sg13g2_decap_8 FILLER_180_1517 ();
 sg13g2_decap_8 FILLER_180_1524 ();
 sg13g2_decap_8 FILLER_180_1531 ();
 sg13g2_decap_8 FILLER_180_1538 ();
 sg13g2_decap_8 FILLER_180_1545 ();
 sg13g2_decap_8 FILLER_180_1552 ();
 sg13g2_decap_8 FILLER_180_1559 ();
 sg13g2_decap_8 FILLER_180_1566 ();
 sg13g2_decap_8 FILLER_180_1573 ();
 sg13g2_decap_8 FILLER_180_1580 ();
 sg13g2_decap_8 FILLER_180_1587 ();
 sg13g2_decap_8 FILLER_180_1594 ();
 sg13g2_decap_8 FILLER_180_1601 ();
 sg13g2_decap_8 FILLER_180_1608 ();
 sg13g2_decap_8 FILLER_180_1615 ();
 sg13g2_decap_8 FILLER_180_1622 ();
 sg13g2_decap_8 FILLER_180_1629 ();
 sg13g2_decap_8 FILLER_180_1636 ();
 sg13g2_decap_8 FILLER_180_1643 ();
 sg13g2_decap_8 FILLER_180_1650 ();
 sg13g2_decap_8 FILLER_180_1657 ();
 sg13g2_decap_8 FILLER_180_1664 ();
 sg13g2_decap_8 FILLER_180_1671 ();
 sg13g2_decap_8 FILLER_180_1678 ();
 sg13g2_decap_8 FILLER_180_1685 ();
 sg13g2_decap_8 FILLER_180_1692 ();
 sg13g2_decap_8 FILLER_180_1699 ();
 sg13g2_decap_8 FILLER_180_1706 ();
 sg13g2_decap_8 FILLER_180_1713 ();
 sg13g2_decap_8 FILLER_180_1720 ();
 sg13g2_decap_8 FILLER_180_1727 ();
 sg13g2_decap_8 FILLER_180_1734 ();
 sg13g2_decap_8 FILLER_180_1741 ();
 sg13g2_decap_8 FILLER_180_1748 ();
 sg13g2_decap_8 FILLER_180_1755 ();
 sg13g2_decap_4 FILLER_180_1762 ();
 sg13g2_fill_2 FILLER_180_1766 ();
 sg13g2_decap_8 FILLER_181_0 ();
 sg13g2_decap_8 FILLER_181_7 ();
 sg13g2_decap_8 FILLER_181_14 ();
 sg13g2_decap_8 FILLER_181_21 ();
 sg13g2_decap_8 FILLER_181_28 ();
 sg13g2_decap_8 FILLER_181_35 ();
 sg13g2_decap_8 FILLER_181_42 ();
 sg13g2_decap_8 FILLER_181_49 ();
 sg13g2_decap_8 FILLER_181_56 ();
 sg13g2_decap_8 FILLER_181_63 ();
 sg13g2_decap_8 FILLER_181_70 ();
 sg13g2_decap_8 FILLER_181_77 ();
 sg13g2_decap_8 FILLER_181_84 ();
 sg13g2_decap_8 FILLER_181_91 ();
 sg13g2_decap_8 FILLER_181_98 ();
 sg13g2_decap_8 FILLER_181_105 ();
 sg13g2_decap_8 FILLER_181_112 ();
 sg13g2_decap_8 FILLER_181_119 ();
 sg13g2_decap_8 FILLER_181_126 ();
 sg13g2_decap_8 FILLER_181_133 ();
 sg13g2_decap_8 FILLER_181_140 ();
 sg13g2_decap_8 FILLER_181_147 ();
 sg13g2_decap_8 FILLER_181_154 ();
 sg13g2_decap_8 FILLER_181_161 ();
 sg13g2_decap_8 FILLER_181_168 ();
 sg13g2_decap_8 FILLER_181_175 ();
 sg13g2_decap_8 FILLER_181_182 ();
 sg13g2_decap_8 FILLER_181_189 ();
 sg13g2_decap_8 FILLER_181_196 ();
 sg13g2_decap_8 FILLER_181_227 ();
 sg13g2_decap_8 FILLER_181_234 ();
 sg13g2_decap_8 FILLER_181_241 ();
 sg13g2_decap_8 FILLER_181_248 ();
 sg13g2_decap_8 FILLER_181_255 ();
 sg13g2_decap_8 FILLER_181_262 ();
 sg13g2_decap_8 FILLER_181_269 ();
 sg13g2_decap_8 FILLER_181_276 ();
 sg13g2_decap_8 FILLER_181_283 ();
 sg13g2_decap_8 FILLER_181_290 ();
 sg13g2_decap_8 FILLER_181_297 ();
 sg13g2_decap_8 FILLER_181_304 ();
 sg13g2_decap_8 FILLER_181_311 ();
 sg13g2_decap_8 FILLER_181_318 ();
 sg13g2_decap_8 FILLER_181_325 ();
 sg13g2_decap_8 FILLER_181_332 ();
 sg13g2_fill_1 FILLER_181_339 ();
 sg13g2_decap_4 FILLER_181_350 ();
 sg13g2_decap_8 FILLER_181_364 ();
 sg13g2_fill_2 FILLER_181_371 ();
 sg13g2_decap_8 FILLER_181_399 ();
 sg13g2_decap_8 FILLER_181_406 ();
 sg13g2_decap_8 FILLER_181_413 ();
 sg13g2_decap_8 FILLER_181_420 ();
 sg13g2_decap_8 FILLER_181_427 ();
 sg13g2_decap_8 FILLER_181_469 ();
 sg13g2_decap_8 FILLER_181_476 ();
 sg13g2_decap_8 FILLER_181_483 ();
 sg13g2_decap_8 FILLER_181_490 ();
 sg13g2_decap_8 FILLER_181_497 ();
 sg13g2_decap_8 FILLER_181_504 ();
 sg13g2_fill_2 FILLER_181_511 ();
 sg13g2_fill_1 FILLER_181_513 ();
 sg13g2_fill_2 FILLER_181_540 ();
 sg13g2_decap_8 FILLER_181_555 ();
 sg13g2_decap_8 FILLER_181_562 ();
 sg13g2_decap_8 FILLER_181_569 ();
 sg13g2_decap_8 FILLER_181_576 ();
 sg13g2_decap_8 FILLER_181_583 ();
 sg13g2_decap_8 FILLER_181_590 ();
 sg13g2_decap_8 FILLER_181_597 ();
 sg13g2_decap_8 FILLER_181_604 ();
 sg13g2_decap_8 FILLER_181_611 ();
 sg13g2_decap_8 FILLER_181_618 ();
 sg13g2_decap_8 FILLER_181_625 ();
 sg13g2_decap_8 FILLER_181_632 ();
 sg13g2_decap_8 FILLER_181_639 ();
 sg13g2_decap_8 FILLER_181_646 ();
 sg13g2_decap_8 FILLER_181_653 ();
 sg13g2_decap_8 FILLER_181_660 ();
 sg13g2_decap_8 FILLER_181_667 ();
 sg13g2_decap_8 FILLER_181_674 ();
 sg13g2_decap_8 FILLER_181_681 ();
 sg13g2_decap_8 FILLER_181_688 ();
 sg13g2_decap_8 FILLER_181_695 ();
 sg13g2_fill_2 FILLER_181_702 ();
 sg13g2_decap_8 FILLER_181_716 ();
 sg13g2_decap_8 FILLER_181_723 ();
 sg13g2_decap_8 FILLER_181_730 ();
 sg13g2_decap_8 FILLER_181_737 ();
 sg13g2_decap_8 FILLER_181_744 ();
 sg13g2_decap_8 FILLER_181_751 ();
 sg13g2_decap_8 FILLER_181_758 ();
 sg13g2_decap_8 FILLER_181_765 ();
 sg13g2_decap_8 FILLER_181_772 ();
 sg13g2_decap_8 FILLER_181_779 ();
 sg13g2_decap_8 FILLER_181_786 ();
 sg13g2_decap_8 FILLER_181_793 ();
 sg13g2_decap_8 FILLER_181_800 ();
 sg13g2_decap_8 FILLER_181_807 ();
 sg13g2_decap_8 FILLER_181_814 ();
 sg13g2_decap_8 FILLER_181_821 ();
 sg13g2_decap_8 FILLER_181_828 ();
 sg13g2_decap_8 FILLER_181_835 ();
 sg13g2_decap_8 FILLER_181_842 ();
 sg13g2_decap_8 FILLER_181_849 ();
 sg13g2_decap_8 FILLER_181_856 ();
 sg13g2_decap_8 FILLER_181_863 ();
 sg13g2_decap_8 FILLER_181_870 ();
 sg13g2_decap_8 FILLER_181_877 ();
 sg13g2_decap_8 FILLER_181_884 ();
 sg13g2_decap_8 FILLER_181_891 ();
 sg13g2_decap_8 FILLER_181_898 ();
 sg13g2_decap_8 FILLER_181_905 ();
 sg13g2_decap_8 FILLER_181_912 ();
 sg13g2_decap_8 FILLER_181_919 ();
 sg13g2_decap_8 FILLER_181_926 ();
 sg13g2_decap_8 FILLER_181_933 ();
 sg13g2_decap_8 FILLER_181_940 ();
 sg13g2_decap_8 FILLER_181_947 ();
 sg13g2_decap_8 FILLER_181_954 ();
 sg13g2_decap_8 FILLER_181_961 ();
 sg13g2_decap_8 FILLER_181_968 ();
 sg13g2_decap_8 FILLER_181_975 ();
 sg13g2_decap_8 FILLER_181_982 ();
 sg13g2_decap_8 FILLER_181_989 ();
 sg13g2_decap_8 FILLER_181_996 ();
 sg13g2_decap_8 FILLER_181_1003 ();
 sg13g2_decap_8 FILLER_181_1010 ();
 sg13g2_decap_8 FILLER_181_1017 ();
 sg13g2_decap_8 FILLER_181_1024 ();
 sg13g2_decap_8 FILLER_181_1031 ();
 sg13g2_decap_8 FILLER_181_1038 ();
 sg13g2_decap_8 FILLER_181_1045 ();
 sg13g2_decap_8 FILLER_181_1052 ();
 sg13g2_decap_8 FILLER_181_1059 ();
 sg13g2_decap_8 FILLER_181_1066 ();
 sg13g2_decap_8 FILLER_181_1073 ();
 sg13g2_decap_8 FILLER_181_1080 ();
 sg13g2_decap_8 FILLER_181_1087 ();
 sg13g2_decap_8 FILLER_181_1094 ();
 sg13g2_decap_8 FILLER_181_1101 ();
 sg13g2_decap_8 FILLER_181_1108 ();
 sg13g2_decap_8 FILLER_181_1115 ();
 sg13g2_decap_8 FILLER_181_1122 ();
 sg13g2_decap_8 FILLER_181_1129 ();
 sg13g2_decap_8 FILLER_181_1136 ();
 sg13g2_decap_8 FILLER_181_1143 ();
 sg13g2_decap_8 FILLER_181_1150 ();
 sg13g2_decap_8 FILLER_181_1157 ();
 sg13g2_decap_8 FILLER_181_1164 ();
 sg13g2_decap_8 FILLER_181_1171 ();
 sg13g2_decap_8 FILLER_181_1178 ();
 sg13g2_decap_8 FILLER_181_1185 ();
 sg13g2_decap_8 FILLER_181_1192 ();
 sg13g2_decap_8 FILLER_181_1199 ();
 sg13g2_decap_8 FILLER_181_1206 ();
 sg13g2_decap_8 FILLER_181_1213 ();
 sg13g2_decap_8 FILLER_181_1220 ();
 sg13g2_decap_8 FILLER_181_1227 ();
 sg13g2_decap_8 FILLER_181_1234 ();
 sg13g2_decap_8 FILLER_181_1241 ();
 sg13g2_decap_8 FILLER_181_1248 ();
 sg13g2_decap_8 FILLER_181_1255 ();
 sg13g2_decap_8 FILLER_181_1262 ();
 sg13g2_decap_8 FILLER_181_1269 ();
 sg13g2_decap_8 FILLER_181_1276 ();
 sg13g2_decap_8 FILLER_181_1283 ();
 sg13g2_decap_8 FILLER_181_1290 ();
 sg13g2_decap_8 FILLER_181_1297 ();
 sg13g2_decap_8 FILLER_181_1304 ();
 sg13g2_decap_8 FILLER_181_1311 ();
 sg13g2_decap_8 FILLER_181_1318 ();
 sg13g2_decap_8 FILLER_181_1325 ();
 sg13g2_decap_8 FILLER_181_1332 ();
 sg13g2_decap_8 FILLER_181_1339 ();
 sg13g2_decap_8 FILLER_181_1346 ();
 sg13g2_decap_8 FILLER_181_1353 ();
 sg13g2_decap_8 FILLER_181_1360 ();
 sg13g2_decap_8 FILLER_181_1367 ();
 sg13g2_decap_8 FILLER_181_1374 ();
 sg13g2_decap_8 FILLER_181_1381 ();
 sg13g2_decap_8 FILLER_181_1388 ();
 sg13g2_decap_8 FILLER_181_1395 ();
 sg13g2_decap_8 FILLER_181_1402 ();
 sg13g2_decap_8 FILLER_181_1409 ();
 sg13g2_decap_8 FILLER_181_1416 ();
 sg13g2_decap_8 FILLER_181_1423 ();
 sg13g2_decap_8 FILLER_181_1430 ();
 sg13g2_decap_8 FILLER_181_1437 ();
 sg13g2_decap_8 FILLER_181_1444 ();
 sg13g2_decap_8 FILLER_181_1451 ();
 sg13g2_decap_8 FILLER_181_1458 ();
 sg13g2_decap_8 FILLER_181_1465 ();
 sg13g2_decap_8 FILLER_181_1472 ();
 sg13g2_decap_8 FILLER_181_1479 ();
 sg13g2_decap_8 FILLER_181_1486 ();
 sg13g2_decap_8 FILLER_181_1493 ();
 sg13g2_decap_8 FILLER_181_1500 ();
 sg13g2_decap_8 FILLER_181_1507 ();
 sg13g2_decap_8 FILLER_181_1514 ();
 sg13g2_decap_8 FILLER_181_1521 ();
 sg13g2_decap_8 FILLER_181_1528 ();
 sg13g2_decap_8 FILLER_181_1535 ();
 sg13g2_decap_8 FILLER_181_1542 ();
 sg13g2_decap_8 FILLER_181_1549 ();
 sg13g2_decap_8 FILLER_181_1556 ();
 sg13g2_decap_8 FILLER_181_1563 ();
 sg13g2_decap_8 FILLER_181_1570 ();
 sg13g2_decap_8 FILLER_181_1577 ();
 sg13g2_decap_8 FILLER_181_1584 ();
 sg13g2_decap_8 FILLER_181_1591 ();
 sg13g2_decap_8 FILLER_181_1598 ();
 sg13g2_decap_8 FILLER_181_1605 ();
 sg13g2_decap_8 FILLER_181_1612 ();
 sg13g2_decap_8 FILLER_181_1619 ();
 sg13g2_decap_8 FILLER_181_1626 ();
 sg13g2_decap_8 FILLER_181_1633 ();
 sg13g2_decap_8 FILLER_181_1640 ();
 sg13g2_decap_8 FILLER_181_1647 ();
 sg13g2_decap_8 FILLER_181_1654 ();
 sg13g2_decap_8 FILLER_181_1661 ();
 sg13g2_decap_8 FILLER_181_1668 ();
 sg13g2_decap_8 FILLER_181_1675 ();
 sg13g2_decap_8 FILLER_181_1682 ();
 sg13g2_decap_8 FILLER_181_1689 ();
 sg13g2_decap_8 FILLER_181_1696 ();
 sg13g2_decap_8 FILLER_181_1703 ();
 sg13g2_decap_8 FILLER_181_1710 ();
 sg13g2_decap_8 FILLER_181_1717 ();
 sg13g2_decap_8 FILLER_181_1724 ();
 sg13g2_decap_8 FILLER_181_1731 ();
 sg13g2_decap_8 FILLER_181_1738 ();
 sg13g2_decap_8 FILLER_181_1745 ();
 sg13g2_decap_8 FILLER_181_1752 ();
 sg13g2_decap_8 FILLER_181_1759 ();
 sg13g2_fill_2 FILLER_181_1766 ();
 sg13g2_decap_8 FILLER_182_0 ();
 sg13g2_decap_8 FILLER_182_7 ();
 sg13g2_decap_8 FILLER_182_14 ();
 sg13g2_decap_8 FILLER_182_21 ();
 sg13g2_decap_8 FILLER_182_28 ();
 sg13g2_decap_8 FILLER_182_35 ();
 sg13g2_decap_8 FILLER_182_42 ();
 sg13g2_decap_8 FILLER_182_49 ();
 sg13g2_decap_8 FILLER_182_56 ();
 sg13g2_decap_8 FILLER_182_63 ();
 sg13g2_decap_8 FILLER_182_70 ();
 sg13g2_decap_8 FILLER_182_77 ();
 sg13g2_decap_8 FILLER_182_84 ();
 sg13g2_decap_8 FILLER_182_91 ();
 sg13g2_decap_8 FILLER_182_98 ();
 sg13g2_decap_8 FILLER_182_105 ();
 sg13g2_decap_8 FILLER_182_112 ();
 sg13g2_decap_8 FILLER_182_119 ();
 sg13g2_decap_8 FILLER_182_126 ();
 sg13g2_decap_8 FILLER_182_133 ();
 sg13g2_decap_8 FILLER_182_140 ();
 sg13g2_decap_8 FILLER_182_147 ();
 sg13g2_decap_8 FILLER_182_154 ();
 sg13g2_decap_8 FILLER_182_161 ();
 sg13g2_decap_8 FILLER_182_168 ();
 sg13g2_decap_8 FILLER_182_175 ();
 sg13g2_decap_8 FILLER_182_182 ();
 sg13g2_decap_8 FILLER_182_189 ();
 sg13g2_decap_8 FILLER_182_196 ();
 sg13g2_decap_8 FILLER_182_203 ();
 sg13g2_decap_4 FILLER_182_210 ();
 sg13g2_decap_8 FILLER_182_219 ();
 sg13g2_decap_8 FILLER_182_226 ();
 sg13g2_decap_8 FILLER_182_233 ();
 sg13g2_decap_8 FILLER_182_240 ();
 sg13g2_decap_8 FILLER_182_247 ();
 sg13g2_decap_8 FILLER_182_254 ();
 sg13g2_decap_8 FILLER_182_261 ();
 sg13g2_decap_8 FILLER_182_268 ();
 sg13g2_decap_8 FILLER_182_275 ();
 sg13g2_decap_8 FILLER_182_282 ();
 sg13g2_decap_8 FILLER_182_289 ();
 sg13g2_decap_8 FILLER_182_296 ();
 sg13g2_decap_8 FILLER_182_303 ();
 sg13g2_decap_8 FILLER_182_310 ();
 sg13g2_decap_8 FILLER_182_317 ();
 sg13g2_decap_4 FILLER_182_324 ();
 sg13g2_fill_2 FILLER_182_328 ();
 sg13g2_fill_1 FILLER_182_356 ();
 sg13g2_decap_8 FILLER_182_366 ();
 sg13g2_decap_4 FILLER_182_373 ();
 sg13g2_fill_1 FILLER_182_377 ();
 sg13g2_decap_8 FILLER_182_392 ();
 sg13g2_fill_2 FILLER_182_399 ();
 sg13g2_fill_1 FILLER_182_401 ();
 sg13g2_decap_8 FILLER_182_406 ();
 sg13g2_decap_8 FILLER_182_413 ();
 sg13g2_decap_8 FILLER_182_420 ();
 sg13g2_decap_8 FILLER_182_427 ();
 sg13g2_decap_8 FILLER_182_437 ();
 sg13g2_decap_8 FILLER_182_444 ();
 sg13g2_decap_4 FILLER_182_451 ();
 sg13g2_decap_8 FILLER_182_481 ();
 sg13g2_decap_8 FILLER_182_488 ();
 sg13g2_decap_8 FILLER_182_495 ();
 sg13g2_decap_8 FILLER_182_502 ();
 sg13g2_decap_8 FILLER_182_509 ();
 sg13g2_decap_8 FILLER_182_516 ();
 sg13g2_decap_8 FILLER_182_523 ();
 sg13g2_decap_8 FILLER_182_530 ();
 sg13g2_decap_4 FILLER_182_537 ();
 sg13g2_fill_2 FILLER_182_541 ();
 sg13g2_decap_8 FILLER_182_548 ();
 sg13g2_decap_8 FILLER_182_555 ();
 sg13g2_decap_8 FILLER_182_562 ();
 sg13g2_decap_8 FILLER_182_569 ();
 sg13g2_decap_8 FILLER_182_576 ();
 sg13g2_fill_2 FILLER_182_583 ();
 sg13g2_fill_1 FILLER_182_585 ();
 sg13g2_decap_8 FILLER_182_611 ();
 sg13g2_decap_8 FILLER_182_618 ();
 sg13g2_decap_8 FILLER_182_625 ();
 sg13g2_decap_8 FILLER_182_632 ();
 sg13g2_decap_8 FILLER_182_639 ();
 sg13g2_decap_8 FILLER_182_646 ();
 sg13g2_decap_8 FILLER_182_653 ();
 sg13g2_decap_8 FILLER_182_660 ();
 sg13g2_decap_8 FILLER_182_667 ();
 sg13g2_decap_8 FILLER_182_674 ();
 sg13g2_decap_8 FILLER_182_681 ();
 sg13g2_decap_8 FILLER_182_688 ();
 sg13g2_decap_8 FILLER_182_695 ();
 sg13g2_decap_8 FILLER_182_702 ();
 sg13g2_decap_8 FILLER_182_709 ();
 sg13g2_decap_8 FILLER_182_716 ();
 sg13g2_decap_8 FILLER_182_723 ();
 sg13g2_decap_8 FILLER_182_730 ();
 sg13g2_decap_8 FILLER_182_737 ();
 sg13g2_decap_8 FILLER_182_744 ();
 sg13g2_decap_8 FILLER_182_751 ();
 sg13g2_decap_8 FILLER_182_758 ();
 sg13g2_decap_8 FILLER_182_765 ();
 sg13g2_decap_8 FILLER_182_772 ();
 sg13g2_decap_8 FILLER_182_779 ();
 sg13g2_decap_8 FILLER_182_786 ();
 sg13g2_decap_8 FILLER_182_793 ();
 sg13g2_decap_8 FILLER_182_800 ();
 sg13g2_decap_8 FILLER_182_807 ();
 sg13g2_decap_8 FILLER_182_814 ();
 sg13g2_decap_8 FILLER_182_821 ();
 sg13g2_decap_8 FILLER_182_828 ();
 sg13g2_decap_8 FILLER_182_835 ();
 sg13g2_decap_8 FILLER_182_842 ();
 sg13g2_decap_8 FILLER_182_849 ();
 sg13g2_decap_8 FILLER_182_856 ();
 sg13g2_decap_8 FILLER_182_863 ();
 sg13g2_decap_8 FILLER_182_870 ();
 sg13g2_decap_8 FILLER_182_877 ();
 sg13g2_decap_8 FILLER_182_884 ();
 sg13g2_decap_8 FILLER_182_891 ();
 sg13g2_decap_8 FILLER_182_898 ();
 sg13g2_decap_8 FILLER_182_905 ();
 sg13g2_decap_8 FILLER_182_912 ();
 sg13g2_decap_8 FILLER_182_919 ();
 sg13g2_decap_8 FILLER_182_926 ();
 sg13g2_decap_8 FILLER_182_933 ();
 sg13g2_decap_8 FILLER_182_940 ();
 sg13g2_decap_8 FILLER_182_947 ();
 sg13g2_decap_8 FILLER_182_954 ();
 sg13g2_decap_8 FILLER_182_961 ();
 sg13g2_decap_8 FILLER_182_968 ();
 sg13g2_decap_8 FILLER_182_975 ();
 sg13g2_decap_8 FILLER_182_982 ();
 sg13g2_decap_8 FILLER_182_989 ();
 sg13g2_decap_8 FILLER_182_996 ();
 sg13g2_decap_8 FILLER_182_1003 ();
 sg13g2_decap_8 FILLER_182_1010 ();
 sg13g2_decap_8 FILLER_182_1017 ();
 sg13g2_decap_8 FILLER_182_1024 ();
 sg13g2_decap_8 FILLER_182_1031 ();
 sg13g2_decap_8 FILLER_182_1038 ();
 sg13g2_decap_8 FILLER_182_1045 ();
 sg13g2_decap_8 FILLER_182_1052 ();
 sg13g2_decap_8 FILLER_182_1059 ();
 sg13g2_decap_8 FILLER_182_1066 ();
 sg13g2_decap_8 FILLER_182_1073 ();
 sg13g2_decap_8 FILLER_182_1080 ();
 sg13g2_decap_8 FILLER_182_1087 ();
 sg13g2_decap_8 FILLER_182_1094 ();
 sg13g2_decap_8 FILLER_182_1101 ();
 sg13g2_decap_8 FILLER_182_1108 ();
 sg13g2_decap_8 FILLER_182_1115 ();
 sg13g2_decap_8 FILLER_182_1122 ();
 sg13g2_decap_8 FILLER_182_1129 ();
 sg13g2_decap_8 FILLER_182_1136 ();
 sg13g2_decap_8 FILLER_182_1143 ();
 sg13g2_decap_8 FILLER_182_1150 ();
 sg13g2_decap_8 FILLER_182_1157 ();
 sg13g2_decap_8 FILLER_182_1164 ();
 sg13g2_decap_8 FILLER_182_1171 ();
 sg13g2_decap_8 FILLER_182_1178 ();
 sg13g2_decap_8 FILLER_182_1185 ();
 sg13g2_decap_8 FILLER_182_1192 ();
 sg13g2_decap_8 FILLER_182_1199 ();
 sg13g2_decap_8 FILLER_182_1206 ();
 sg13g2_decap_8 FILLER_182_1213 ();
 sg13g2_decap_8 FILLER_182_1220 ();
 sg13g2_decap_8 FILLER_182_1227 ();
 sg13g2_decap_8 FILLER_182_1234 ();
 sg13g2_decap_8 FILLER_182_1241 ();
 sg13g2_decap_8 FILLER_182_1248 ();
 sg13g2_decap_8 FILLER_182_1255 ();
 sg13g2_decap_8 FILLER_182_1262 ();
 sg13g2_decap_8 FILLER_182_1269 ();
 sg13g2_decap_8 FILLER_182_1276 ();
 sg13g2_decap_8 FILLER_182_1283 ();
 sg13g2_decap_8 FILLER_182_1290 ();
 sg13g2_decap_8 FILLER_182_1297 ();
 sg13g2_decap_8 FILLER_182_1304 ();
 sg13g2_decap_8 FILLER_182_1311 ();
 sg13g2_decap_8 FILLER_182_1318 ();
 sg13g2_decap_8 FILLER_182_1325 ();
 sg13g2_decap_8 FILLER_182_1332 ();
 sg13g2_decap_8 FILLER_182_1339 ();
 sg13g2_decap_8 FILLER_182_1346 ();
 sg13g2_decap_8 FILLER_182_1353 ();
 sg13g2_decap_8 FILLER_182_1360 ();
 sg13g2_decap_8 FILLER_182_1367 ();
 sg13g2_decap_8 FILLER_182_1374 ();
 sg13g2_decap_8 FILLER_182_1381 ();
 sg13g2_decap_8 FILLER_182_1388 ();
 sg13g2_decap_8 FILLER_182_1395 ();
 sg13g2_decap_8 FILLER_182_1402 ();
 sg13g2_decap_8 FILLER_182_1409 ();
 sg13g2_decap_8 FILLER_182_1416 ();
 sg13g2_decap_8 FILLER_182_1423 ();
 sg13g2_decap_8 FILLER_182_1430 ();
 sg13g2_decap_8 FILLER_182_1437 ();
 sg13g2_decap_8 FILLER_182_1444 ();
 sg13g2_decap_8 FILLER_182_1451 ();
 sg13g2_decap_8 FILLER_182_1458 ();
 sg13g2_decap_8 FILLER_182_1465 ();
 sg13g2_decap_8 FILLER_182_1472 ();
 sg13g2_decap_8 FILLER_182_1479 ();
 sg13g2_decap_8 FILLER_182_1486 ();
 sg13g2_decap_8 FILLER_182_1493 ();
 sg13g2_decap_8 FILLER_182_1500 ();
 sg13g2_decap_8 FILLER_182_1507 ();
 sg13g2_decap_8 FILLER_182_1514 ();
 sg13g2_decap_8 FILLER_182_1521 ();
 sg13g2_decap_8 FILLER_182_1528 ();
 sg13g2_decap_8 FILLER_182_1535 ();
 sg13g2_decap_8 FILLER_182_1542 ();
 sg13g2_decap_8 FILLER_182_1549 ();
 sg13g2_decap_8 FILLER_182_1556 ();
 sg13g2_decap_8 FILLER_182_1563 ();
 sg13g2_decap_8 FILLER_182_1570 ();
 sg13g2_decap_8 FILLER_182_1577 ();
 sg13g2_decap_8 FILLER_182_1584 ();
 sg13g2_decap_8 FILLER_182_1591 ();
 sg13g2_decap_8 FILLER_182_1598 ();
 sg13g2_decap_8 FILLER_182_1605 ();
 sg13g2_decap_8 FILLER_182_1612 ();
 sg13g2_decap_8 FILLER_182_1619 ();
 sg13g2_decap_8 FILLER_182_1626 ();
 sg13g2_decap_8 FILLER_182_1633 ();
 sg13g2_decap_8 FILLER_182_1640 ();
 sg13g2_decap_8 FILLER_182_1647 ();
 sg13g2_decap_8 FILLER_182_1654 ();
 sg13g2_decap_8 FILLER_182_1661 ();
 sg13g2_decap_8 FILLER_182_1668 ();
 sg13g2_decap_8 FILLER_182_1675 ();
 sg13g2_decap_8 FILLER_182_1682 ();
 sg13g2_decap_8 FILLER_182_1689 ();
 sg13g2_decap_8 FILLER_182_1696 ();
 sg13g2_decap_8 FILLER_182_1703 ();
 sg13g2_decap_8 FILLER_182_1710 ();
 sg13g2_decap_8 FILLER_182_1717 ();
 sg13g2_decap_8 FILLER_182_1724 ();
 sg13g2_decap_8 FILLER_182_1731 ();
 sg13g2_decap_8 FILLER_182_1738 ();
 sg13g2_decap_8 FILLER_182_1745 ();
 sg13g2_decap_8 FILLER_182_1752 ();
 sg13g2_decap_8 FILLER_182_1759 ();
 sg13g2_fill_2 FILLER_182_1766 ();
 sg13g2_decap_8 FILLER_183_0 ();
 sg13g2_decap_8 FILLER_183_7 ();
 sg13g2_decap_8 FILLER_183_14 ();
 sg13g2_decap_8 FILLER_183_21 ();
 sg13g2_decap_8 FILLER_183_28 ();
 sg13g2_decap_8 FILLER_183_35 ();
 sg13g2_decap_8 FILLER_183_42 ();
 sg13g2_decap_8 FILLER_183_49 ();
 sg13g2_decap_8 FILLER_183_56 ();
 sg13g2_decap_8 FILLER_183_63 ();
 sg13g2_decap_8 FILLER_183_70 ();
 sg13g2_decap_8 FILLER_183_77 ();
 sg13g2_decap_8 FILLER_183_84 ();
 sg13g2_decap_8 FILLER_183_91 ();
 sg13g2_decap_8 FILLER_183_98 ();
 sg13g2_decap_8 FILLER_183_105 ();
 sg13g2_decap_8 FILLER_183_112 ();
 sg13g2_decap_8 FILLER_183_119 ();
 sg13g2_decap_8 FILLER_183_126 ();
 sg13g2_decap_8 FILLER_183_133 ();
 sg13g2_decap_8 FILLER_183_140 ();
 sg13g2_decap_8 FILLER_183_147 ();
 sg13g2_decap_8 FILLER_183_154 ();
 sg13g2_decap_8 FILLER_183_161 ();
 sg13g2_decap_8 FILLER_183_168 ();
 sg13g2_decap_8 FILLER_183_175 ();
 sg13g2_decap_8 FILLER_183_182 ();
 sg13g2_decap_8 FILLER_183_189 ();
 sg13g2_decap_8 FILLER_183_196 ();
 sg13g2_decap_8 FILLER_183_203 ();
 sg13g2_decap_8 FILLER_183_210 ();
 sg13g2_decap_8 FILLER_183_217 ();
 sg13g2_decap_8 FILLER_183_224 ();
 sg13g2_decap_8 FILLER_183_231 ();
 sg13g2_decap_8 FILLER_183_238 ();
 sg13g2_decap_8 FILLER_183_245 ();
 sg13g2_decap_8 FILLER_183_252 ();
 sg13g2_decap_8 FILLER_183_259 ();
 sg13g2_decap_8 FILLER_183_266 ();
 sg13g2_decap_8 FILLER_183_273 ();
 sg13g2_decap_8 FILLER_183_280 ();
 sg13g2_decap_8 FILLER_183_287 ();
 sg13g2_decap_8 FILLER_183_294 ();
 sg13g2_decap_8 FILLER_183_301 ();
 sg13g2_decap_8 FILLER_183_308 ();
 sg13g2_decap_8 FILLER_183_315 ();
 sg13g2_decap_8 FILLER_183_322 ();
 sg13g2_decap_8 FILLER_183_329 ();
 sg13g2_decap_4 FILLER_183_336 ();
 sg13g2_fill_1 FILLER_183_340 ();
 sg13g2_decap_8 FILLER_183_345 ();
 sg13g2_decap_8 FILLER_183_352 ();
 sg13g2_decap_8 FILLER_183_359 ();
 sg13g2_decap_8 FILLER_183_366 ();
 sg13g2_decap_8 FILLER_183_373 ();
 sg13g2_decap_8 FILLER_183_380 ();
 sg13g2_decap_4 FILLER_183_387 ();
 sg13g2_decap_8 FILLER_183_417 ();
 sg13g2_decap_4 FILLER_183_424 ();
 sg13g2_fill_1 FILLER_183_428 ();
 sg13g2_decap_8 FILLER_183_454 ();
 sg13g2_decap_4 FILLER_183_461 ();
 sg13g2_fill_1 FILLER_183_465 ();
 sg13g2_decap_8 FILLER_183_470 ();
 sg13g2_decap_8 FILLER_183_477 ();
 sg13g2_decap_8 FILLER_183_484 ();
 sg13g2_decap_8 FILLER_183_491 ();
 sg13g2_decap_8 FILLER_183_498 ();
 sg13g2_decap_8 FILLER_183_505 ();
 sg13g2_decap_8 FILLER_183_512 ();
 sg13g2_decap_8 FILLER_183_519 ();
 sg13g2_decap_8 FILLER_183_526 ();
 sg13g2_decap_8 FILLER_183_533 ();
 sg13g2_decap_8 FILLER_183_540 ();
 sg13g2_decap_8 FILLER_183_547 ();
 sg13g2_decap_8 FILLER_183_554 ();
 sg13g2_decap_8 FILLER_183_561 ();
 sg13g2_decap_8 FILLER_183_568 ();
 sg13g2_decap_8 FILLER_183_575 ();
 sg13g2_decap_8 FILLER_183_582 ();
 sg13g2_decap_8 FILLER_183_589 ();
 sg13g2_decap_8 FILLER_183_596 ();
 sg13g2_decap_8 FILLER_183_603 ();
 sg13g2_decap_8 FILLER_183_610 ();
 sg13g2_decap_8 FILLER_183_617 ();
 sg13g2_decap_8 FILLER_183_624 ();
 sg13g2_decap_8 FILLER_183_631 ();
 sg13g2_decap_8 FILLER_183_638 ();
 sg13g2_decap_8 FILLER_183_645 ();
 sg13g2_decap_8 FILLER_183_652 ();
 sg13g2_decap_8 FILLER_183_659 ();
 sg13g2_decap_8 FILLER_183_666 ();
 sg13g2_decap_8 FILLER_183_673 ();
 sg13g2_decap_8 FILLER_183_680 ();
 sg13g2_decap_8 FILLER_183_687 ();
 sg13g2_decap_8 FILLER_183_694 ();
 sg13g2_decap_8 FILLER_183_701 ();
 sg13g2_decap_8 FILLER_183_708 ();
 sg13g2_decap_8 FILLER_183_715 ();
 sg13g2_decap_8 FILLER_183_722 ();
 sg13g2_decap_8 FILLER_183_729 ();
 sg13g2_decap_8 FILLER_183_736 ();
 sg13g2_decap_8 FILLER_183_743 ();
 sg13g2_decap_8 FILLER_183_750 ();
 sg13g2_decap_8 FILLER_183_757 ();
 sg13g2_decap_8 FILLER_183_764 ();
 sg13g2_decap_8 FILLER_183_771 ();
 sg13g2_decap_8 FILLER_183_778 ();
 sg13g2_decap_8 FILLER_183_785 ();
 sg13g2_decap_8 FILLER_183_792 ();
 sg13g2_decap_8 FILLER_183_799 ();
 sg13g2_decap_8 FILLER_183_806 ();
 sg13g2_decap_8 FILLER_183_813 ();
 sg13g2_decap_8 FILLER_183_820 ();
 sg13g2_decap_8 FILLER_183_827 ();
 sg13g2_decap_8 FILLER_183_834 ();
 sg13g2_decap_8 FILLER_183_841 ();
 sg13g2_decap_8 FILLER_183_848 ();
 sg13g2_decap_8 FILLER_183_855 ();
 sg13g2_decap_8 FILLER_183_862 ();
 sg13g2_decap_8 FILLER_183_869 ();
 sg13g2_decap_8 FILLER_183_876 ();
 sg13g2_decap_8 FILLER_183_883 ();
 sg13g2_decap_8 FILLER_183_890 ();
 sg13g2_decap_8 FILLER_183_897 ();
 sg13g2_decap_8 FILLER_183_904 ();
 sg13g2_decap_8 FILLER_183_911 ();
 sg13g2_decap_8 FILLER_183_918 ();
 sg13g2_decap_8 FILLER_183_925 ();
 sg13g2_decap_8 FILLER_183_932 ();
 sg13g2_decap_8 FILLER_183_939 ();
 sg13g2_decap_8 FILLER_183_946 ();
 sg13g2_decap_8 FILLER_183_953 ();
 sg13g2_decap_8 FILLER_183_960 ();
 sg13g2_decap_8 FILLER_183_967 ();
 sg13g2_decap_8 FILLER_183_974 ();
 sg13g2_decap_8 FILLER_183_981 ();
 sg13g2_decap_8 FILLER_183_988 ();
 sg13g2_decap_8 FILLER_183_995 ();
 sg13g2_decap_8 FILLER_183_1002 ();
 sg13g2_decap_8 FILLER_183_1009 ();
 sg13g2_decap_8 FILLER_183_1016 ();
 sg13g2_decap_8 FILLER_183_1023 ();
 sg13g2_decap_8 FILLER_183_1030 ();
 sg13g2_decap_8 FILLER_183_1037 ();
 sg13g2_decap_8 FILLER_183_1044 ();
 sg13g2_decap_8 FILLER_183_1051 ();
 sg13g2_decap_8 FILLER_183_1058 ();
 sg13g2_decap_8 FILLER_183_1065 ();
 sg13g2_decap_8 FILLER_183_1072 ();
 sg13g2_decap_8 FILLER_183_1079 ();
 sg13g2_decap_8 FILLER_183_1086 ();
 sg13g2_decap_8 FILLER_183_1093 ();
 sg13g2_decap_8 FILLER_183_1100 ();
 sg13g2_decap_8 FILLER_183_1107 ();
 sg13g2_decap_8 FILLER_183_1114 ();
 sg13g2_decap_8 FILLER_183_1121 ();
 sg13g2_decap_8 FILLER_183_1128 ();
 sg13g2_decap_8 FILLER_183_1135 ();
 sg13g2_decap_8 FILLER_183_1142 ();
 sg13g2_decap_8 FILLER_183_1149 ();
 sg13g2_decap_8 FILLER_183_1156 ();
 sg13g2_decap_8 FILLER_183_1163 ();
 sg13g2_decap_8 FILLER_183_1170 ();
 sg13g2_decap_8 FILLER_183_1177 ();
 sg13g2_decap_8 FILLER_183_1184 ();
 sg13g2_decap_8 FILLER_183_1191 ();
 sg13g2_decap_8 FILLER_183_1198 ();
 sg13g2_decap_8 FILLER_183_1205 ();
 sg13g2_decap_8 FILLER_183_1212 ();
 sg13g2_decap_8 FILLER_183_1219 ();
 sg13g2_decap_8 FILLER_183_1226 ();
 sg13g2_decap_8 FILLER_183_1233 ();
 sg13g2_decap_8 FILLER_183_1240 ();
 sg13g2_decap_8 FILLER_183_1247 ();
 sg13g2_decap_8 FILLER_183_1254 ();
 sg13g2_decap_8 FILLER_183_1261 ();
 sg13g2_decap_8 FILLER_183_1268 ();
 sg13g2_decap_8 FILLER_183_1275 ();
 sg13g2_decap_8 FILLER_183_1282 ();
 sg13g2_decap_8 FILLER_183_1289 ();
 sg13g2_decap_8 FILLER_183_1296 ();
 sg13g2_decap_8 FILLER_183_1303 ();
 sg13g2_decap_8 FILLER_183_1310 ();
 sg13g2_decap_8 FILLER_183_1317 ();
 sg13g2_decap_8 FILLER_183_1324 ();
 sg13g2_decap_8 FILLER_183_1331 ();
 sg13g2_decap_8 FILLER_183_1338 ();
 sg13g2_decap_8 FILLER_183_1345 ();
 sg13g2_decap_8 FILLER_183_1352 ();
 sg13g2_decap_8 FILLER_183_1359 ();
 sg13g2_decap_8 FILLER_183_1366 ();
 sg13g2_decap_8 FILLER_183_1373 ();
 sg13g2_decap_8 FILLER_183_1380 ();
 sg13g2_decap_8 FILLER_183_1387 ();
 sg13g2_decap_8 FILLER_183_1394 ();
 sg13g2_decap_8 FILLER_183_1401 ();
 sg13g2_decap_8 FILLER_183_1408 ();
 sg13g2_decap_8 FILLER_183_1415 ();
 sg13g2_decap_8 FILLER_183_1422 ();
 sg13g2_decap_8 FILLER_183_1429 ();
 sg13g2_decap_8 FILLER_183_1436 ();
 sg13g2_decap_8 FILLER_183_1443 ();
 sg13g2_decap_8 FILLER_183_1450 ();
 sg13g2_decap_8 FILLER_183_1457 ();
 sg13g2_decap_8 FILLER_183_1464 ();
 sg13g2_decap_8 FILLER_183_1471 ();
 sg13g2_decap_8 FILLER_183_1478 ();
 sg13g2_decap_8 FILLER_183_1485 ();
 sg13g2_decap_8 FILLER_183_1492 ();
 sg13g2_decap_8 FILLER_183_1499 ();
 sg13g2_decap_8 FILLER_183_1506 ();
 sg13g2_decap_8 FILLER_183_1513 ();
 sg13g2_decap_8 FILLER_183_1520 ();
 sg13g2_decap_8 FILLER_183_1527 ();
 sg13g2_decap_8 FILLER_183_1534 ();
 sg13g2_decap_8 FILLER_183_1541 ();
 sg13g2_decap_8 FILLER_183_1548 ();
 sg13g2_decap_8 FILLER_183_1555 ();
 sg13g2_decap_8 FILLER_183_1562 ();
 sg13g2_decap_8 FILLER_183_1569 ();
 sg13g2_decap_8 FILLER_183_1576 ();
 sg13g2_decap_8 FILLER_183_1583 ();
 sg13g2_decap_8 FILLER_183_1590 ();
 sg13g2_decap_8 FILLER_183_1597 ();
 sg13g2_decap_8 FILLER_183_1604 ();
 sg13g2_decap_8 FILLER_183_1611 ();
 sg13g2_decap_8 FILLER_183_1618 ();
 sg13g2_decap_8 FILLER_183_1625 ();
 sg13g2_decap_8 FILLER_183_1632 ();
 sg13g2_decap_8 FILLER_183_1639 ();
 sg13g2_decap_8 FILLER_183_1646 ();
 sg13g2_decap_8 FILLER_183_1653 ();
 sg13g2_decap_8 FILLER_183_1660 ();
 sg13g2_decap_8 FILLER_183_1667 ();
 sg13g2_decap_8 FILLER_183_1674 ();
 sg13g2_decap_8 FILLER_183_1681 ();
 sg13g2_decap_8 FILLER_183_1688 ();
 sg13g2_decap_8 FILLER_183_1695 ();
 sg13g2_decap_8 FILLER_183_1702 ();
 sg13g2_decap_8 FILLER_183_1709 ();
 sg13g2_decap_8 FILLER_183_1716 ();
 sg13g2_decap_8 FILLER_183_1723 ();
 sg13g2_decap_8 FILLER_183_1730 ();
 sg13g2_decap_8 FILLER_183_1737 ();
 sg13g2_decap_8 FILLER_183_1744 ();
 sg13g2_decap_8 FILLER_183_1751 ();
 sg13g2_decap_8 FILLER_183_1758 ();
 sg13g2_fill_2 FILLER_183_1765 ();
 sg13g2_fill_1 FILLER_183_1767 ();
 sg13g2_decap_8 FILLER_184_0 ();
 sg13g2_decap_8 FILLER_184_7 ();
 sg13g2_decap_8 FILLER_184_14 ();
 sg13g2_decap_8 FILLER_184_21 ();
 sg13g2_decap_8 FILLER_184_28 ();
 sg13g2_decap_8 FILLER_184_35 ();
 sg13g2_decap_8 FILLER_184_42 ();
 sg13g2_decap_8 FILLER_184_49 ();
 sg13g2_decap_8 FILLER_184_56 ();
 sg13g2_decap_8 FILLER_184_63 ();
 sg13g2_decap_8 FILLER_184_70 ();
 sg13g2_decap_8 FILLER_184_77 ();
 sg13g2_decap_8 FILLER_184_84 ();
 sg13g2_decap_8 FILLER_184_91 ();
 sg13g2_decap_8 FILLER_184_98 ();
 sg13g2_decap_8 FILLER_184_105 ();
 sg13g2_decap_8 FILLER_184_112 ();
 sg13g2_decap_8 FILLER_184_119 ();
 sg13g2_decap_8 FILLER_184_126 ();
 sg13g2_decap_8 FILLER_184_133 ();
 sg13g2_decap_8 FILLER_184_140 ();
 sg13g2_decap_8 FILLER_184_147 ();
 sg13g2_decap_8 FILLER_184_154 ();
 sg13g2_decap_8 FILLER_184_161 ();
 sg13g2_decap_8 FILLER_184_168 ();
 sg13g2_decap_8 FILLER_184_175 ();
 sg13g2_decap_8 FILLER_184_182 ();
 sg13g2_decap_8 FILLER_184_189 ();
 sg13g2_decap_8 FILLER_184_196 ();
 sg13g2_decap_8 FILLER_184_203 ();
 sg13g2_decap_8 FILLER_184_210 ();
 sg13g2_decap_8 FILLER_184_217 ();
 sg13g2_decap_8 FILLER_184_224 ();
 sg13g2_decap_8 FILLER_184_231 ();
 sg13g2_decap_8 FILLER_184_238 ();
 sg13g2_decap_8 FILLER_184_245 ();
 sg13g2_decap_8 FILLER_184_252 ();
 sg13g2_decap_8 FILLER_184_259 ();
 sg13g2_decap_8 FILLER_184_266 ();
 sg13g2_decap_8 FILLER_184_273 ();
 sg13g2_decap_8 FILLER_184_280 ();
 sg13g2_decap_8 FILLER_184_287 ();
 sg13g2_decap_8 FILLER_184_294 ();
 sg13g2_decap_8 FILLER_184_301 ();
 sg13g2_decap_8 FILLER_184_308 ();
 sg13g2_decap_8 FILLER_184_315 ();
 sg13g2_decap_8 FILLER_184_322 ();
 sg13g2_decap_8 FILLER_184_329 ();
 sg13g2_decap_8 FILLER_184_336 ();
 sg13g2_decap_8 FILLER_184_343 ();
 sg13g2_decap_8 FILLER_184_350 ();
 sg13g2_decap_8 FILLER_184_357 ();
 sg13g2_decap_8 FILLER_184_364 ();
 sg13g2_decap_8 FILLER_184_371 ();
 sg13g2_decap_8 FILLER_184_378 ();
 sg13g2_decap_8 FILLER_184_385 ();
 sg13g2_decap_8 FILLER_184_392 ();
 sg13g2_decap_8 FILLER_184_399 ();
 sg13g2_decap_8 FILLER_184_406 ();
 sg13g2_decap_8 FILLER_184_413 ();
 sg13g2_decap_8 FILLER_184_420 ();
 sg13g2_decap_8 FILLER_184_427 ();
 sg13g2_decap_8 FILLER_184_434 ();
 sg13g2_decap_8 FILLER_184_441 ();
 sg13g2_decap_8 FILLER_184_448 ();
 sg13g2_decap_8 FILLER_184_455 ();
 sg13g2_decap_8 FILLER_184_462 ();
 sg13g2_decap_8 FILLER_184_469 ();
 sg13g2_decap_8 FILLER_184_476 ();
 sg13g2_decap_8 FILLER_184_483 ();
 sg13g2_decap_8 FILLER_184_490 ();
 sg13g2_decap_8 FILLER_184_497 ();
 sg13g2_decap_8 FILLER_184_504 ();
 sg13g2_decap_8 FILLER_184_511 ();
 sg13g2_decap_8 FILLER_184_518 ();
 sg13g2_decap_8 FILLER_184_525 ();
 sg13g2_decap_8 FILLER_184_532 ();
 sg13g2_decap_8 FILLER_184_539 ();
 sg13g2_decap_8 FILLER_184_546 ();
 sg13g2_decap_8 FILLER_184_553 ();
 sg13g2_decap_8 FILLER_184_560 ();
 sg13g2_decap_8 FILLER_184_567 ();
 sg13g2_decap_8 FILLER_184_574 ();
 sg13g2_decap_8 FILLER_184_581 ();
 sg13g2_decap_8 FILLER_184_588 ();
 sg13g2_decap_8 FILLER_184_595 ();
 sg13g2_decap_8 FILLER_184_602 ();
 sg13g2_decap_8 FILLER_184_609 ();
 sg13g2_decap_8 FILLER_184_616 ();
 sg13g2_decap_8 FILLER_184_623 ();
 sg13g2_decap_8 FILLER_184_630 ();
 sg13g2_decap_8 FILLER_184_637 ();
 sg13g2_decap_8 FILLER_184_644 ();
 sg13g2_decap_8 FILLER_184_651 ();
 sg13g2_decap_8 FILLER_184_658 ();
 sg13g2_decap_8 FILLER_184_665 ();
 sg13g2_decap_8 FILLER_184_672 ();
 sg13g2_decap_8 FILLER_184_679 ();
 sg13g2_decap_8 FILLER_184_686 ();
 sg13g2_decap_8 FILLER_184_693 ();
 sg13g2_decap_8 FILLER_184_700 ();
 sg13g2_decap_8 FILLER_184_707 ();
 sg13g2_decap_8 FILLER_184_714 ();
 sg13g2_decap_8 FILLER_184_721 ();
 sg13g2_decap_8 FILLER_184_728 ();
 sg13g2_decap_8 FILLER_184_735 ();
 sg13g2_decap_8 FILLER_184_742 ();
 sg13g2_decap_8 FILLER_184_749 ();
 sg13g2_decap_8 FILLER_184_756 ();
 sg13g2_decap_8 FILLER_184_763 ();
 sg13g2_decap_8 FILLER_184_770 ();
 sg13g2_decap_8 FILLER_184_777 ();
 sg13g2_decap_8 FILLER_184_784 ();
 sg13g2_decap_8 FILLER_184_791 ();
 sg13g2_decap_8 FILLER_184_798 ();
 sg13g2_decap_8 FILLER_184_805 ();
 sg13g2_decap_8 FILLER_184_812 ();
 sg13g2_decap_8 FILLER_184_819 ();
 sg13g2_decap_8 FILLER_184_826 ();
 sg13g2_decap_8 FILLER_184_833 ();
 sg13g2_decap_8 FILLER_184_840 ();
 sg13g2_decap_8 FILLER_184_847 ();
 sg13g2_decap_8 FILLER_184_854 ();
 sg13g2_decap_8 FILLER_184_861 ();
 sg13g2_decap_8 FILLER_184_868 ();
 sg13g2_decap_8 FILLER_184_875 ();
 sg13g2_decap_8 FILLER_184_882 ();
 sg13g2_decap_8 FILLER_184_889 ();
 sg13g2_decap_8 FILLER_184_896 ();
 sg13g2_decap_8 FILLER_184_903 ();
 sg13g2_decap_8 FILLER_184_910 ();
 sg13g2_decap_8 FILLER_184_917 ();
 sg13g2_decap_8 FILLER_184_924 ();
 sg13g2_decap_8 FILLER_184_931 ();
 sg13g2_decap_8 FILLER_184_938 ();
 sg13g2_decap_8 FILLER_184_945 ();
 sg13g2_decap_8 FILLER_184_952 ();
 sg13g2_decap_8 FILLER_184_959 ();
 sg13g2_decap_8 FILLER_184_966 ();
 sg13g2_decap_8 FILLER_184_973 ();
 sg13g2_decap_8 FILLER_184_980 ();
 sg13g2_decap_8 FILLER_184_987 ();
 sg13g2_decap_8 FILLER_184_994 ();
 sg13g2_decap_8 FILLER_184_1001 ();
 sg13g2_decap_8 FILLER_184_1008 ();
 sg13g2_decap_8 FILLER_184_1015 ();
 sg13g2_decap_8 FILLER_184_1022 ();
 sg13g2_decap_8 FILLER_184_1029 ();
 sg13g2_decap_8 FILLER_184_1036 ();
 sg13g2_decap_8 FILLER_184_1043 ();
 sg13g2_decap_8 FILLER_184_1050 ();
 sg13g2_decap_8 FILLER_184_1057 ();
 sg13g2_decap_8 FILLER_184_1064 ();
 sg13g2_decap_8 FILLER_184_1071 ();
 sg13g2_decap_8 FILLER_184_1078 ();
 sg13g2_decap_8 FILLER_184_1085 ();
 sg13g2_decap_8 FILLER_184_1092 ();
 sg13g2_decap_8 FILLER_184_1099 ();
 sg13g2_decap_8 FILLER_184_1106 ();
 sg13g2_decap_8 FILLER_184_1113 ();
 sg13g2_decap_8 FILLER_184_1120 ();
 sg13g2_decap_8 FILLER_184_1127 ();
 sg13g2_decap_8 FILLER_184_1134 ();
 sg13g2_decap_8 FILLER_184_1141 ();
 sg13g2_decap_8 FILLER_184_1148 ();
 sg13g2_decap_8 FILLER_184_1155 ();
 sg13g2_decap_8 FILLER_184_1162 ();
 sg13g2_decap_8 FILLER_184_1169 ();
 sg13g2_decap_8 FILLER_184_1176 ();
 sg13g2_decap_8 FILLER_184_1183 ();
 sg13g2_decap_8 FILLER_184_1190 ();
 sg13g2_decap_8 FILLER_184_1197 ();
 sg13g2_decap_8 FILLER_184_1204 ();
 sg13g2_decap_8 FILLER_184_1211 ();
 sg13g2_decap_8 FILLER_184_1218 ();
 sg13g2_decap_8 FILLER_184_1225 ();
 sg13g2_decap_8 FILLER_184_1232 ();
 sg13g2_decap_8 FILLER_184_1239 ();
 sg13g2_decap_8 FILLER_184_1246 ();
 sg13g2_decap_8 FILLER_184_1253 ();
 sg13g2_decap_8 FILLER_184_1260 ();
 sg13g2_decap_8 FILLER_184_1267 ();
 sg13g2_decap_8 FILLER_184_1274 ();
 sg13g2_decap_8 FILLER_184_1281 ();
 sg13g2_decap_8 FILLER_184_1288 ();
 sg13g2_decap_8 FILLER_184_1295 ();
 sg13g2_decap_8 FILLER_184_1302 ();
 sg13g2_decap_8 FILLER_184_1309 ();
 sg13g2_decap_8 FILLER_184_1316 ();
 sg13g2_decap_8 FILLER_184_1323 ();
 sg13g2_decap_8 FILLER_184_1330 ();
 sg13g2_decap_8 FILLER_184_1337 ();
 sg13g2_decap_8 FILLER_184_1344 ();
 sg13g2_decap_8 FILLER_184_1351 ();
 sg13g2_decap_8 FILLER_184_1358 ();
 sg13g2_decap_8 FILLER_184_1365 ();
 sg13g2_decap_8 FILLER_184_1372 ();
 sg13g2_decap_8 FILLER_184_1379 ();
 sg13g2_decap_8 FILLER_184_1386 ();
 sg13g2_decap_8 FILLER_184_1393 ();
 sg13g2_decap_8 FILLER_184_1400 ();
 sg13g2_decap_8 FILLER_184_1407 ();
 sg13g2_decap_8 FILLER_184_1414 ();
 sg13g2_decap_8 FILLER_184_1421 ();
 sg13g2_decap_8 FILLER_184_1428 ();
 sg13g2_decap_8 FILLER_184_1435 ();
 sg13g2_decap_8 FILLER_184_1442 ();
 sg13g2_decap_8 FILLER_184_1449 ();
 sg13g2_decap_8 FILLER_184_1456 ();
 sg13g2_decap_8 FILLER_184_1463 ();
 sg13g2_decap_8 FILLER_184_1470 ();
 sg13g2_decap_8 FILLER_184_1477 ();
 sg13g2_decap_8 FILLER_184_1484 ();
 sg13g2_decap_8 FILLER_184_1491 ();
 sg13g2_decap_8 FILLER_184_1498 ();
 sg13g2_decap_8 FILLER_184_1505 ();
 sg13g2_decap_8 FILLER_184_1512 ();
 sg13g2_decap_8 FILLER_184_1519 ();
 sg13g2_decap_8 FILLER_184_1526 ();
 sg13g2_decap_8 FILLER_184_1533 ();
 sg13g2_decap_8 FILLER_184_1540 ();
 sg13g2_decap_8 FILLER_184_1547 ();
 sg13g2_decap_8 FILLER_184_1554 ();
 sg13g2_decap_8 FILLER_184_1561 ();
 sg13g2_decap_8 FILLER_184_1568 ();
 sg13g2_decap_8 FILLER_184_1575 ();
 sg13g2_decap_8 FILLER_184_1582 ();
 sg13g2_decap_8 FILLER_184_1589 ();
 sg13g2_decap_8 FILLER_184_1596 ();
 sg13g2_decap_8 FILLER_184_1603 ();
 sg13g2_decap_8 FILLER_184_1610 ();
 sg13g2_decap_8 FILLER_184_1617 ();
 sg13g2_decap_8 FILLER_184_1624 ();
 sg13g2_decap_8 FILLER_184_1631 ();
 sg13g2_decap_8 FILLER_184_1638 ();
 sg13g2_decap_8 FILLER_184_1645 ();
 sg13g2_decap_8 FILLER_184_1652 ();
 sg13g2_decap_8 FILLER_184_1659 ();
 sg13g2_decap_8 FILLER_184_1666 ();
 sg13g2_decap_8 FILLER_184_1673 ();
 sg13g2_decap_8 FILLER_184_1680 ();
 sg13g2_decap_8 FILLER_184_1687 ();
 sg13g2_decap_8 FILLER_184_1694 ();
 sg13g2_decap_8 FILLER_184_1701 ();
 sg13g2_decap_8 FILLER_184_1708 ();
 sg13g2_decap_8 FILLER_184_1715 ();
 sg13g2_decap_8 FILLER_184_1722 ();
 sg13g2_decap_8 FILLER_184_1729 ();
 sg13g2_decap_8 FILLER_184_1736 ();
 sg13g2_decap_8 FILLER_184_1743 ();
 sg13g2_decap_8 FILLER_184_1750 ();
 sg13g2_decap_8 FILLER_184_1757 ();
 sg13g2_decap_4 FILLER_184_1764 ();
 sg13g2_decap_8 FILLER_185_0 ();
 sg13g2_decap_8 FILLER_185_7 ();
 sg13g2_decap_8 FILLER_185_14 ();
 sg13g2_decap_8 FILLER_185_21 ();
 sg13g2_decap_8 FILLER_185_28 ();
 sg13g2_decap_8 FILLER_185_35 ();
 sg13g2_decap_8 FILLER_185_42 ();
 sg13g2_decap_8 FILLER_185_49 ();
 sg13g2_decap_4 FILLER_185_60 ();
 sg13g2_decap_4 FILLER_185_68 ();
 sg13g2_decap_4 FILLER_185_76 ();
 sg13g2_decap_4 FILLER_185_84 ();
 sg13g2_decap_4 FILLER_185_92 ();
 sg13g2_decap_4 FILLER_185_100 ();
 sg13g2_decap_4 FILLER_185_108 ();
 sg13g2_decap_4 FILLER_185_116 ();
 sg13g2_decap_8 FILLER_185_124 ();
 sg13g2_decap_8 FILLER_185_131 ();
 sg13g2_decap_8 FILLER_185_138 ();
 sg13g2_decap_8 FILLER_185_145 ();
 sg13g2_decap_8 FILLER_185_152 ();
 sg13g2_decap_8 FILLER_185_159 ();
 sg13g2_decap_8 FILLER_185_166 ();
 sg13g2_decap_8 FILLER_185_173 ();
 sg13g2_decap_8 FILLER_185_180 ();
 sg13g2_decap_8 FILLER_185_187 ();
 sg13g2_decap_8 FILLER_185_194 ();
 sg13g2_decap_8 FILLER_185_201 ();
 sg13g2_decap_8 FILLER_185_208 ();
 sg13g2_decap_8 FILLER_185_215 ();
 sg13g2_decap_8 FILLER_185_222 ();
 sg13g2_decap_8 FILLER_185_229 ();
 sg13g2_decap_8 FILLER_185_236 ();
 sg13g2_decap_8 FILLER_185_243 ();
 sg13g2_decap_8 FILLER_185_250 ();
 sg13g2_decap_8 FILLER_185_257 ();
 sg13g2_decap_8 FILLER_185_264 ();
 sg13g2_decap_8 FILLER_185_271 ();
 sg13g2_decap_8 FILLER_185_278 ();
 sg13g2_decap_8 FILLER_185_285 ();
 sg13g2_decap_8 FILLER_185_292 ();
 sg13g2_decap_8 FILLER_185_299 ();
 sg13g2_decap_4 FILLER_185_306 ();
 sg13g2_fill_2 FILLER_185_310 ();
 sg13g2_decap_4 FILLER_185_316 ();
 sg13g2_decap_4 FILLER_185_324 ();
 sg13g2_decap_4 FILLER_185_332 ();
 sg13g2_fill_2 FILLER_185_341 ();
 sg13g2_fill_1 FILLER_185_343 ();
 sg13g2_decap_4 FILLER_185_348 ();
 sg13g2_fill_2 FILLER_185_357 ();
 sg13g2_fill_1 FILLER_185_359 ();
 sg13g2_fill_2 FILLER_185_365 ();
 sg13g2_fill_1 FILLER_185_367 ();
 sg13g2_decap_8 FILLER_185_372 ();
 sg13g2_decap_8 FILLER_185_379 ();
 sg13g2_decap_8 FILLER_185_386 ();
 sg13g2_decap_8 FILLER_185_393 ();
 sg13g2_decap_8 FILLER_185_400 ();
 sg13g2_decap_8 FILLER_185_407 ();
 sg13g2_decap_8 FILLER_185_414 ();
 sg13g2_decap_8 FILLER_185_421 ();
 sg13g2_decap_8 FILLER_185_428 ();
 sg13g2_decap_8 FILLER_185_435 ();
 sg13g2_decap_8 FILLER_185_442 ();
 sg13g2_decap_8 FILLER_185_449 ();
 sg13g2_decap_8 FILLER_185_456 ();
 sg13g2_decap_8 FILLER_185_463 ();
 sg13g2_decap_8 FILLER_185_470 ();
 sg13g2_decap_8 FILLER_185_477 ();
 sg13g2_decap_8 FILLER_185_484 ();
 sg13g2_decap_8 FILLER_185_491 ();
 sg13g2_decap_8 FILLER_185_498 ();
 sg13g2_decap_8 FILLER_185_505 ();
 sg13g2_decap_8 FILLER_185_512 ();
 sg13g2_decap_8 FILLER_185_519 ();
 sg13g2_decap_8 FILLER_185_526 ();
 sg13g2_decap_8 FILLER_185_533 ();
 sg13g2_decap_8 FILLER_185_540 ();
 sg13g2_decap_8 FILLER_185_547 ();
 sg13g2_decap_8 FILLER_185_554 ();
 sg13g2_decap_8 FILLER_185_561 ();
 sg13g2_decap_8 FILLER_185_568 ();
 sg13g2_decap_8 FILLER_185_575 ();
 sg13g2_decap_8 FILLER_185_582 ();
 sg13g2_decap_8 FILLER_185_589 ();
 sg13g2_decap_8 FILLER_185_596 ();
 sg13g2_decap_8 FILLER_185_603 ();
 sg13g2_decap_8 FILLER_185_610 ();
 sg13g2_decap_8 FILLER_185_617 ();
 sg13g2_decap_8 FILLER_185_624 ();
 sg13g2_decap_8 FILLER_185_631 ();
 sg13g2_decap_8 FILLER_185_638 ();
 sg13g2_decap_8 FILLER_185_645 ();
 sg13g2_decap_8 FILLER_185_652 ();
 sg13g2_decap_8 FILLER_185_659 ();
 sg13g2_decap_8 FILLER_185_666 ();
 sg13g2_decap_8 FILLER_185_673 ();
 sg13g2_decap_8 FILLER_185_680 ();
 sg13g2_decap_8 FILLER_185_687 ();
 sg13g2_decap_8 FILLER_185_694 ();
 sg13g2_decap_8 FILLER_185_701 ();
 sg13g2_decap_8 FILLER_185_708 ();
 sg13g2_decap_8 FILLER_185_715 ();
 sg13g2_decap_8 FILLER_185_722 ();
 sg13g2_decap_8 FILLER_185_729 ();
 sg13g2_decap_8 FILLER_185_736 ();
 sg13g2_decap_8 FILLER_185_743 ();
 sg13g2_decap_8 FILLER_185_750 ();
 sg13g2_decap_8 FILLER_185_757 ();
 sg13g2_decap_8 FILLER_185_764 ();
 sg13g2_decap_8 FILLER_185_771 ();
 sg13g2_decap_8 FILLER_185_778 ();
 sg13g2_decap_8 FILLER_185_785 ();
 sg13g2_decap_8 FILLER_185_792 ();
 sg13g2_decap_8 FILLER_185_799 ();
 sg13g2_decap_8 FILLER_185_806 ();
 sg13g2_decap_8 FILLER_185_813 ();
 sg13g2_decap_8 FILLER_185_820 ();
 sg13g2_decap_8 FILLER_185_827 ();
 sg13g2_decap_8 FILLER_185_834 ();
 sg13g2_decap_8 FILLER_185_841 ();
 sg13g2_decap_8 FILLER_185_848 ();
 sg13g2_decap_8 FILLER_185_855 ();
 sg13g2_decap_8 FILLER_185_862 ();
 sg13g2_decap_8 FILLER_185_869 ();
 sg13g2_decap_8 FILLER_185_876 ();
 sg13g2_decap_8 FILLER_185_883 ();
 sg13g2_decap_8 FILLER_185_890 ();
 sg13g2_decap_8 FILLER_185_897 ();
 sg13g2_decap_8 FILLER_185_904 ();
 sg13g2_decap_8 FILLER_185_911 ();
 sg13g2_decap_8 FILLER_185_918 ();
 sg13g2_decap_8 FILLER_185_925 ();
 sg13g2_decap_8 FILLER_185_932 ();
 sg13g2_decap_8 FILLER_185_939 ();
 sg13g2_decap_8 FILLER_185_946 ();
 sg13g2_decap_8 FILLER_185_953 ();
 sg13g2_decap_8 FILLER_185_960 ();
 sg13g2_decap_8 FILLER_185_967 ();
 sg13g2_decap_8 FILLER_185_974 ();
 sg13g2_decap_8 FILLER_185_981 ();
 sg13g2_decap_8 FILLER_185_988 ();
 sg13g2_decap_8 FILLER_185_995 ();
 sg13g2_decap_8 FILLER_185_1002 ();
 sg13g2_decap_8 FILLER_185_1009 ();
 sg13g2_decap_8 FILLER_185_1016 ();
 sg13g2_decap_8 FILLER_185_1023 ();
 sg13g2_decap_8 FILLER_185_1030 ();
 sg13g2_decap_8 FILLER_185_1037 ();
 sg13g2_decap_8 FILLER_185_1044 ();
 sg13g2_decap_8 FILLER_185_1051 ();
 sg13g2_decap_8 FILLER_185_1058 ();
 sg13g2_decap_8 FILLER_185_1065 ();
 sg13g2_decap_8 FILLER_185_1072 ();
 sg13g2_decap_8 FILLER_185_1079 ();
 sg13g2_decap_8 FILLER_185_1086 ();
 sg13g2_decap_8 FILLER_185_1093 ();
 sg13g2_decap_8 FILLER_185_1100 ();
 sg13g2_decap_8 FILLER_185_1107 ();
 sg13g2_decap_8 FILLER_185_1114 ();
 sg13g2_decap_8 FILLER_185_1121 ();
 sg13g2_decap_8 FILLER_185_1128 ();
 sg13g2_decap_8 FILLER_185_1135 ();
 sg13g2_decap_8 FILLER_185_1142 ();
 sg13g2_decap_8 FILLER_185_1149 ();
 sg13g2_decap_8 FILLER_185_1156 ();
 sg13g2_decap_8 FILLER_185_1163 ();
 sg13g2_decap_8 FILLER_185_1170 ();
 sg13g2_decap_8 FILLER_185_1177 ();
 sg13g2_decap_8 FILLER_185_1184 ();
 sg13g2_decap_8 FILLER_185_1191 ();
 sg13g2_decap_8 FILLER_185_1198 ();
 sg13g2_decap_8 FILLER_185_1205 ();
 sg13g2_decap_8 FILLER_185_1212 ();
 sg13g2_decap_8 FILLER_185_1219 ();
 sg13g2_decap_8 FILLER_185_1226 ();
 sg13g2_decap_8 FILLER_185_1233 ();
 sg13g2_decap_8 FILLER_185_1240 ();
 sg13g2_decap_8 FILLER_185_1247 ();
 sg13g2_decap_8 FILLER_185_1254 ();
 sg13g2_decap_8 FILLER_185_1261 ();
 sg13g2_decap_8 FILLER_185_1268 ();
 sg13g2_decap_8 FILLER_185_1275 ();
 sg13g2_decap_8 FILLER_185_1282 ();
 sg13g2_decap_8 FILLER_185_1289 ();
 sg13g2_decap_8 FILLER_185_1296 ();
 sg13g2_decap_8 FILLER_185_1303 ();
 sg13g2_decap_8 FILLER_185_1310 ();
 sg13g2_decap_8 FILLER_185_1317 ();
 sg13g2_decap_8 FILLER_185_1324 ();
 sg13g2_decap_8 FILLER_185_1331 ();
 sg13g2_decap_8 FILLER_185_1338 ();
 sg13g2_decap_8 FILLER_185_1345 ();
 sg13g2_decap_8 FILLER_185_1352 ();
 sg13g2_decap_8 FILLER_185_1359 ();
 sg13g2_decap_8 FILLER_185_1366 ();
 sg13g2_decap_8 FILLER_185_1373 ();
 sg13g2_decap_8 FILLER_185_1380 ();
 sg13g2_decap_8 FILLER_185_1387 ();
 sg13g2_decap_8 FILLER_185_1394 ();
 sg13g2_decap_8 FILLER_185_1401 ();
 sg13g2_decap_8 FILLER_185_1408 ();
 sg13g2_decap_8 FILLER_185_1415 ();
 sg13g2_decap_8 FILLER_185_1422 ();
 sg13g2_decap_8 FILLER_185_1429 ();
 sg13g2_decap_8 FILLER_185_1436 ();
 sg13g2_decap_8 FILLER_185_1443 ();
 sg13g2_decap_8 FILLER_185_1450 ();
 sg13g2_decap_8 FILLER_185_1457 ();
 sg13g2_decap_8 FILLER_185_1464 ();
 sg13g2_decap_8 FILLER_185_1471 ();
 sg13g2_decap_8 FILLER_185_1478 ();
 sg13g2_decap_8 FILLER_185_1485 ();
 sg13g2_decap_8 FILLER_185_1492 ();
 sg13g2_decap_8 FILLER_185_1499 ();
 sg13g2_decap_8 FILLER_185_1506 ();
 sg13g2_decap_8 FILLER_185_1513 ();
 sg13g2_decap_8 FILLER_185_1520 ();
 sg13g2_decap_8 FILLER_185_1527 ();
 sg13g2_decap_8 FILLER_185_1534 ();
 sg13g2_decap_8 FILLER_185_1541 ();
 sg13g2_decap_8 FILLER_185_1548 ();
 sg13g2_decap_8 FILLER_185_1555 ();
 sg13g2_decap_8 FILLER_185_1562 ();
 sg13g2_decap_8 FILLER_185_1569 ();
 sg13g2_decap_8 FILLER_185_1576 ();
 sg13g2_decap_8 FILLER_185_1583 ();
 sg13g2_decap_8 FILLER_185_1590 ();
 sg13g2_decap_8 FILLER_185_1597 ();
 sg13g2_decap_8 FILLER_185_1604 ();
 sg13g2_decap_8 FILLER_185_1611 ();
 sg13g2_decap_8 FILLER_185_1618 ();
 sg13g2_decap_8 FILLER_185_1625 ();
 sg13g2_decap_8 FILLER_185_1632 ();
 sg13g2_decap_8 FILLER_185_1639 ();
 sg13g2_decap_8 FILLER_185_1646 ();
 sg13g2_decap_8 FILLER_185_1653 ();
 sg13g2_decap_8 FILLER_185_1660 ();
 sg13g2_decap_8 FILLER_185_1667 ();
 sg13g2_decap_8 FILLER_185_1674 ();
 sg13g2_decap_8 FILLER_185_1681 ();
 sg13g2_decap_8 FILLER_185_1688 ();
 sg13g2_decap_8 FILLER_185_1695 ();
 sg13g2_decap_8 FILLER_185_1702 ();
 sg13g2_decap_8 FILLER_185_1709 ();
 sg13g2_decap_8 FILLER_185_1716 ();
 sg13g2_decap_8 FILLER_185_1723 ();
 sg13g2_decap_8 FILLER_185_1730 ();
 sg13g2_decap_8 FILLER_185_1737 ();
 sg13g2_decap_8 FILLER_185_1744 ();
 sg13g2_decap_8 FILLER_185_1751 ();
 sg13g2_decap_8 FILLER_185_1758 ();
 sg13g2_fill_2 FILLER_185_1765 ();
 sg13g2_fill_1 FILLER_185_1767 ();
 assign uio_oe[0] = net266;
 assign uio_oe[1] = net267;
 assign uio_oe[2] = net268;
 assign uio_oe[3] = net269;
 assign uio_oe[4] = net270;
 assign uio_oe[5] = net271;
 assign uio_oe[6] = net272;
 assign uio_oe[7] = net10;
 assign uio_out[7] = net11;
endmodule
